magic
tech sky130A
magscale 1 2
timestamp 1732488445
<< obsli1 >>
rect 1104 1071 24840 43537
<< obsm1 >>
rect 14 484 25930 43852
<< metal2 >>
rect 202 44463 258 44623
rect 478 44463 534 44623
rect 754 44463 810 44623
rect 1030 44463 1086 44623
rect 1306 44463 1362 44623
rect 1582 44463 1638 44623
rect 1858 44463 1914 44623
rect 2134 44463 2190 44623
rect 2410 44463 2466 44623
rect 2686 44463 2742 44623
rect 2962 44463 3018 44623
rect 3238 44463 3294 44623
rect 3514 44463 3570 44623
rect 3790 44463 3846 44623
rect 4066 44463 4122 44623
rect 4342 44463 4398 44623
rect 4618 44463 4674 44623
rect 4894 44463 4950 44623
rect 5170 44463 5226 44623
rect 5446 44463 5502 44623
rect 5722 44463 5778 44623
rect 5998 44463 6054 44623
rect 6274 44463 6330 44623
rect 6550 44463 6606 44623
rect 6826 44463 6882 44623
rect 7102 44463 7158 44623
rect 7378 44463 7434 44623
rect 7654 44463 7710 44623
rect 7930 44463 7986 44623
rect 8206 44463 8262 44623
rect 8482 44463 8538 44623
rect 8758 44463 8814 44623
rect 9034 44463 9090 44623
rect 9310 44463 9366 44623
rect 9586 44463 9642 44623
rect 9862 44463 9918 44623
rect 10138 44463 10194 44623
rect 10414 44463 10470 44623
rect 10690 44463 10746 44623
rect 10966 44463 11022 44623
rect 11242 44463 11298 44623
rect 11518 44463 11574 44623
rect 11794 44463 11850 44623
rect 12070 44463 12126 44623
rect 12346 44463 12402 44623
rect 12622 44463 12678 44623
rect 12898 44463 12954 44623
rect 13174 44463 13230 44623
rect 13450 44463 13506 44623
rect 13726 44463 13782 44623
rect 14002 44463 14058 44623
rect 14278 44463 14334 44623
rect 14554 44463 14610 44623
rect 14830 44463 14886 44623
rect 15106 44463 15162 44623
rect 15382 44463 15438 44623
rect 15658 44463 15714 44623
rect 15934 44463 15990 44623
rect 16210 44463 16266 44623
rect 16486 44463 16542 44623
rect 16762 44463 16818 44623
rect 17038 44463 17094 44623
rect 17314 44463 17370 44623
rect 17590 44463 17646 44623
rect 17866 44463 17922 44623
rect 18142 44463 18198 44623
rect 18418 44463 18474 44623
rect 18694 44463 18750 44623
rect 18970 44463 19026 44623
rect 19246 44463 19302 44623
rect 19522 44463 19578 44623
rect 19798 44463 19854 44623
rect 20074 44463 20130 44623
rect 20350 44463 20406 44623
rect 20626 44463 20682 44623
rect 20902 44463 20958 44623
rect 21178 44463 21234 44623
rect 21454 44463 21510 44623
rect 21730 44463 21786 44623
rect 22006 44463 22062 44623
rect 22282 44463 22338 44623
rect 22558 44463 22614 44623
rect 22834 44463 22890 44623
rect 23110 44463 23166 44623
rect 23386 44463 23442 44623
rect 23662 44463 23718 44623
rect 23938 44463 23994 44623
rect 24214 44463 24270 44623
rect 24490 44463 24546 44623
rect 24766 44463 24822 44623
rect 25042 44463 25098 44623
rect 25318 44463 25374 44623
rect 25594 44463 25650 44623
rect 202 0 258 160
rect 478 0 534 160
rect 754 0 810 160
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 0 1638 160
rect 1858 0 1914 160
rect 2134 0 2190 160
rect 2410 0 2466 160
rect 2686 0 2742 160
rect 2962 0 3018 160
rect 3238 0 3294 160
rect 3514 0 3570 160
rect 3790 0 3846 160
rect 4066 0 4122 160
rect 4342 0 4398 160
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5170 0 5226 160
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11242 0 11298 160
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 0 14610 160
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 0 19854 160
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20902 0 20958 160
rect 21178 0 21234 160
rect 21454 0 21510 160
rect 21730 0 21786 160
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 0 22614 160
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24766 0 24822 160
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
<< obsm2 >>
rect 20 44407 146 44577
rect 314 44407 422 44577
rect 590 44407 698 44577
rect 866 44407 974 44577
rect 1142 44407 1250 44577
rect 1418 44407 1526 44577
rect 1694 44407 1802 44577
rect 1970 44407 2078 44577
rect 2246 44407 2354 44577
rect 2522 44407 2630 44577
rect 2798 44407 2906 44577
rect 3074 44407 3182 44577
rect 3350 44407 3458 44577
rect 3626 44407 3734 44577
rect 3902 44407 4010 44577
rect 4178 44407 4286 44577
rect 4454 44407 4562 44577
rect 4730 44407 4838 44577
rect 5006 44407 5114 44577
rect 5282 44407 5390 44577
rect 5558 44407 5666 44577
rect 5834 44407 5942 44577
rect 6110 44407 6218 44577
rect 6386 44407 6494 44577
rect 6662 44407 6770 44577
rect 6938 44407 7046 44577
rect 7214 44407 7322 44577
rect 7490 44407 7598 44577
rect 7766 44407 7874 44577
rect 8042 44407 8150 44577
rect 8318 44407 8426 44577
rect 8594 44407 8702 44577
rect 8870 44407 8978 44577
rect 9146 44407 9254 44577
rect 9422 44407 9530 44577
rect 9698 44407 9806 44577
rect 9974 44407 10082 44577
rect 10250 44407 10358 44577
rect 10526 44407 10634 44577
rect 10802 44407 10910 44577
rect 11078 44407 11186 44577
rect 11354 44407 11462 44577
rect 11630 44407 11738 44577
rect 11906 44407 12014 44577
rect 12182 44407 12290 44577
rect 12458 44407 12566 44577
rect 12734 44407 12842 44577
rect 13010 44407 13118 44577
rect 13286 44407 13394 44577
rect 13562 44407 13670 44577
rect 13838 44407 13946 44577
rect 14114 44407 14222 44577
rect 14390 44407 14498 44577
rect 14666 44407 14774 44577
rect 14942 44407 15050 44577
rect 15218 44407 15326 44577
rect 15494 44407 15602 44577
rect 15770 44407 15878 44577
rect 16046 44407 16154 44577
rect 16322 44407 16430 44577
rect 16598 44407 16706 44577
rect 16874 44407 16982 44577
rect 17150 44407 17258 44577
rect 17426 44407 17534 44577
rect 17702 44407 17810 44577
rect 17978 44407 18086 44577
rect 18254 44407 18362 44577
rect 18530 44407 18638 44577
rect 18806 44407 18914 44577
rect 19082 44407 19190 44577
rect 19358 44407 19466 44577
rect 19634 44407 19742 44577
rect 19910 44407 20018 44577
rect 20186 44407 20294 44577
rect 20462 44407 20570 44577
rect 20738 44407 20846 44577
rect 21014 44407 21122 44577
rect 21290 44407 21398 44577
rect 21566 44407 21674 44577
rect 21842 44407 21950 44577
rect 22118 44407 22226 44577
rect 22394 44407 22502 44577
rect 22670 44407 22778 44577
rect 22946 44407 23054 44577
rect 23222 44407 23330 44577
rect 23498 44407 23606 44577
rect 23774 44407 23882 44577
rect 24050 44407 24158 44577
rect 24326 44407 24434 44577
rect 24602 44407 24710 44577
rect 24878 44407 24986 44577
rect 25154 44407 25262 44577
rect 25430 44407 25538 44577
rect 25706 44407 25924 44577
rect 20 216 25924 44407
rect 20 54 146 216
rect 314 54 422 216
rect 590 54 698 216
rect 866 54 974 216
rect 1142 54 1250 216
rect 1418 54 1526 216
rect 1694 54 1802 216
rect 1970 54 2078 216
rect 2246 54 2354 216
rect 2522 54 2630 216
rect 2798 54 2906 216
rect 3074 54 3182 216
rect 3350 54 3458 216
rect 3626 54 3734 216
rect 3902 54 4010 216
rect 4178 54 4286 216
rect 4454 54 4562 216
rect 4730 54 4838 216
rect 5006 54 5114 216
rect 5282 54 5390 216
rect 5558 54 5666 216
rect 5834 54 5942 216
rect 6110 54 6218 216
rect 6386 54 6494 216
rect 6662 54 6770 216
rect 6938 54 7046 216
rect 7214 54 7322 216
rect 7490 54 7598 216
rect 7766 54 7874 216
rect 8042 54 8150 216
rect 8318 54 8426 216
rect 8594 54 8702 216
rect 8870 54 8978 216
rect 9146 54 9254 216
rect 9422 54 9530 216
rect 9698 54 9806 216
rect 9974 54 10082 216
rect 10250 54 10358 216
rect 10526 54 10634 216
rect 10802 54 10910 216
rect 11078 54 11186 216
rect 11354 54 11462 216
rect 11630 54 11738 216
rect 11906 54 12014 216
rect 12182 54 12290 216
rect 12458 54 12566 216
rect 12734 54 12842 216
rect 13010 54 13118 216
rect 13286 54 13394 216
rect 13562 54 13670 216
rect 13838 54 13946 216
rect 14114 54 14222 216
rect 14390 54 14498 216
rect 14666 54 14774 216
rect 14942 54 15050 216
rect 15218 54 15326 216
rect 15494 54 15602 216
rect 15770 54 15878 216
rect 16046 54 16154 216
rect 16322 54 16430 216
rect 16598 54 16706 216
rect 16874 54 16982 216
rect 17150 54 17258 216
rect 17426 54 17534 216
rect 17702 54 17810 216
rect 17978 54 18086 216
rect 18254 54 18362 216
rect 18530 54 18638 216
rect 18806 54 18914 216
rect 19082 54 19190 216
rect 19358 54 19466 216
rect 19634 54 19742 216
rect 19910 54 20018 216
rect 20186 54 20294 216
rect 20462 54 20570 216
rect 20738 54 20846 216
rect 21014 54 21122 216
rect 21290 54 21398 216
rect 21566 54 21674 216
rect 21842 54 21950 216
rect 22118 54 22226 216
rect 22394 54 22502 216
rect 22670 54 22778 216
rect 22946 54 23054 216
rect 23222 54 23330 216
rect 23498 54 23606 216
rect 23774 54 23882 216
rect 24050 54 24158 216
rect 24326 54 24434 216
rect 24602 54 24710 216
rect 24878 54 24986 216
rect 25154 54 25262 216
rect 25430 54 25538 216
rect 25706 54 25924 216
<< metal3 >>
rect 25840 43528 26000 43648
rect 25840 42984 26000 43104
rect 25840 42440 26000 42560
rect 25840 41896 26000 42016
rect 25840 41352 26000 41472
rect 25840 40808 26000 40928
rect 25840 40264 26000 40384
rect 25840 39720 26000 39840
rect 0 39448 160 39568
rect 0 39176 160 39296
rect 25840 39176 26000 39296
rect 0 38904 160 39024
rect 0 38632 160 38752
rect 25840 38632 26000 38752
rect 0 38360 160 38480
rect 0 38088 160 38208
rect 25840 38088 26000 38208
rect 0 37816 160 37936
rect 0 37544 160 37664
rect 25840 37544 26000 37664
rect 0 37272 160 37392
rect 0 37000 160 37120
rect 25840 37000 26000 37120
rect 0 36728 160 36848
rect 0 36456 160 36576
rect 25840 36456 26000 36576
rect 0 36184 160 36304
rect 0 35912 160 36032
rect 25840 35912 26000 36032
rect 0 35640 160 35760
rect 0 35368 160 35488
rect 25840 35368 26000 35488
rect 0 35096 160 35216
rect 0 34824 160 34944
rect 25840 34824 26000 34944
rect 0 34552 160 34672
rect 0 34280 160 34400
rect 25840 34280 26000 34400
rect 0 34008 160 34128
rect 0 33736 160 33856
rect 25840 33736 26000 33856
rect 0 33464 160 33584
rect 0 33192 160 33312
rect 25840 33192 26000 33312
rect 0 32920 160 33040
rect 0 32648 160 32768
rect 25840 32648 26000 32768
rect 0 32376 160 32496
rect 0 32104 160 32224
rect 25840 32104 26000 32224
rect 0 31832 160 31952
rect 0 31560 160 31680
rect 25840 31560 26000 31680
rect 0 31288 160 31408
rect 0 31016 160 31136
rect 25840 31016 26000 31136
rect 0 30744 160 30864
rect 0 30472 160 30592
rect 25840 30472 26000 30592
rect 0 30200 160 30320
rect 0 29928 160 30048
rect 25840 29928 26000 30048
rect 0 29656 160 29776
rect 0 29384 160 29504
rect 25840 29384 26000 29504
rect 0 29112 160 29232
rect 0 28840 160 28960
rect 25840 28840 26000 28960
rect 0 28568 160 28688
rect 0 28296 160 28416
rect 25840 28296 26000 28416
rect 0 28024 160 28144
rect 0 27752 160 27872
rect 25840 27752 26000 27872
rect 0 27480 160 27600
rect 0 27208 160 27328
rect 25840 27208 26000 27328
rect 0 26936 160 27056
rect 0 26664 160 26784
rect 25840 26664 26000 26784
rect 0 26392 160 26512
rect 0 26120 160 26240
rect 25840 26120 26000 26240
rect 0 25848 160 25968
rect 0 25576 160 25696
rect 25840 25576 26000 25696
rect 0 25304 160 25424
rect 0 25032 160 25152
rect 25840 25032 26000 25152
rect 0 24760 160 24880
rect 0 24488 160 24608
rect 25840 24488 26000 24608
rect 0 24216 160 24336
rect 0 23944 160 24064
rect 25840 23944 26000 24064
rect 0 23672 160 23792
rect 0 23400 160 23520
rect 25840 23400 26000 23520
rect 0 23128 160 23248
rect 0 22856 160 22976
rect 25840 22856 26000 22976
rect 0 22584 160 22704
rect 0 22312 160 22432
rect 25840 22312 26000 22432
rect 0 22040 160 22160
rect 0 21768 160 21888
rect 25840 21768 26000 21888
rect 0 21496 160 21616
rect 0 21224 160 21344
rect 25840 21224 26000 21344
rect 0 20952 160 21072
rect 0 20680 160 20800
rect 25840 20680 26000 20800
rect 0 20408 160 20528
rect 0 20136 160 20256
rect 25840 20136 26000 20256
rect 0 19864 160 19984
rect 0 19592 160 19712
rect 25840 19592 26000 19712
rect 0 19320 160 19440
rect 0 19048 160 19168
rect 25840 19048 26000 19168
rect 0 18776 160 18896
rect 0 18504 160 18624
rect 25840 18504 26000 18624
rect 0 18232 160 18352
rect 0 17960 160 18080
rect 25840 17960 26000 18080
rect 0 17688 160 17808
rect 0 17416 160 17536
rect 25840 17416 26000 17536
rect 0 17144 160 17264
rect 0 16872 160 16992
rect 25840 16872 26000 16992
rect 0 16600 160 16720
rect 0 16328 160 16448
rect 25840 16328 26000 16448
rect 0 16056 160 16176
rect 0 15784 160 15904
rect 25840 15784 26000 15904
rect 0 15512 160 15632
rect 0 15240 160 15360
rect 25840 15240 26000 15360
rect 0 14968 160 15088
rect 0 14696 160 14816
rect 25840 14696 26000 14816
rect 0 14424 160 14544
rect 0 14152 160 14272
rect 25840 14152 26000 14272
rect 0 13880 160 14000
rect 0 13608 160 13728
rect 25840 13608 26000 13728
rect 0 13336 160 13456
rect 0 13064 160 13184
rect 25840 13064 26000 13184
rect 0 12792 160 12912
rect 0 12520 160 12640
rect 25840 12520 26000 12640
rect 0 12248 160 12368
rect 0 11976 160 12096
rect 25840 11976 26000 12096
rect 0 11704 160 11824
rect 0 11432 160 11552
rect 25840 11432 26000 11552
rect 0 11160 160 11280
rect 0 10888 160 11008
rect 25840 10888 26000 11008
rect 0 10616 160 10736
rect 0 10344 160 10464
rect 25840 10344 26000 10464
rect 0 10072 160 10192
rect 0 9800 160 9920
rect 25840 9800 26000 9920
rect 0 9528 160 9648
rect 0 9256 160 9376
rect 25840 9256 26000 9376
rect 0 8984 160 9104
rect 0 8712 160 8832
rect 25840 8712 26000 8832
rect 0 8440 160 8560
rect 0 8168 160 8288
rect 25840 8168 26000 8288
rect 0 7896 160 8016
rect 0 7624 160 7744
rect 25840 7624 26000 7744
rect 0 7352 160 7472
rect 0 7080 160 7200
rect 25840 7080 26000 7200
rect 0 6808 160 6928
rect 0 6536 160 6656
rect 25840 6536 26000 6656
rect 0 6264 160 6384
rect 0 5992 160 6112
rect 25840 5992 26000 6112
rect 0 5720 160 5840
rect 0 5448 160 5568
rect 25840 5448 26000 5568
rect 0 5176 160 5296
rect 0 4904 160 5024
rect 25840 4904 26000 5024
rect 25840 4360 26000 4480
rect 25840 3816 26000 3936
rect 25840 3272 26000 3392
rect 25840 2728 26000 2848
rect 25840 2184 26000 2304
rect 25840 1640 26000 1760
rect 25840 1096 26000 1216
rect 25840 552 26000 672
<< obsm3 >>
rect 160 43728 25840 44573
rect 160 43448 25760 43728
rect 160 43184 25840 43448
rect 160 42904 25760 43184
rect 160 42640 25840 42904
rect 160 42360 25760 42640
rect 160 42096 25840 42360
rect 160 41816 25760 42096
rect 160 41552 25840 41816
rect 160 41272 25760 41552
rect 160 41008 25840 41272
rect 160 40728 25760 41008
rect 160 40464 25840 40728
rect 160 40184 25760 40464
rect 160 39920 25840 40184
rect 160 39648 25760 39920
rect 240 39640 25760 39648
rect 240 39376 25840 39640
rect 240 39096 25760 39376
rect 240 38832 25840 39096
rect 240 38552 25760 38832
rect 240 38288 25840 38552
rect 240 38008 25760 38288
rect 240 37744 25840 38008
rect 240 37464 25760 37744
rect 240 37200 25840 37464
rect 240 36920 25760 37200
rect 240 36656 25840 36920
rect 240 36376 25760 36656
rect 240 36112 25840 36376
rect 240 35832 25760 36112
rect 240 35568 25840 35832
rect 240 35288 25760 35568
rect 240 35024 25840 35288
rect 240 34744 25760 35024
rect 240 34480 25840 34744
rect 240 34200 25760 34480
rect 240 33936 25840 34200
rect 240 33656 25760 33936
rect 240 33392 25840 33656
rect 240 33112 25760 33392
rect 240 32848 25840 33112
rect 240 32568 25760 32848
rect 240 32304 25840 32568
rect 240 32024 25760 32304
rect 240 31760 25840 32024
rect 240 31480 25760 31760
rect 240 31216 25840 31480
rect 240 30936 25760 31216
rect 240 30672 25840 30936
rect 240 30392 25760 30672
rect 240 30128 25840 30392
rect 240 29848 25760 30128
rect 240 29584 25840 29848
rect 240 29304 25760 29584
rect 240 29040 25840 29304
rect 240 28760 25760 29040
rect 240 28496 25840 28760
rect 240 28216 25760 28496
rect 240 27952 25840 28216
rect 240 27672 25760 27952
rect 240 27408 25840 27672
rect 240 27128 25760 27408
rect 240 26864 25840 27128
rect 240 26584 25760 26864
rect 240 26320 25840 26584
rect 240 26040 25760 26320
rect 240 25776 25840 26040
rect 240 25496 25760 25776
rect 240 25232 25840 25496
rect 240 24952 25760 25232
rect 240 24688 25840 24952
rect 240 24408 25760 24688
rect 240 24144 25840 24408
rect 240 23864 25760 24144
rect 240 23600 25840 23864
rect 240 23320 25760 23600
rect 240 23056 25840 23320
rect 240 22776 25760 23056
rect 240 22512 25840 22776
rect 240 22232 25760 22512
rect 240 21968 25840 22232
rect 240 21688 25760 21968
rect 240 21424 25840 21688
rect 240 21144 25760 21424
rect 240 20880 25840 21144
rect 240 20600 25760 20880
rect 240 20336 25840 20600
rect 240 20056 25760 20336
rect 240 19792 25840 20056
rect 240 19512 25760 19792
rect 240 19248 25840 19512
rect 240 18968 25760 19248
rect 240 18704 25840 18968
rect 240 18424 25760 18704
rect 240 18160 25840 18424
rect 240 17880 25760 18160
rect 240 17616 25840 17880
rect 240 17336 25760 17616
rect 240 17072 25840 17336
rect 240 16792 25760 17072
rect 240 16528 25840 16792
rect 240 16248 25760 16528
rect 240 15984 25840 16248
rect 240 15704 25760 15984
rect 240 15440 25840 15704
rect 240 15160 25760 15440
rect 240 14896 25840 15160
rect 240 14616 25760 14896
rect 240 14352 25840 14616
rect 240 14072 25760 14352
rect 240 13808 25840 14072
rect 240 13528 25760 13808
rect 240 13264 25840 13528
rect 240 12984 25760 13264
rect 240 12720 25840 12984
rect 240 12440 25760 12720
rect 240 12176 25840 12440
rect 240 11896 25760 12176
rect 240 11632 25840 11896
rect 240 11352 25760 11632
rect 240 11088 25840 11352
rect 240 10808 25760 11088
rect 240 10544 25840 10808
rect 240 10264 25760 10544
rect 240 10000 25840 10264
rect 240 9720 25760 10000
rect 240 9456 25840 9720
rect 240 9176 25760 9456
rect 240 8912 25840 9176
rect 240 8632 25760 8912
rect 240 8368 25840 8632
rect 240 8088 25760 8368
rect 240 7824 25840 8088
rect 240 7544 25760 7824
rect 240 7280 25840 7544
rect 240 7000 25760 7280
rect 240 6736 25840 7000
rect 240 6456 25760 6736
rect 240 6192 25840 6456
rect 240 5912 25760 6192
rect 240 5648 25840 5912
rect 240 5368 25760 5648
rect 240 5104 25840 5368
rect 240 4824 25760 5104
rect 160 4560 25840 4824
rect 160 4280 25760 4560
rect 160 4016 25840 4280
rect 160 3736 25760 4016
rect 160 3472 25840 3736
rect 160 3192 25760 3472
rect 160 2928 25840 3192
rect 160 2648 25760 2928
rect 160 2384 25840 2648
rect 160 2104 25760 2384
rect 160 1840 25840 2104
rect 160 1560 25760 1840
rect 160 1296 25840 1560
rect 160 1016 25760 1296
rect 160 752 25840 1016
rect 160 579 25760 752
<< metal4 >>
rect 3911 1040 4231 43568
rect 6878 1040 7198 43568
rect 9845 1040 10165 43568
rect 12812 1040 13132 43568
rect 15779 1040 16099 43568
rect 18746 1040 19066 43568
rect 21713 1040 22033 43568
rect 24680 1040 25000 43568
<< obsm4 >>
rect 611 43648 23309 44573
rect 611 960 3831 43648
rect 4311 960 6798 43648
rect 7278 960 9765 43648
rect 10245 960 12732 43648
rect 13212 960 15699 43648
rect 16179 960 18666 43648
rect 19146 960 21633 43648
rect 22113 960 23309 43648
rect 611 851 23309 960
<< obsm5 >>
rect 3060 21940 12764 22260
<< labels >>
rlabel metal3 s 25840 9256 26000 9376 6 Config_accessC_bit0
port 1 nsew signal output
rlabel metal3 s 25840 9800 26000 9920 6 Config_accessC_bit1
port 2 nsew signal output
rlabel metal3 s 25840 10344 26000 10464 6 Config_accessC_bit2
port 3 nsew signal output
rlabel metal3 s 25840 10888 26000 11008 6 Config_accessC_bit3
port 4 nsew signal output
rlabel metal3 s 0 17960 160 18080 6 E1END[0]
port 5 nsew signal input
rlabel metal3 s 0 18232 160 18352 6 E1END[1]
port 6 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 E1END[2]
port 7 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 E1END[3]
port 8 nsew signal input
rlabel metal3 s 0 21224 160 21344 6 E2END[0]
port 9 nsew signal input
rlabel metal3 s 0 21496 160 21616 6 E2END[1]
port 10 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 E2END[2]
port 11 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 E2END[3]
port 12 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 E2END[4]
port 13 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 E2END[5]
port 14 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 E2END[6]
port 15 nsew signal input
rlabel metal3 s 0 23128 160 23248 6 E2END[7]
port 16 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 E2MID[0]
port 17 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 E2MID[1]
port 18 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 E2MID[2]
port 19 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 E2MID[3]
port 20 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 E2MID[4]
port 21 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 E2MID[5]
port 22 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 E2MID[6]
port 23 nsew signal input
rlabel metal3 s 0 20952 160 21072 6 E2MID[7]
port 24 nsew signal input
rlabel metal3 s 0 27752 160 27872 6 E6END[0]
port 25 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 E6END[10]
port 26 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 E6END[11]
port 27 nsew signal input
rlabel metal3 s 0 28024 160 28144 6 E6END[1]
port 28 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 E6END[2]
port 29 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 E6END[3]
port 30 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 E6END[4]
port 31 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 E6END[5]
port 32 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 E6END[6]
port 33 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 E6END[7]
port 34 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 E6END[8]
port 35 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 E6END[9]
port 36 nsew signal input
rlabel metal3 s 0 23400 160 23520 6 EE4END[0]
port 37 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 EE4END[10]
port 38 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 EE4END[11]
port 39 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 EE4END[12]
port 40 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 EE4END[13]
port 41 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 EE4END[14]
port 42 nsew signal input
rlabel metal3 s 0 27480 160 27600 6 EE4END[15]
port 43 nsew signal input
rlabel metal3 s 0 23672 160 23792 6 EE4END[1]
port 44 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 EE4END[2]
port 45 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 EE4END[3]
port 46 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 EE4END[4]
port 47 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 EE4END[5]
port 48 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 EE4END[6]
port 49 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 EE4END[7]
port 50 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 EE4END[8]
port 51 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 EE4END[9]
port 52 nsew signal input
rlabel metal3 s 25840 15784 26000 15904 6 FAB2RAM_A0_O0
port 53 nsew signal output
rlabel metal3 s 25840 16328 26000 16448 6 FAB2RAM_A0_O1
port 54 nsew signal output
rlabel metal3 s 25840 16872 26000 16992 6 FAB2RAM_A0_O2
port 55 nsew signal output
rlabel metal3 s 25840 17416 26000 17536 6 FAB2RAM_A0_O3
port 56 nsew signal output
rlabel metal3 s 25840 13608 26000 13728 6 FAB2RAM_A1_O0
port 57 nsew signal output
rlabel metal3 s 25840 14152 26000 14272 6 FAB2RAM_A1_O1
port 58 nsew signal output
rlabel metal3 s 25840 14696 26000 14816 6 FAB2RAM_A1_O2
port 59 nsew signal output
rlabel metal3 s 25840 15240 26000 15360 6 FAB2RAM_A1_O3
port 60 nsew signal output
rlabel metal3 s 25840 11432 26000 11552 6 FAB2RAM_C_O0
port 61 nsew signal output
rlabel metal3 s 25840 11976 26000 12096 6 FAB2RAM_C_O1
port 62 nsew signal output
rlabel metal3 s 25840 12520 26000 12640 6 FAB2RAM_C_O2
port 63 nsew signal output
rlabel metal3 s 25840 13064 26000 13184 6 FAB2RAM_C_O3
port 64 nsew signal output
rlabel metal3 s 25840 24488 26000 24608 6 FAB2RAM_D0_O0
port 65 nsew signal output
rlabel metal3 s 25840 25032 26000 25152 6 FAB2RAM_D0_O1
port 66 nsew signal output
rlabel metal3 s 25840 25576 26000 25696 6 FAB2RAM_D0_O2
port 67 nsew signal output
rlabel metal3 s 25840 26120 26000 26240 6 FAB2RAM_D0_O3
port 68 nsew signal output
rlabel metal3 s 25840 22312 26000 22432 6 FAB2RAM_D1_O0
port 69 nsew signal output
rlabel metal3 s 25840 22856 26000 22976 6 FAB2RAM_D1_O1
port 70 nsew signal output
rlabel metal3 s 25840 23400 26000 23520 6 FAB2RAM_D1_O2
port 71 nsew signal output
rlabel metal3 s 25840 23944 26000 24064 6 FAB2RAM_D1_O3
port 72 nsew signal output
rlabel metal3 s 25840 20136 26000 20256 6 FAB2RAM_D2_O0
port 73 nsew signal output
rlabel metal3 s 25840 20680 26000 20800 6 FAB2RAM_D2_O1
port 74 nsew signal output
rlabel metal3 s 25840 21224 26000 21344 6 FAB2RAM_D2_O2
port 75 nsew signal output
rlabel metal3 s 25840 21768 26000 21888 6 FAB2RAM_D2_O3
port 76 nsew signal output
rlabel metal3 s 25840 17960 26000 18080 6 FAB2RAM_D3_O0
port 77 nsew signal output
rlabel metal3 s 25840 18504 26000 18624 6 FAB2RAM_D3_O1
port 78 nsew signal output
rlabel metal3 s 25840 19048 26000 19168 6 FAB2RAM_D3_O2
port 79 nsew signal output
rlabel metal3 s 25840 19592 26000 19712 6 FAB2RAM_D3_O3
port 80 nsew signal output
rlabel metal3 s 0 31016 160 31136 6 FrameData[0]
port 81 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 FrameData[10]
port 82 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 FrameData[11]
port 83 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 FrameData[12]
port 84 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 FrameData[13]
port 85 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 FrameData[14]
port 86 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 FrameData[15]
port 87 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 FrameData[16]
port 88 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 FrameData[17]
port 89 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 FrameData[18]
port 90 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 FrameData[19]
port 91 nsew signal input
rlabel metal3 s 0 31288 160 31408 6 FrameData[1]
port 92 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 FrameData[20]
port 93 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 FrameData[21]
port 94 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 FrameData[22]
port 95 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 FrameData[23]
port 96 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 FrameData[24]
port 97 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 FrameData[25]
port 98 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 FrameData[26]
port 99 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 FrameData[27]
port 100 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 FrameData[28]
port 101 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 FrameData[29]
port 102 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 FrameData[2]
port 103 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 FrameData[30]
port 104 nsew signal input
rlabel metal3 s 0 39448 160 39568 6 FrameData[31]
port 105 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 FrameData[3]
port 106 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 FrameData[4]
port 107 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 FrameData[5]
port 108 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 FrameData[6]
port 109 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 FrameData[7]
port 110 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 FrameData[8]
port 111 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 FrameData[9]
port 112 nsew signal input
rlabel metal3 s 25840 26664 26000 26784 6 FrameData_O[0]
port 113 nsew signal output
rlabel metal3 s 25840 32104 26000 32224 6 FrameData_O[10]
port 114 nsew signal output
rlabel metal3 s 25840 32648 26000 32768 6 FrameData_O[11]
port 115 nsew signal output
rlabel metal3 s 25840 33192 26000 33312 6 FrameData_O[12]
port 116 nsew signal output
rlabel metal3 s 25840 33736 26000 33856 6 FrameData_O[13]
port 117 nsew signal output
rlabel metal3 s 25840 34280 26000 34400 6 FrameData_O[14]
port 118 nsew signal output
rlabel metal3 s 25840 34824 26000 34944 6 FrameData_O[15]
port 119 nsew signal output
rlabel metal3 s 25840 35368 26000 35488 6 FrameData_O[16]
port 120 nsew signal output
rlabel metal3 s 25840 35912 26000 36032 6 FrameData_O[17]
port 121 nsew signal output
rlabel metal3 s 25840 36456 26000 36576 6 FrameData_O[18]
port 122 nsew signal output
rlabel metal3 s 25840 37000 26000 37120 6 FrameData_O[19]
port 123 nsew signal output
rlabel metal3 s 25840 27208 26000 27328 6 FrameData_O[1]
port 124 nsew signal output
rlabel metal3 s 25840 37544 26000 37664 6 FrameData_O[20]
port 125 nsew signal output
rlabel metal3 s 25840 38088 26000 38208 6 FrameData_O[21]
port 126 nsew signal output
rlabel metal3 s 25840 38632 26000 38752 6 FrameData_O[22]
port 127 nsew signal output
rlabel metal3 s 25840 39176 26000 39296 6 FrameData_O[23]
port 128 nsew signal output
rlabel metal3 s 25840 39720 26000 39840 6 FrameData_O[24]
port 129 nsew signal output
rlabel metal3 s 25840 40264 26000 40384 6 FrameData_O[25]
port 130 nsew signal output
rlabel metal3 s 25840 40808 26000 40928 6 FrameData_O[26]
port 131 nsew signal output
rlabel metal3 s 25840 41352 26000 41472 6 FrameData_O[27]
port 132 nsew signal output
rlabel metal3 s 25840 41896 26000 42016 6 FrameData_O[28]
port 133 nsew signal output
rlabel metal3 s 25840 42440 26000 42560 6 FrameData_O[29]
port 134 nsew signal output
rlabel metal3 s 25840 27752 26000 27872 6 FrameData_O[2]
port 135 nsew signal output
rlabel metal3 s 25840 42984 26000 43104 6 FrameData_O[30]
port 136 nsew signal output
rlabel metal3 s 25840 43528 26000 43648 6 FrameData_O[31]
port 137 nsew signal output
rlabel metal3 s 25840 28296 26000 28416 6 FrameData_O[3]
port 138 nsew signal output
rlabel metal3 s 25840 28840 26000 28960 6 FrameData_O[4]
port 139 nsew signal output
rlabel metal3 s 25840 29384 26000 29504 6 FrameData_O[5]
port 140 nsew signal output
rlabel metal3 s 25840 29928 26000 30048 6 FrameData_O[6]
port 141 nsew signal output
rlabel metal3 s 25840 30472 26000 30592 6 FrameData_O[7]
port 142 nsew signal output
rlabel metal3 s 25840 31016 26000 31136 6 FrameData_O[8]
port 143 nsew signal output
rlabel metal3 s 25840 31560 26000 31680 6 FrameData_O[9]
port 144 nsew signal output
rlabel metal2 s 20350 0 20406 160 6 FrameStrobe[0]
port 145 nsew signal input
rlabel metal2 s 23110 0 23166 160 6 FrameStrobe[10]
port 146 nsew signal input
rlabel metal2 s 23386 0 23442 160 6 FrameStrobe[11]
port 147 nsew signal input
rlabel metal2 s 23662 0 23718 160 6 FrameStrobe[12]
port 148 nsew signal input
rlabel metal2 s 23938 0 23994 160 6 FrameStrobe[13]
port 149 nsew signal input
rlabel metal2 s 24214 0 24270 160 6 FrameStrobe[14]
port 150 nsew signal input
rlabel metal2 s 24490 0 24546 160 6 FrameStrobe[15]
port 151 nsew signal input
rlabel metal2 s 24766 0 24822 160 6 FrameStrobe[16]
port 152 nsew signal input
rlabel metal2 s 25042 0 25098 160 6 FrameStrobe[17]
port 153 nsew signal input
rlabel metal2 s 25318 0 25374 160 6 FrameStrobe[18]
port 154 nsew signal input
rlabel metal2 s 25594 0 25650 160 6 FrameStrobe[19]
port 155 nsew signal input
rlabel metal2 s 20626 0 20682 160 6 FrameStrobe[1]
port 156 nsew signal input
rlabel metal2 s 20902 0 20958 160 6 FrameStrobe[2]
port 157 nsew signal input
rlabel metal2 s 21178 0 21234 160 6 FrameStrobe[3]
port 158 nsew signal input
rlabel metal2 s 21454 0 21510 160 6 FrameStrobe[4]
port 159 nsew signal input
rlabel metal2 s 21730 0 21786 160 6 FrameStrobe[5]
port 160 nsew signal input
rlabel metal2 s 22006 0 22062 160 6 FrameStrobe[6]
port 161 nsew signal input
rlabel metal2 s 22282 0 22338 160 6 FrameStrobe[7]
port 162 nsew signal input
rlabel metal2 s 22558 0 22614 160 6 FrameStrobe[8]
port 163 nsew signal input
rlabel metal2 s 22834 0 22890 160 6 FrameStrobe[9]
port 164 nsew signal input
rlabel metal2 s 20350 44463 20406 44623 6 FrameStrobe_O[0]
port 165 nsew signal output
rlabel metal2 s 23110 44463 23166 44623 6 FrameStrobe_O[10]
port 166 nsew signal output
rlabel metal2 s 23386 44463 23442 44623 6 FrameStrobe_O[11]
port 167 nsew signal output
rlabel metal2 s 23662 44463 23718 44623 6 FrameStrobe_O[12]
port 168 nsew signal output
rlabel metal2 s 23938 44463 23994 44623 6 FrameStrobe_O[13]
port 169 nsew signal output
rlabel metal2 s 24214 44463 24270 44623 6 FrameStrobe_O[14]
port 170 nsew signal output
rlabel metal2 s 24490 44463 24546 44623 6 FrameStrobe_O[15]
port 171 nsew signal output
rlabel metal2 s 24766 44463 24822 44623 6 FrameStrobe_O[16]
port 172 nsew signal output
rlabel metal2 s 25042 44463 25098 44623 6 FrameStrobe_O[17]
port 173 nsew signal output
rlabel metal2 s 25318 44463 25374 44623 6 FrameStrobe_O[18]
port 174 nsew signal output
rlabel metal2 s 25594 44463 25650 44623 6 FrameStrobe_O[19]
port 175 nsew signal output
rlabel metal2 s 20626 44463 20682 44623 6 FrameStrobe_O[1]
port 176 nsew signal output
rlabel metal2 s 20902 44463 20958 44623 6 FrameStrobe_O[2]
port 177 nsew signal output
rlabel metal2 s 21178 44463 21234 44623 6 FrameStrobe_O[3]
port 178 nsew signal output
rlabel metal2 s 21454 44463 21510 44623 6 FrameStrobe_O[4]
port 179 nsew signal output
rlabel metal2 s 21730 44463 21786 44623 6 FrameStrobe_O[5]
port 180 nsew signal output
rlabel metal2 s 22006 44463 22062 44623 6 FrameStrobe_O[6]
port 181 nsew signal output
rlabel metal2 s 22282 44463 22338 44623 6 FrameStrobe_O[7]
port 182 nsew signal output
rlabel metal2 s 22558 44463 22614 44623 6 FrameStrobe_O[8]
port 183 nsew signal output
rlabel metal2 s 22834 44463 22890 44623 6 FrameStrobe_O[9]
port 184 nsew signal output
rlabel metal2 s 202 44463 258 44623 6 N1BEG[0]
port 185 nsew signal output
rlabel metal2 s 478 44463 534 44623 6 N1BEG[1]
port 186 nsew signal output
rlabel metal2 s 754 44463 810 44623 6 N1BEG[2]
port 187 nsew signal output
rlabel metal2 s 1030 44463 1086 44623 6 N1BEG[3]
port 188 nsew signal output
rlabel metal2 s 202 0 258 160 6 N1END[0]
port 189 nsew signal input
rlabel metal2 s 478 0 534 160 6 N1END[1]
port 190 nsew signal input
rlabel metal2 s 754 0 810 160 6 N1END[2]
port 191 nsew signal input
rlabel metal2 s 1030 0 1086 160 6 N1END[3]
port 192 nsew signal input
rlabel metal2 s 1306 44463 1362 44623 6 N2BEG[0]
port 193 nsew signal output
rlabel metal2 s 1582 44463 1638 44623 6 N2BEG[1]
port 194 nsew signal output
rlabel metal2 s 1858 44463 1914 44623 6 N2BEG[2]
port 195 nsew signal output
rlabel metal2 s 2134 44463 2190 44623 6 N2BEG[3]
port 196 nsew signal output
rlabel metal2 s 2410 44463 2466 44623 6 N2BEG[4]
port 197 nsew signal output
rlabel metal2 s 2686 44463 2742 44623 6 N2BEG[5]
port 198 nsew signal output
rlabel metal2 s 2962 44463 3018 44623 6 N2BEG[6]
port 199 nsew signal output
rlabel metal2 s 3238 44463 3294 44623 6 N2BEG[7]
port 200 nsew signal output
rlabel metal2 s 3514 44463 3570 44623 6 N2BEGb[0]
port 201 nsew signal output
rlabel metal2 s 3790 44463 3846 44623 6 N2BEGb[1]
port 202 nsew signal output
rlabel metal2 s 4066 44463 4122 44623 6 N2BEGb[2]
port 203 nsew signal output
rlabel metal2 s 4342 44463 4398 44623 6 N2BEGb[3]
port 204 nsew signal output
rlabel metal2 s 4618 44463 4674 44623 6 N2BEGb[4]
port 205 nsew signal output
rlabel metal2 s 4894 44463 4950 44623 6 N2BEGb[5]
port 206 nsew signal output
rlabel metal2 s 5170 44463 5226 44623 6 N2BEGb[6]
port 207 nsew signal output
rlabel metal2 s 5446 44463 5502 44623 6 N2BEGb[7]
port 208 nsew signal output
rlabel metal2 s 3514 0 3570 160 6 N2END[0]
port 209 nsew signal input
rlabel metal2 s 3790 0 3846 160 6 N2END[1]
port 210 nsew signal input
rlabel metal2 s 4066 0 4122 160 6 N2END[2]
port 211 nsew signal input
rlabel metal2 s 4342 0 4398 160 6 N2END[3]
port 212 nsew signal input
rlabel metal2 s 4618 0 4674 160 6 N2END[4]
port 213 nsew signal input
rlabel metal2 s 4894 0 4950 160 6 N2END[5]
port 214 nsew signal input
rlabel metal2 s 5170 0 5226 160 6 N2END[6]
port 215 nsew signal input
rlabel metal2 s 5446 0 5502 160 6 N2END[7]
port 216 nsew signal input
rlabel metal2 s 1306 0 1362 160 6 N2MID[0]
port 217 nsew signal input
rlabel metal2 s 1582 0 1638 160 6 N2MID[1]
port 218 nsew signal input
rlabel metal2 s 1858 0 1914 160 6 N2MID[2]
port 219 nsew signal input
rlabel metal2 s 2134 0 2190 160 6 N2MID[3]
port 220 nsew signal input
rlabel metal2 s 2410 0 2466 160 6 N2MID[4]
port 221 nsew signal input
rlabel metal2 s 2686 0 2742 160 6 N2MID[5]
port 222 nsew signal input
rlabel metal2 s 2962 0 3018 160 6 N2MID[6]
port 223 nsew signal input
rlabel metal2 s 3238 0 3294 160 6 N2MID[7]
port 224 nsew signal input
rlabel metal2 s 5722 44463 5778 44623 6 N4BEG[0]
port 225 nsew signal output
rlabel metal2 s 8482 44463 8538 44623 6 N4BEG[10]
port 226 nsew signal output
rlabel metal2 s 8758 44463 8814 44623 6 N4BEG[11]
port 227 nsew signal output
rlabel metal2 s 9034 44463 9090 44623 6 N4BEG[12]
port 228 nsew signal output
rlabel metal2 s 9310 44463 9366 44623 6 N4BEG[13]
port 229 nsew signal output
rlabel metal2 s 9586 44463 9642 44623 6 N4BEG[14]
port 230 nsew signal output
rlabel metal2 s 9862 44463 9918 44623 6 N4BEG[15]
port 231 nsew signal output
rlabel metal2 s 5998 44463 6054 44623 6 N4BEG[1]
port 232 nsew signal output
rlabel metal2 s 6274 44463 6330 44623 6 N4BEG[2]
port 233 nsew signal output
rlabel metal2 s 6550 44463 6606 44623 6 N4BEG[3]
port 234 nsew signal output
rlabel metal2 s 6826 44463 6882 44623 6 N4BEG[4]
port 235 nsew signal output
rlabel metal2 s 7102 44463 7158 44623 6 N4BEG[5]
port 236 nsew signal output
rlabel metal2 s 7378 44463 7434 44623 6 N4BEG[6]
port 237 nsew signal output
rlabel metal2 s 7654 44463 7710 44623 6 N4BEG[7]
port 238 nsew signal output
rlabel metal2 s 7930 44463 7986 44623 6 N4BEG[8]
port 239 nsew signal output
rlabel metal2 s 8206 44463 8262 44623 6 N4BEG[9]
port 240 nsew signal output
rlabel metal2 s 5722 0 5778 160 6 N4END[0]
port 241 nsew signal input
rlabel metal2 s 8482 0 8538 160 6 N4END[10]
port 242 nsew signal input
rlabel metal2 s 8758 0 8814 160 6 N4END[11]
port 243 nsew signal input
rlabel metal2 s 9034 0 9090 160 6 N4END[12]
port 244 nsew signal input
rlabel metal2 s 9310 0 9366 160 6 N4END[13]
port 245 nsew signal input
rlabel metal2 s 9586 0 9642 160 6 N4END[14]
port 246 nsew signal input
rlabel metal2 s 9862 0 9918 160 6 N4END[15]
port 247 nsew signal input
rlabel metal2 s 5998 0 6054 160 6 N4END[1]
port 248 nsew signal input
rlabel metal2 s 6274 0 6330 160 6 N4END[2]
port 249 nsew signal input
rlabel metal2 s 6550 0 6606 160 6 N4END[3]
port 250 nsew signal input
rlabel metal2 s 6826 0 6882 160 6 N4END[4]
port 251 nsew signal input
rlabel metal2 s 7102 0 7158 160 6 N4END[5]
port 252 nsew signal input
rlabel metal2 s 7378 0 7434 160 6 N4END[6]
port 253 nsew signal input
rlabel metal2 s 7654 0 7710 160 6 N4END[7]
port 254 nsew signal input
rlabel metal2 s 7930 0 7986 160 6 N4END[8]
port 255 nsew signal input
rlabel metal2 s 8206 0 8262 160 6 N4END[9]
port 256 nsew signal input
rlabel metal3 s 25840 7080 26000 7200 6 RAM2FAB_D0_I0
port 257 nsew signal input
rlabel metal3 s 25840 7624 26000 7744 6 RAM2FAB_D0_I1
port 258 nsew signal input
rlabel metal3 s 25840 8168 26000 8288 6 RAM2FAB_D0_I2
port 259 nsew signal input
rlabel metal3 s 25840 8712 26000 8832 6 RAM2FAB_D0_I3
port 260 nsew signal input
rlabel metal3 s 25840 4904 26000 5024 6 RAM2FAB_D1_I0
port 261 nsew signal input
rlabel metal3 s 25840 5448 26000 5568 6 RAM2FAB_D1_I1
port 262 nsew signal input
rlabel metal3 s 25840 5992 26000 6112 6 RAM2FAB_D1_I2
port 263 nsew signal input
rlabel metal3 s 25840 6536 26000 6656 6 RAM2FAB_D1_I3
port 264 nsew signal input
rlabel metal3 s 25840 2728 26000 2848 6 RAM2FAB_D2_I0
port 265 nsew signal input
rlabel metal3 s 25840 3272 26000 3392 6 RAM2FAB_D2_I1
port 266 nsew signal input
rlabel metal3 s 25840 3816 26000 3936 6 RAM2FAB_D2_I2
port 267 nsew signal input
rlabel metal3 s 25840 4360 26000 4480 6 RAM2FAB_D2_I3
port 268 nsew signal input
rlabel metal3 s 25840 552 26000 672 6 RAM2FAB_D3_I0
port 269 nsew signal input
rlabel metal3 s 25840 1096 26000 1216 6 RAM2FAB_D3_I1
port 270 nsew signal input
rlabel metal3 s 25840 1640 26000 1760 6 RAM2FAB_D3_I2
port 271 nsew signal input
rlabel metal3 s 25840 2184 26000 2304 6 RAM2FAB_D3_I3
port 272 nsew signal input
rlabel metal2 s 10138 0 10194 160 6 S1BEG[0]
port 273 nsew signal output
rlabel metal2 s 10414 0 10470 160 6 S1BEG[1]
port 274 nsew signal output
rlabel metal2 s 10690 0 10746 160 6 S1BEG[2]
port 275 nsew signal output
rlabel metal2 s 10966 0 11022 160 6 S1BEG[3]
port 276 nsew signal output
rlabel metal2 s 10138 44463 10194 44623 6 S1END[0]
port 277 nsew signal input
rlabel metal2 s 10414 44463 10470 44623 6 S1END[1]
port 278 nsew signal input
rlabel metal2 s 10690 44463 10746 44623 6 S1END[2]
port 279 nsew signal input
rlabel metal2 s 10966 44463 11022 44623 6 S1END[3]
port 280 nsew signal input
rlabel metal2 s 13450 0 13506 160 6 S2BEG[0]
port 281 nsew signal output
rlabel metal2 s 13726 0 13782 160 6 S2BEG[1]
port 282 nsew signal output
rlabel metal2 s 14002 0 14058 160 6 S2BEG[2]
port 283 nsew signal output
rlabel metal2 s 14278 0 14334 160 6 S2BEG[3]
port 284 nsew signal output
rlabel metal2 s 14554 0 14610 160 6 S2BEG[4]
port 285 nsew signal output
rlabel metal2 s 14830 0 14886 160 6 S2BEG[5]
port 286 nsew signal output
rlabel metal2 s 15106 0 15162 160 6 S2BEG[6]
port 287 nsew signal output
rlabel metal2 s 15382 0 15438 160 6 S2BEG[7]
port 288 nsew signal output
rlabel metal2 s 11242 0 11298 160 6 S2BEGb[0]
port 289 nsew signal output
rlabel metal2 s 11518 0 11574 160 6 S2BEGb[1]
port 290 nsew signal output
rlabel metal2 s 11794 0 11850 160 6 S2BEGb[2]
port 291 nsew signal output
rlabel metal2 s 12070 0 12126 160 6 S2BEGb[3]
port 292 nsew signal output
rlabel metal2 s 12346 0 12402 160 6 S2BEGb[4]
port 293 nsew signal output
rlabel metal2 s 12622 0 12678 160 6 S2BEGb[5]
port 294 nsew signal output
rlabel metal2 s 12898 0 12954 160 6 S2BEGb[6]
port 295 nsew signal output
rlabel metal2 s 13174 0 13230 160 6 S2BEGb[7]
port 296 nsew signal output
rlabel metal2 s 11242 44463 11298 44623 6 S2END[0]
port 297 nsew signal input
rlabel metal2 s 11518 44463 11574 44623 6 S2END[1]
port 298 nsew signal input
rlabel metal2 s 11794 44463 11850 44623 6 S2END[2]
port 299 nsew signal input
rlabel metal2 s 12070 44463 12126 44623 6 S2END[3]
port 300 nsew signal input
rlabel metal2 s 12346 44463 12402 44623 6 S2END[4]
port 301 nsew signal input
rlabel metal2 s 12622 44463 12678 44623 6 S2END[5]
port 302 nsew signal input
rlabel metal2 s 12898 44463 12954 44623 6 S2END[6]
port 303 nsew signal input
rlabel metal2 s 13174 44463 13230 44623 6 S2END[7]
port 304 nsew signal input
rlabel metal2 s 13450 44463 13506 44623 6 S2MID[0]
port 305 nsew signal input
rlabel metal2 s 13726 44463 13782 44623 6 S2MID[1]
port 306 nsew signal input
rlabel metal2 s 14002 44463 14058 44623 6 S2MID[2]
port 307 nsew signal input
rlabel metal2 s 14278 44463 14334 44623 6 S2MID[3]
port 308 nsew signal input
rlabel metal2 s 14554 44463 14610 44623 6 S2MID[4]
port 309 nsew signal input
rlabel metal2 s 14830 44463 14886 44623 6 S2MID[5]
port 310 nsew signal input
rlabel metal2 s 15106 44463 15162 44623 6 S2MID[6]
port 311 nsew signal input
rlabel metal2 s 15382 44463 15438 44623 6 S2MID[7]
port 312 nsew signal input
rlabel metal2 s 15658 0 15714 160 6 S4BEG[0]
port 313 nsew signal output
rlabel metal2 s 18418 0 18474 160 6 S4BEG[10]
port 314 nsew signal output
rlabel metal2 s 18694 0 18750 160 6 S4BEG[11]
port 315 nsew signal output
rlabel metal2 s 18970 0 19026 160 6 S4BEG[12]
port 316 nsew signal output
rlabel metal2 s 19246 0 19302 160 6 S4BEG[13]
port 317 nsew signal output
rlabel metal2 s 19522 0 19578 160 6 S4BEG[14]
port 318 nsew signal output
rlabel metal2 s 19798 0 19854 160 6 S4BEG[15]
port 319 nsew signal output
rlabel metal2 s 15934 0 15990 160 6 S4BEG[1]
port 320 nsew signal output
rlabel metal2 s 16210 0 16266 160 6 S4BEG[2]
port 321 nsew signal output
rlabel metal2 s 16486 0 16542 160 6 S4BEG[3]
port 322 nsew signal output
rlabel metal2 s 16762 0 16818 160 6 S4BEG[4]
port 323 nsew signal output
rlabel metal2 s 17038 0 17094 160 6 S4BEG[5]
port 324 nsew signal output
rlabel metal2 s 17314 0 17370 160 6 S4BEG[6]
port 325 nsew signal output
rlabel metal2 s 17590 0 17646 160 6 S4BEG[7]
port 326 nsew signal output
rlabel metal2 s 17866 0 17922 160 6 S4BEG[8]
port 327 nsew signal output
rlabel metal2 s 18142 0 18198 160 6 S4BEG[9]
port 328 nsew signal output
rlabel metal2 s 15658 44463 15714 44623 6 S4END[0]
port 329 nsew signal input
rlabel metal2 s 18418 44463 18474 44623 6 S4END[10]
port 330 nsew signal input
rlabel metal2 s 18694 44463 18750 44623 6 S4END[11]
port 331 nsew signal input
rlabel metal2 s 18970 44463 19026 44623 6 S4END[12]
port 332 nsew signal input
rlabel metal2 s 19246 44463 19302 44623 6 S4END[13]
port 333 nsew signal input
rlabel metal2 s 19522 44463 19578 44623 6 S4END[14]
port 334 nsew signal input
rlabel metal2 s 19798 44463 19854 44623 6 S4END[15]
port 335 nsew signal input
rlabel metal2 s 15934 44463 15990 44623 6 S4END[1]
port 336 nsew signal input
rlabel metal2 s 16210 44463 16266 44623 6 S4END[2]
port 337 nsew signal input
rlabel metal2 s 16486 44463 16542 44623 6 S4END[3]
port 338 nsew signal input
rlabel metal2 s 16762 44463 16818 44623 6 S4END[4]
port 339 nsew signal input
rlabel metal2 s 17038 44463 17094 44623 6 S4END[5]
port 340 nsew signal input
rlabel metal2 s 17314 44463 17370 44623 6 S4END[6]
port 341 nsew signal input
rlabel metal2 s 17590 44463 17646 44623 6 S4END[7]
port 342 nsew signal input
rlabel metal2 s 17866 44463 17922 44623 6 S4END[8]
port 343 nsew signal input
rlabel metal2 s 18142 44463 18198 44623 6 S4END[9]
port 344 nsew signal input
rlabel metal2 s 20074 0 20130 160 6 UserCLK
port 345 nsew signal input
rlabel metal2 s 20074 44463 20130 44623 6 UserCLKo
port 346 nsew signal output
rlabel metal4 s 6878 1040 7198 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 12812 1040 13132 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 18746 1040 19066 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 24680 1040 25000 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 3911 1040 4231 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 9845 1040 10165 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 15779 1040 16099 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 21713 1040 22033 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal3 s 0 4904 160 5024 6 W1BEG[0]
port 349 nsew signal output
rlabel metal3 s 0 5176 160 5296 6 W1BEG[1]
port 350 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 W1BEG[2]
port 351 nsew signal output
rlabel metal3 s 0 5720 160 5840 6 W1BEG[3]
port 352 nsew signal output
rlabel metal3 s 0 5992 160 6112 6 W2BEG[0]
port 353 nsew signal output
rlabel metal3 s 0 6264 160 6384 6 W2BEG[1]
port 354 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 W2BEG[2]
port 355 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 W2BEG[3]
port 356 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 W2BEG[4]
port 357 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 W2BEG[5]
port 358 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 W2BEG[6]
port 359 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 W2BEG[7]
port 360 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 W2BEGb[0]
port 361 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 W2BEGb[1]
port 362 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 W2BEGb[2]
port 363 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 W2BEGb[3]
port 364 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 W2BEGb[4]
port 365 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 W2BEGb[5]
port 366 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 W2BEGb[6]
port 367 nsew signal output
rlabel metal3 s 0 10072 160 10192 6 W2BEGb[7]
port 368 nsew signal output
rlabel metal3 s 0 14696 160 14816 6 W6BEG[0]
port 369 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 W6BEG[10]
port 370 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 W6BEG[11]
port 371 nsew signal output
rlabel metal3 s 0 14968 160 15088 6 W6BEG[1]
port 372 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 W6BEG[2]
port 373 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 W6BEG[3]
port 374 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 W6BEG[4]
port 375 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 W6BEG[5]
port 376 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 W6BEG[6]
port 377 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 W6BEG[7]
port 378 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 W6BEG[8]
port 379 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 W6BEG[9]
port 380 nsew signal output
rlabel metal3 s 0 10344 160 10464 6 WW4BEG[0]
port 381 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 WW4BEG[10]
port 382 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 WW4BEG[11]
port 383 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 WW4BEG[12]
port 384 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 WW4BEG[13]
port 385 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 WW4BEG[14]
port 386 nsew signal output
rlabel metal3 s 0 14424 160 14544 6 WW4BEG[15]
port 387 nsew signal output
rlabel metal3 s 0 10616 160 10736 6 WW4BEG[1]
port 388 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 WW4BEG[2]
port 389 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 WW4BEG[3]
port 390 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 WW4BEG[4]
port 391 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 WW4BEG[5]
port 392 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 WW4BEG[6]
port 393 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 WW4BEG[7]
port 394 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 WW4BEG[8]
port 395 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 WW4BEG[9]
port 396 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 26000 44623
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4310154
string GDS_FILE /home/asma/Desktop/FPGA_IGNITE_2024/openlane/RAM_IO_redo/runs/24_11_24_22_44/results/signoff/RAM_IO.magic.gds
string GDS_START 173598
<< end >>

