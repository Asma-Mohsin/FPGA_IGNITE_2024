magic
tech sky130A
magscale 1 2
timestamp 1732405133
<< viali >>
rect 1869 7497 1903 7531
rect 2789 7497 2823 7531
rect 3341 7497 3375 7531
rect 4261 7497 4295 7531
rect 4813 7497 4847 7531
rect 5549 7497 5583 7531
rect 5917 7497 5951 7531
rect 7021 7497 7055 7531
rect 7389 7497 7423 7531
rect 8033 7497 8067 7531
rect 9229 7497 9263 7531
rect 9965 7497 9999 7531
rect 10517 7497 10551 7531
rect 11069 7497 11103 7531
rect 12173 7497 12207 7531
rect 12909 7497 12943 7531
rect 13829 7497 13863 7531
rect 14381 7497 14415 7531
rect 15301 7497 15335 7531
rect 15853 7497 15887 7531
rect 16313 7497 16347 7531
rect 16865 7497 16899 7531
rect 19349 7497 19383 7531
rect 19809 7497 19843 7531
rect 22753 7497 22787 7531
rect 23489 7497 23523 7531
rect 24961 7497 24995 7531
rect 25697 7497 25731 7531
rect 26249 7497 26283 7531
rect 28181 7497 28215 7531
rect 28917 7497 28951 7531
rect 31309 7497 31343 7531
rect 32321 7497 32355 7531
rect 32873 7497 32907 7531
rect 33517 7497 33551 7531
rect 34253 7497 34287 7531
rect 34989 7497 35023 7531
rect 35909 7497 35943 7531
rect 36461 7497 36495 7531
rect 36829 7497 36863 7531
rect 37473 7497 37507 7531
rect 38025 7497 38059 7531
rect 38669 7497 38703 7531
rect 39405 7497 39439 7531
rect 40141 7497 40175 7531
rect 40877 7497 40911 7531
rect 41613 7497 41647 7531
rect 42625 7497 42659 7531
rect 43177 7497 43211 7531
rect 43821 7497 43855 7531
rect 5273 7429 5307 7463
rect 8309 7429 8343 7463
rect 8677 7429 8711 7463
rect 32229 7429 32263 7463
rect 36369 7429 36403 7463
rect 40785 7429 40819 7463
rect 43085 7429 43119 7463
rect 1777 7361 1811 7395
rect 2513 7361 2547 7395
rect 3249 7361 3283 7395
rect 3985 7361 4019 7395
rect 4721 7361 4755 7395
rect 5825 7361 5859 7395
rect 6745 7361 6779 7395
rect 7297 7361 7331 7395
rect 9137 7361 9171 7395
rect 9873 7361 9907 7395
rect 10425 7361 10459 7395
rect 10977 7361 11011 7395
rect 12081 7361 12115 7395
rect 12817 7361 12851 7395
rect 13553 7361 13587 7395
rect 14289 7361 14323 7395
rect 15025 7361 15059 7395
rect 15761 7361 15795 7395
rect 16497 7361 16531 7395
rect 16681 7361 16715 7395
rect 17325 7361 17359 7395
rect 17877 7361 17911 7395
rect 18797 7361 18831 7395
rect 19533 7361 19567 7395
rect 19625 7361 19659 7395
rect 20269 7361 20303 7395
rect 20361 7361 20395 7395
rect 21005 7361 21039 7395
rect 22017 7361 22051 7395
rect 22477 7361 22511 7395
rect 22569 7361 22603 7395
rect 23213 7361 23247 7395
rect 23305 7361 23339 7395
rect 23949 7361 23983 7395
rect 24685 7361 24719 7395
rect 24777 7361 24811 7395
rect 25421 7361 25455 7395
rect 25605 7361 25639 7395
rect 26157 7361 26191 7395
rect 26433 7361 26467 7395
rect 27169 7361 27203 7395
rect 27629 7361 27663 7395
rect 28365 7361 28399 7395
rect 28641 7361 28675 7395
rect 29101 7361 29135 7395
rect 29837 7361 29871 7395
rect 30573 7361 30607 7395
rect 31217 7361 31251 7395
rect 32781 7361 32815 7395
rect 33425 7361 33459 7395
rect 34161 7361 34195 7395
rect 34897 7361 34931 7395
rect 35633 7361 35667 7395
rect 37013 7361 37047 7395
rect 37381 7361 37415 7395
rect 37933 7361 37967 7395
rect 38577 7361 38611 7395
rect 39313 7361 39347 7395
rect 40049 7361 40083 7395
rect 41521 7361 41555 7395
rect 42533 7361 42567 7395
rect 43729 7361 43763 7395
rect 18613 7225 18647 7259
rect 20545 7225 20579 7259
rect 21833 7225 21867 7259
rect 23029 7225 23063 7259
rect 25237 7225 25271 7259
rect 25973 7225 26007 7259
rect 17141 7157 17175 7191
rect 18061 7157 18095 7191
rect 20085 7157 20119 7191
rect 20821 7157 20855 7191
rect 22293 7157 22327 7191
rect 23765 7157 23799 7191
rect 24501 7157 24535 7191
rect 26985 7157 27019 7191
rect 27445 7157 27479 7191
rect 28457 7157 28491 7191
rect 29653 7157 29687 7191
rect 30389 7157 30423 7191
rect 33793 6953 33827 6987
rect 34713 6953 34747 6987
rect 35265 6953 35299 6987
rect 37105 6953 37139 6987
rect 37841 6953 37875 6987
rect 38577 6953 38611 6987
rect 44281 6953 44315 6987
rect 1777 6817 1811 6851
rect 43913 6817 43947 6851
rect 33977 6749 34011 6783
rect 34897 6749 34931 6783
rect 35449 6725 35483 6759
rect 36553 6749 36587 6783
rect 37289 6749 37323 6783
rect 38025 6749 38059 6783
rect 38761 6749 38795 6783
rect 44189 6749 44223 6783
rect 1501 6681 1535 6715
rect 43637 6681 43671 6715
rect 36369 6613 36403 6647
rect 18981 4097 19015 4131
rect 19257 4097 19291 4131
rect 21373 4097 21407 4131
rect 21649 4097 21683 4131
rect 22017 4097 22051 4131
rect 26341 4097 26375 4131
rect 26801 4097 26835 4131
rect 32689 4097 32723 4131
rect 19073 3961 19107 3995
rect 26525 3961 26559 3995
rect 18797 3893 18831 3927
rect 21189 3893 21223 3927
rect 21465 3893 21499 3927
rect 21833 3893 21867 3927
rect 26617 3893 26651 3927
rect 32505 3893 32539 3927
rect 18705 3689 18739 3723
rect 19257 3689 19291 3723
rect 20269 3689 20303 3723
rect 21005 3689 21039 3723
rect 21649 3689 21683 3723
rect 29837 3689 29871 3723
rect 30849 3689 30883 3723
rect 33057 3689 33091 3723
rect 16773 3621 16807 3655
rect 16865 3621 16899 3655
rect 17325 3621 17359 3655
rect 23029 3621 23063 3655
rect 23765 3621 23799 3655
rect 23857 3621 23891 3655
rect 25881 3621 25915 3655
rect 26617 3621 26651 3655
rect 26985 3621 27019 3655
rect 27353 3621 27387 3655
rect 27445 3621 27479 3655
rect 28365 3621 28399 3655
rect 31585 3621 31619 3655
rect 16589 3485 16623 3519
rect 17049 3485 17083 3519
rect 17141 3485 17175 3519
rect 17417 3485 17451 3519
rect 17877 3485 17911 3519
rect 18153 3485 18187 3519
rect 18429 3485 18463 3519
rect 18521 3485 18555 3519
rect 19073 3485 19107 3519
rect 19441 3485 19475 3519
rect 19717 3485 19751 3519
rect 19993 3485 20027 3519
rect 20085 3485 20119 3519
rect 20545 3485 20579 3519
rect 20821 3485 20855 3519
rect 21281 3485 21315 3519
rect 21465 3485 21499 3519
rect 21925 3485 21959 3519
rect 22201 3485 22235 3519
rect 22477 3485 22511 3519
rect 22569 3485 22603 3519
rect 23213 3485 23247 3519
rect 23489 3485 23523 3519
rect 23581 3485 23615 3519
rect 24041 3485 24075 3519
rect 24685 3485 24719 3519
rect 24961 3485 24995 3519
rect 25237 3485 25271 3519
rect 25513 3485 25547 3519
rect 25697 3485 25731 3519
rect 26157 3485 26191 3519
rect 27169 3485 27203 3519
rect 27629 3485 27663 3519
rect 27905 3485 27939 3519
rect 28549 3485 28583 3519
rect 28825 3485 28859 3519
rect 29101 3485 29135 3519
rect 29377 3485 29411 3519
rect 30205 3485 30239 3519
rect 30481 3485 30515 3519
rect 30757 3485 30791 3519
rect 31217 3485 31251 3519
rect 31493 3485 31527 3519
rect 31769 3485 31803 3519
rect 32045 3485 32079 3519
rect 32321 3485 32355 3519
rect 32597 3485 32631 3519
rect 26433 3417 26467 3451
rect 26801 3417 26835 3451
rect 28089 3417 28123 3451
rect 29745 3417 29779 3451
rect 32965 3417 32999 3451
rect 17601 3349 17635 3383
rect 17693 3349 17727 3383
rect 17969 3349 18003 3383
rect 18245 3349 18279 3383
rect 18889 3349 18923 3383
rect 19533 3349 19567 3383
rect 19809 3349 19843 3383
rect 20361 3349 20395 3383
rect 21097 3349 21131 3383
rect 21741 3349 21775 3383
rect 22017 3349 22051 3383
rect 22293 3349 22327 3383
rect 22753 3349 22787 3383
rect 23305 3349 23339 3383
rect 24501 3349 24535 3383
rect 24777 3349 24811 3383
rect 25053 3349 25087 3383
rect 25329 3349 25363 3383
rect 25973 3349 26007 3383
rect 27721 3349 27755 3383
rect 28181 3349 28215 3383
rect 28641 3349 28675 3383
rect 28917 3349 28951 3383
rect 29193 3349 29227 3383
rect 30021 3349 30055 3383
rect 30297 3349 30331 3383
rect 31033 3349 31067 3383
rect 31309 3349 31343 3383
rect 31861 3349 31895 3383
rect 32137 3349 32171 3383
rect 32413 3349 32447 3383
rect 13737 3145 13771 3179
rect 14565 3145 14599 3179
rect 17233 3145 17267 3179
rect 17325 3145 17359 3179
rect 18153 3145 18187 3179
rect 24041 3145 24075 3179
rect 28273 3145 28307 3179
rect 30481 3145 30515 3179
rect 34529 3145 34563 3179
rect 35449 3145 35483 3179
rect 39129 3145 39163 3179
rect 17695 3077 17729 3111
rect 18061 3077 18095 3111
rect 18797 3077 18831 3111
rect 19717 3077 19751 3111
rect 20177 3077 20211 3111
rect 22753 3077 22787 3111
rect 23305 3077 23339 3111
rect 25237 3077 25271 3111
rect 25789 3077 25823 3111
rect 26341 3077 26375 3111
rect 27077 3077 27111 3111
rect 27629 3077 27663 3111
rect 29837 3077 29871 3111
rect 30389 3077 30423 3111
rect 32229 3077 32263 3111
rect 32781 3077 32815 3111
rect 34437 3077 34471 3111
rect 9137 3009 9171 3043
rect 13553 3009 13587 3043
rect 14381 3009 14415 3043
rect 15945 3009 15979 3043
rect 16957 3009 16991 3043
rect 17049 3009 17083 3043
rect 17509 3009 17543 3043
rect 18429 3009 18463 3043
rect 19165 3009 19199 3043
rect 20729 3009 20763 3043
rect 21281 3009 21315 3043
rect 22017 3009 22051 3043
rect 22201 3009 22235 3043
rect 23949 3009 23983 3043
rect 24225 3009 24259 3043
rect 24501 3009 24535 3043
rect 24685 3009 24719 3043
rect 28181 3009 28215 3043
rect 28733 3009 28767 3043
rect 29285 3009 29319 3043
rect 30941 3009 30975 3043
rect 31493 3009 31527 3043
rect 33333 3009 33367 3043
rect 33885 3009 33919 3043
rect 34989 3009 35023 3043
rect 35633 3009 35667 3043
rect 38945 3009 38979 3043
rect 15669 2941 15703 2975
rect 19349 2941 19383 2975
rect 19901 2941 19935 2975
rect 9321 2873 9355 2907
rect 23765 2873 23799 2907
rect 32965 2873 32999 2907
rect 16773 2805 16807 2839
rect 17785 2805 17819 2839
rect 18521 2805 18555 2839
rect 18889 2805 18923 2839
rect 20269 2805 20303 2839
rect 20821 2805 20855 2839
rect 21373 2805 21407 2839
rect 21833 2805 21867 2839
rect 22293 2805 22327 2839
rect 22845 2805 22879 2839
rect 23397 2805 23431 2839
rect 24317 2805 24351 2839
rect 24777 2805 24811 2839
rect 25329 2805 25363 2839
rect 25881 2805 25915 2839
rect 26433 2805 26467 2839
rect 27169 2805 27203 2839
rect 27721 2805 27755 2839
rect 28825 2805 28859 2839
rect 29377 2805 29411 2839
rect 29929 2805 29963 2839
rect 31033 2805 31067 2839
rect 31585 2805 31619 2839
rect 32321 2805 32355 2839
rect 33425 2805 33459 2839
rect 33977 2805 34011 2839
rect 35081 2805 35115 2839
rect 6561 2601 6595 2635
rect 9689 2601 9723 2635
rect 9965 2601 9999 2635
rect 13185 2601 13219 2635
rect 15117 2601 15151 2635
rect 15393 2601 15427 2635
rect 18337 2601 18371 2635
rect 18889 2601 18923 2635
rect 25145 2601 25179 2635
rect 26249 2601 26283 2635
rect 26801 2601 26835 2635
rect 27721 2601 27755 2635
rect 29745 2601 29779 2635
rect 30849 2601 30883 2635
rect 32321 2601 32355 2635
rect 34897 2601 34931 2635
rect 36093 2601 36127 2635
rect 36645 2601 36679 2635
rect 37105 2601 37139 2635
rect 37473 2601 37507 2635
rect 38025 2601 38059 2635
rect 39129 2601 39163 2635
rect 5917 2533 5951 2567
rect 7113 2533 7147 2567
rect 10333 2533 10367 2567
rect 11069 2533 11103 2567
rect 11345 2533 11379 2567
rect 11989 2533 12023 2567
rect 12265 2533 12299 2567
rect 14565 2533 14599 2567
rect 30389 2533 30423 2567
rect 31769 2533 31803 2567
rect 34345 2533 34379 2567
rect 36001 2533 36035 2567
rect 38301 2533 38335 2567
rect 15945 2465 15979 2499
rect 16957 2465 16991 2499
rect 17969 2465 18003 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 29009 2465 29043 2499
rect 33609 2465 33643 2499
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7205 2397 7239 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 8033 2397 8067 2431
rect 8309 2397 8343 2431
rect 8585 2397 8619 2431
rect 8953 2397 8987 2431
rect 9229 2397 9263 2431
rect 9505 2397 9539 2431
rect 9781 2397 9815 2431
rect 10057 2397 10091 2431
rect 10517 2397 10551 2431
rect 10793 2397 10827 2431
rect 10885 2397 10919 2431
rect 11161 2397 11195 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 12081 2397 12115 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 13369 2397 13403 2431
rect 13461 2397 13495 2431
rect 13737 2397 13771 2431
rect 14473 2397 14507 2431
rect 14749 2397 14783 2431
rect 15025 2397 15059 2431
rect 15301 2397 15335 2431
rect 15577 2397 15611 2431
rect 15669 2397 15703 2431
rect 16681 2397 16715 2431
rect 17785 2397 17819 2431
rect 18245 2397 18279 2431
rect 18521 2397 18555 2431
rect 18797 2397 18831 2431
rect 19073 2397 19107 2431
rect 19441 2397 19475 2431
rect 19625 2397 19659 2431
rect 21281 2397 21315 2431
rect 22017 2397 22051 2431
rect 22201 2397 22235 2431
rect 23305 2397 23339 2431
rect 23857 2397 23891 2431
rect 25053 2397 25087 2431
rect 25605 2397 25639 2431
rect 26617 2397 26651 2431
rect 27629 2397 27663 2431
rect 28181 2397 28215 2431
rect 28733 2397 28767 2431
rect 29377 2397 29411 2431
rect 29653 2397 29687 2431
rect 30757 2397 30791 2431
rect 31953 2397 31987 2431
rect 32781 2397 32815 2431
rect 33333 2397 33367 2431
rect 34529 2397 34563 2431
rect 35817 2397 35851 2431
rect 36277 2397 36311 2431
rect 36369 2397 36403 2431
rect 36829 2397 36863 2431
rect 36921 2397 36955 2431
rect 37289 2397 37323 2431
rect 37565 2397 37599 2431
rect 37841 2397 37875 2431
rect 38117 2397 38151 2431
rect 38393 2397 38427 2431
rect 38669 2397 38703 2431
rect 38945 2397 38979 2431
rect 39221 2397 39255 2431
rect 39497 2397 39531 2431
rect 39865 2397 39899 2431
rect 40141 2397 40175 2431
rect 40417 2397 40451 2431
rect 40693 2397 40727 2431
rect 40969 2397 41003 2431
rect 20177 2329 20211 2363
rect 20729 2329 20763 2363
rect 21097 2329 21131 2363
rect 21649 2329 21683 2363
rect 22569 2329 22603 2363
rect 22753 2329 22787 2363
rect 24501 2329 24535 2363
rect 26157 2329 26191 2363
rect 27077 2329 27111 2363
rect 30205 2329 30239 2363
rect 31309 2329 31343 2363
rect 32229 2329 32263 2363
rect 33885 2329 33919 2363
rect 34805 2329 34839 2363
rect 35357 2329 35391 2363
rect 5641 2261 5675 2295
rect 6193 2261 6227 2295
rect 6837 2261 6871 2295
rect 7389 2261 7423 2295
rect 7665 2261 7699 2295
rect 7941 2261 7975 2295
rect 8217 2261 8251 2295
rect 8493 2261 8527 2295
rect 8769 2261 8803 2295
rect 9137 2261 9171 2295
rect 9413 2261 9447 2295
rect 10241 2261 10275 2295
rect 10609 2261 10643 2295
rect 11713 2261 11747 2295
rect 12541 2261 12575 2295
rect 12817 2261 12851 2295
rect 13093 2261 13127 2295
rect 13645 2261 13679 2295
rect 13921 2261 13955 2295
rect 14289 2261 14323 2295
rect 14841 2261 14875 2295
rect 18061 2261 18095 2295
rect 18613 2261 18647 2295
rect 19257 2261 19291 2295
rect 21833 2261 21867 2295
rect 22845 2261 22879 2295
rect 23581 2261 23615 2295
rect 23949 2261 23983 2295
rect 24593 2261 24627 2295
rect 25697 2261 25731 2295
rect 27169 2261 27203 2295
rect 28273 2261 28307 2295
rect 29193 2261 29227 2295
rect 31401 2261 31435 2295
rect 32873 2261 32907 2295
rect 33977 2261 34011 2295
rect 35449 2261 35483 2295
rect 36553 2261 36587 2295
rect 37749 2261 37783 2295
rect 38577 2261 38611 2295
rect 38853 2261 38887 2295
rect 39405 2261 39439 2295
rect 39681 2261 39715 2295
rect 40049 2261 40083 2295
rect 40325 2261 40359 2295
rect 40601 2261 40635 2295
rect 40877 2261 40911 2295
rect 41153 2261 41187 2295
<< metal1 >>
rect 20530 8168 20536 8220
rect 20588 8208 20594 8220
rect 30742 8208 30748 8220
rect 20588 8180 30748 8208
rect 20588 8168 20594 8180
rect 30742 8168 30748 8180
rect 30800 8168 30806 8220
rect 18322 8100 18328 8152
rect 18380 8140 18386 8152
rect 18380 8112 31754 8140
rect 18380 8100 18386 8112
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 20990 8072 20996 8084
rect 10836 8044 20996 8072
rect 10836 8032 10842 8044
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 23474 8004 23480 8016
rect 9876 7976 23480 8004
rect 9876 7744 9904 7976
rect 23474 7964 23480 7976
rect 23532 7964 23538 8016
rect 19518 7896 19524 7948
rect 19576 7936 19582 7948
rect 19576 7908 31524 7936
rect 19576 7896 19582 7908
rect 31496 7880 31524 7908
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 25682 7868 25688 7880
rect 17276 7840 25688 7868
rect 17276 7828 17282 7840
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 31478 7828 31484 7880
rect 31536 7828 31542 7880
rect 31726 7868 31754 8112
rect 42702 7868 42708 7880
rect 31726 7840 42708 7868
rect 42702 7828 42708 7840
rect 42760 7828 42766 7880
rect 19794 7760 19800 7812
rect 19852 7800 19858 7812
rect 36906 7800 36912 7812
rect 19852 7772 36912 7800
rect 19852 7760 19858 7772
rect 36906 7760 36912 7772
rect 36964 7760 36970 7812
rect 9858 7692 9864 7744
rect 9916 7692 9922 7744
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 29270 7732 29276 7744
rect 18656 7704 29276 7732
rect 18656 7692 18662 7704
rect 29270 7692 29276 7704
rect 29328 7692 29334 7744
rect 1104 7642 45051 7664
rect 1104 7590 11896 7642
rect 11948 7590 11960 7642
rect 12012 7590 12024 7642
rect 12076 7590 12088 7642
rect 12140 7590 12152 7642
rect 12204 7590 22843 7642
rect 22895 7590 22907 7642
rect 22959 7590 22971 7642
rect 23023 7590 23035 7642
rect 23087 7590 23099 7642
rect 23151 7590 33790 7642
rect 33842 7590 33854 7642
rect 33906 7590 33918 7642
rect 33970 7590 33982 7642
rect 34034 7590 34046 7642
rect 34098 7590 44737 7642
rect 44789 7590 44801 7642
rect 44853 7590 44865 7642
rect 44917 7590 44929 7642
rect 44981 7590 44993 7642
rect 45045 7590 45051 7642
rect 1104 7568 45051 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 1857 7531 1915 7537
rect 1857 7528 1869 7531
rect 1636 7500 1869 7528
rect 1636 7488 1642 7500
rect 1857 7497 1869 7500
rect 1903 7497 1915 7531
rect 1857 7491 1915 7497
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 3108 7500 3341 7528
rect 3108 7488 3114 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 3970 7488 3976 7540
rect 4028 7528 4034 7540
rect 4249 7531 4307 7537
rect 4249 7528 4261 7531
rect 4028 7500 4261 7528
rect 4028 7488 4034 7500
rect 4249 7497 4261 7500
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4580 7500 4813 7528
rect 4580 7488 4586 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 5534 7488 5540 7540
rect 5592 7488 5598 7540
rect 5902 7488 5908 7540
rect 5960 7488 5966 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 7009 7531 7067 7537
rect 7009 7528 7021 7531
rect 6880 7500 7021 7528
rect 6880 7488 6886 7500
rect 7009 7497 7021 7500
rect 7055 7497 7067 7531
rect 7009 7491 7067 7497
rect 7374 7488 7380 7540
rect 7432 7488 7438 7540
rect 8021 7531 8079 7537
rect 8021 7497 8033 7531
rect 8067 7528 8079 7531
rect 8067 7500 8708 7528
rect 8067 7497 8079 7500
rect 8021 7491 8079 7497
rect 8680 7472 8708 7500
rect 8938 7488 8944 7540
rect 8996 7528 9002 7540
rect 9217 7531 9275 7537
rect 9217 7528 9229 7531
rect 8996 7500 9229 7528
rect 8996 7488 9002 7500
rect 9217 7497 9229 7500
rect 9263 7497 9275 7531
rect 9217 7491 9275 7497
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 9953 7531 10011 7537
rect 9953 7528 9965 7531
rect 9732 7500 9965 7528
rect 9732 7488 9738 7500
rect 9953 7497 9965 7500
rect 9999 7497 10011 7531
rect 9953 7491 10011 7497
rect 10502 7488 10508 7540
rect 10560 7488 10566 7540
rect 11054 7488 11060 7540
rect 11112 7488 11118 7540
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11940 7500 12173 7528
rect 11940 7488 11946 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12897 7531 12955 7537
rect 12897 7528 12909 7531
rect 12676 7500 12909 7528
rect 12676 7488 12682 7500
rect 12897 7497 12909 7500
rect 12943 7497 12955 7531
rect 12897 7491 12955 7497
rect 13814 7488 13820 7540
rect 13872 7488 13878 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 14369 7531 14427 7537
rect 14369 7528 14381 7531
rect 14148 7500 14381 7528
rect 14148 7488 14154 7500
rect 14369 7497 14381 7500
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 15010 7488 15016 7540
rect 15068 7528 15074 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15068 7500 15301 7528
rect 15068 7488 15074 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 15841 7531 15899 7537
rect 15841 7528 15853 7531
rect 15620 7500 15853 7528
rect 15620 7488 15626 7500
rect 15841 7497 15853 7500
rect 15887 7497 15899 7531
rect 15841 7491 15899 7497
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 16853 7531 16911 7537
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 19150 7528 19156 7540
rect 16899 7500 19156 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 5261 7463 5319 7469
rect 3252 7432 5028 7460
rect 1762 7352 1768 7404
rect 1820 7352 1826 7404
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 3142 7392 3148 7404
rect 2547 7364 3148 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3252 7401 3280 7432
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 4614 7392 4620 7404
rect 4019 7364 4620 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 4724 7188 4752 7355
rect 5000 7256 5028 7432
rect 5261 7429 5273 7463
rect 5307 7460 5319 7463
rect 5307 7432 8248 7460
rect 5307 7429 5319 7432
rect 5261 7423 5319 7429
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5828 7324 5856 7355
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 8220 7392 8248 7432
rect 8294 7420 8300 7472
rect 8352 7420 8358 7472
rect 8662 7460 8668 7472
rect 8623 7432 8668 7460
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 11698 7460 11704 7472
rect 8772 7432 11704 7460
rect 8772 7392 8800 7432
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 16316 7460 16344 7491
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19242 7488 19248 7540
rect 19300 7488 19306 7540
rect 19334 7488 19340 7540
rect 19392 7488 19398 7540
rect 19794 7488 19800 7540
rect 19852 7488 19858 7540
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 22741 7531 22799 7537
rect 22741 7528 22753 7531
rect 19944 7500 22753 7528
rect 19944 7488 19950 7500
rect 22741 7497 22753 7500
rect 22787 7497 22799 7531
rect 22741 7491 22799 7497
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 24946 7488 24952 7540
rect 25004 7488 25010 7540
rect 25682 7488 25688 7540
rect 25740 7488 25746 7540
rect 26237 7531 26295 7537
rect 26237 7497 26249 7531
rect 26283 7528 26295 7531
rect 27890 7528 27896 7540
rect 26283 7500 27896 7528
rect 26283 7497 26295 7500
rect 26237 7491 26295 7497
rect 27890 7488 27896 7500
rect 27948 7488 27954 7540
rect 28169 7531 28227 7537
rect 28169 7497 28181 7531
rect 28215 7497 28227 7531
rect 28169 7491 28227 7497
rect 28905 7531 28963 7537
rect 28905 7497 28917 7531
rect 28951 7497 28963 7531
rect 28905 7491 28963 7497
rect 29012 7500 30696 7528
rect 16316 7432 16712 7460
rect 8220 7364 8800 7392
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9858 7352 9864 7404
rect 9916 7352 9922 7404
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 10778 7392 10784 7404
rect 10459 7364 10784 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 13262 7392 13268 7404
rect 12851 7364 13268 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 10870 7324 10876 7336
rect 5828 7296 10876 7324
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 8294 7256 8300 7268
rect 5000 7228 8300 7256
rect 8294 7216 8300 7228
rect 8352 7216 8358 7268
rect 12084 7256 12112 7355
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 13170 7284 13176 7336
rect 13228 7324 13234 7336
rect 13556 7324 13584 7355
rect 14274 7352 14280 7404
rect 14332 7352 14338 7404
rect 14642 7352 14648 7404
rect 14700 7392 14706 7404
rect 15013 7395 15071 7401
rect 15013 7392 15025 7395
rect 14700 7364 15025 7392
rect 14700 7352 14706 7364
rect 15013 7361 15025 7364
rect 15059 7361 15071 7395
rect 15013 7355 15071 7361
rect 15102 7352 15108 7404
rect 15160 7392 15166 7404
rect 15749 7395 15807 7401
rect 15749 7392 15761 7395
rect 15160 7364 15761 7392
rect 15160 7352 15166 7364
rect 15749 7361 15761 7364
rect 15795 7361 15807 7395
rect 15749 7355 15807 7361
rect 16482 7352 16488 7404
rect 16540 7352 16546 7404
rect 16684 7401 16712 7432
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 17092 7364 17325 7392
rect 17092 7352 17098 7364
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17862 7352 17868 7404
rect 17920 7352 17926 7404
rect 18506 7352 18512 7404
rect 18564 7392 18570 7404
rect 18785 7395 18843 7401
rect 18785 7392 18797 7395
rect 18564 7364 18797 7392
rect 18564 7352 18570 7364
rect 18785 7361 18797 7364
rect 18831 7361 18843 7395
rect 19260 7392 19288 7488
rect 20456 7432 26464 7460
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19260 7364 19533 7392
rect 18785 7355 18843 7361
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 13228 7296 13584 7324
rect 13228 7284 13234 7296
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 19628 7324 19656 7355
rect 19978 7352 19984 7404
rect 20036 7392 20042 7404
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 20036 7364 20269 7392
rect 20036 7352 20042 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7361 20407 7395
rect 20349 7355 20407 7361
rect 19116 7296 19656 7324
rect 19116 7284 19122 7296
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 20364 7324 20392 7355
rect 19852 7296 20392 7324
rect 19852 7284 19858 7296
rect 18601 7259 18659 7265
rect 12084 7228 18184 7256
rect 8386 7188 8392 7200
rect 4724 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 14458 7188 14464 7200
rect 8720 7160 14464 7188
rect 8720 7148 8726 7160
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 17126 7148 17132 7200
rect 17184 7148 17190 7200
rect 18046 7148 18052 7200
rect 18104 7148 18110 7200
rect 18156 7188 18184 7228
rect 18601 7225 18613 7259
rect 18647 7256 18659 7259
rect 20456 7256 20484 7432
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 20993 7395 21051 7401
rect 20993 7392 21005 7395
rect 20772 7364 21005 7392
rect 20772 7352 20778 7364
rect 20993 7361 21005 7364
rect 21039 7361 21051 7395
rect 20993 7355 21051 7361
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21508 7364 22017 7392
rect 21508 7352 21514 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22465 7395 22523 7401
rect 22465 7392 22477 7395
rect 22244 7364 22477 7392
rect 22244 7352 22250 7364
rect 22465 7361 22477 7364
rect 22511 7361 22523 7395
rect 22465 7355 22523 7361
rect 22554 7352 22560 7404
rect 22612 7352 22618 7404
rect 23198 7352 23204 7404
rect 23256 7352 23262 7404
rect 23290 7352 23296 7404
rect 23348 7352 23354 7404
rect 23658 7352 23664 7404
rect 23716 7392 23722 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23716 7364 23949 7392
rect 23716 7352 23722 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24394 7352 24400 7404
rect 24452 7392 24458 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24452 7364 24685 7392
rect 24452 7352 24458 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24765 7395 24823 7401
rect 24765 7361 24777 7395
rect 24811 7392 24823 7395
rect 25038 7392 25044 7404
rect 24811 7364 25044 7392
rect 24811 7361 24823 7364
rect 24765 7355 24823 7361
rect 25038 7352 25044 7364
rect 25096 7352 25102 7404
rect 25130 7352 25136 7404
rect 25188 7392 25194 7404
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 25188 7364 25421 7392
rect 25188 7352 25194 7364
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25409 7355 25467 7361
rect 25590 7352 25596 7404
rect 25648 7352 25654 7404
rect 25866 7352 25872 7404
rect 25924 7392 25930 7404
rect 26436 7401 26464 7432
rect 27798 7420 27804 7472
rect 27856 7460 27862 7472
rect 28184 7460 28212 7491
rect 27856 7432 28212 7460
rect 27856 7420 27862 7432
rect 26145 7395 26203 7401
rect 26145 7392 26157 7395
rect 25924 7364 26157 7392
rect 25924 7352 25930 7364
rect 26145 7361 26157 7364
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 26421 7395 26479 7401
rect 26421 7361 26433 7395
rect 26467 7361 26479 7395
rect 26421 7355 26479 7361
rect 26602 7352 26608 7404
rect 26660 7392 26666 7404
rect 27157 7395 27215 7401
rect 27157 7392 27169 7395
rect 26660 7364 27169 7392
rect 26660 7352 26666 7364
rect 27157 7361 27169 7364
rect 27203 7361 27215 7395
rect 27157 7355 27215 7361
rect 27338 7352 27344 7404
rect 27396 7392 27402 7404
rect 27617 7395 27675 7401
rect 27617 7392 27629 7395
rect 27396 7364 27629 7392
rect 27396 7352 27402 7364
rect 27617 7361 27629 7364
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 28074 7352 28080 7404
rect 28132 7392 28138 7404
rect 28353 7395 28411 7401
rect 28353 7392 28365 7395
rect 28132 7364 28365 7392
rect 28132 7352 28138 7364
rect 28353 7361 28365 7364
rect 28399 7361 28411 7395
rect 28353 7355 28411 7361
rect 28629 7395 28687 7401
rect 28629 7361 28641 7395
rect 28675 7392 28687 7395
rect 28920 7392 28948 7491
rect 29012 7472 29040 7500
rect 28994 7420 29000 7472
rect 29052 7420 29058 7472
rect 28675 7364 28948 7392
rect 28675 7361 28687 7364
rect 28629 7355 28687 7361
rect 29086 7352 29092 7404
rect 29144 7352 29150 7404
rect 29546 7352 29552 7404
rect 29604 7392 29610 7404
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 29604 7364 29837 7392
rect 29604 7352 29610 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 29825 7355 29883 7361
rect 30374 7352 30380 7404
rect 30432 7392 30438 7404
rect 30561 7395 30619 7401
rect 30561 7392 30573 7395
rect 30432 7364 30573 7392
rect 30432 7352 30438 7364
rect 30561 7361 30573 7364
rect 30607 7361 30619 7395
rect 30668 7392 30696 7500
rect 31018 7488 31024 7540
rect 31076 7528 31082 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 31076 7500 31309 7528
rect 31076 7488 31082 7500
rect 31297 7497 31309 7500
rect 31343 7497 31355 7531
rect 31297 7491 31355 7497
rect 31754 7488 31760 7540
rect 31812 7528 31818 7540
rect 32309 7531 32367 7537
rect 32309 7528 32321 7531
rect 31812 7500 32321 7528
rect 31812 7488 31818 7500
rect 32309 7497 32321 7500
rect 32355 7497 32367 7531
rect 32309 7491 32367 7497
rect 32490 7488 32496 7540
rect 32548 7528 32554 7540
rect 32861 7531 32919 7537
rect 32861 7528 32873 7531
rect 32548 7500 32873 7528
rect 32548 7488 32554 7500
rect 32861 7497 32873 7500
rect 32907 7497 32919 7531
rect 32861 7491 32919 7497
rect 33226 7488 33232 7540
rect 33284 7528 33290 7540
rect 33505 7531 33563 7537
rect 33505 7528 33517 7531
rect 33284 7500 33517 7528
rect 33284 7488 33290 7500
rect 33505 7497 33517 7500
rect 33551 7497 33563 7531
rect 33505 7491 33563 7497
rect 34238 7488 34244 7540
rect 34296 7488 34302 7540
rect 34698 7488 34704 7540
rect 34756 7528 34762 7540
rect 34977 7531 35035 7537
rect 34977 7528 34989 7531
rect 34756 7500 34989 7528
rect 34756 7488 34762 7500
rect 34977 7497 34989 7500
rect 35023 7497 35035 7531
rect 34977 7491 35035 7497
rect 35894 7488 35900 7540
rect 35952 7488 35958 7540
rect 36170 7488 36176 7540
rect 36228 7528 36234 7540
rect 36449 7531 36507 7537
rect 36449 7528 36461 7531
rect 36228 7500 36461 7528
rect 36228 7488 36234 7500
rect 36449 7497 36461 7500
rect 36495 7497 36507 7531
rect 36449 7491 36507 7497
rect 36817 7531 36875 7537
rect 36817 7497 36829 7531
rect 36863 7497 36875 7531
rect 36817 7491 36875 7497
rect 30742 7420 30748 7472
rect 30800 7460 30806 7472
rect 32217 7463 32275 7469
rect 32217 7460 32229 7463
rect 30800 7432 32229 7460
rect 30800 7420 30806 7432
rect 32217 7429 32229 7432
rect 32263 7429 32275 7463
rect 32217 7423 32275 7429
rect 36357 7463 36415 7469
rect 36357 7429 36369 7463
rect 36403 7460 36415 7463
rect 36832 7460 36860 7491
rect 36906 7488 36912 7540
rect 36964 7488 36970 7540
rect 37182 7488 37188 7540
rect 37240 7528 37246 7540
rect 37461 7531 37519 7537
rect 37461 7528 37473 7531
rect 37240 7500 37473 7528
rect 37240 7488 37246 7500
rect 37461 7497 37473 7500
rect 37507 7497 37519 7531
rect 37461 7491 37519 7497
rect 37642 7488 37648 7540
rect 37700 7528 37706 7540
rect 38013 7531 38071 7537
rect 38013 7528 38025 7531
rect 37700 7500 38025 7528
rect 37700 7488 37706 7500
rect 38013 7497 38025 7500
rect 38059 7497 38071 7531
rect 38013 7491 38071 7497
rect 38654 7488 38660 7540
rect 38712 7488 38718 7540
rect 39114 7488 39120 7540
rect 39172 7528 39178 7540
rect 39393 7531 39451 7537
rect 39393 7528 39405 7531
rect 39172 7500 39405 7528
rect 39172 7488 39178 7500
rect 39393 7497 39405 7500
rect 39439 7497 39451 7531
rect 39393 7491 39451 7497
rect 39850 7488 39856 7540
rect 39908 7528 39914 7540
rect 40129 7531 40187 7537
rect 40129 7528 40141 7531
rect 39908 7500 40141 7528
rect 39908 7488 39914 7500
rect 40129 7497 40141 7500
rect 40175 7497 40187 7531
rect 40129 7491 40187 7497
rect 40586 7488 40592 7540
rect 40644 7528 40650 7540
rect 40865 7531 40923 7537
rect 40865 7528 40877 7531
rect 40644 7500 40877 7528
rect 40644 7488 40650 7500
rect 40865 7497 40877 7500
rect 40911 7497 40923 7531
rect 40865 7491 40923 7497
rect 41322 7488 41328 7540
rect 41380 7528 41386 7540
rect 41601 7531 41659 7537
rect 41601 7528 41613 7531
rect 41380 7500 41613 7528
rect 41380 7488 41386 7500
rect 41601 7497 41613 7500
rect 41647 7497 41659 7531
rect 41601 7491 41659 7497
rect 42610 7488 42616 7540
rect 42668 7488 42674 7540
rect 42702 7488 42708 7540
rect 42760 7488 42766 7540
rect 42794 7488 42800 7540
rect 42852 7528 42858 7540
rect 43165 7531 43223 7537
rect 43165 7528 43177 7531
rect 42852 7500 43177 7528
rect 42852 7488 42858 7500
rect 43165 7497 43177 7500
rect 43211 7497 43223 7531
rect 43165 7491 43223 7497
rect 43530 7488 43536 7540
rect 43588 7528 43594 7540
rect 43809 7531 43867 7537
rect 43809 7528 43821 7531
rect 43588 7500 43821 7528
rect 43588 7488 43594 7500
rect 43809 7497 43821 7500
rect 43855 7497 43867 7531
rect 43809 7491 43867 7497
rect 36403 7432 36860 7460
rect 36924 7460 36952 7488
rect 40773 7463 40831 7469
rect 40773 7460 40785 7463
rect 36924 7432 40785 7460
rect 36403 7429 36415 7432
rect 36357 7423 36415 7429
rect 40773 7429 40785 7432
rect 40819 7429 40831 7463
rect 42720 7460 42748 7488
rect 43073 7463 43131 7469
rect 43073 7460 43085 7463
rect 40773 7423 40831 7429
rect 41386 7432 42564 7460
rect 42720 7432 43085 7460
rect 31205 7395 31263 7401
rect 31205 7392 31217 7395
rect 30668 7364 31217 7392
rect 30561 7355 30619 7361
rect 31205 7361 31217 7364
rect 31251 7361 31263 7395
rect 31205 7355 31263 7361
rect 32766 7352 32772 7404
rect 32824 7352 32830 7404
rect 33410 7352 33416 7404
rect 33468 7352 33474 7404
rect 34146 7352 34152 7404
rect 34204 7352 34210 7404
rect 34882 7352 34888 7404
rect 34940 7352 34946 7404
rect 35618 7352 35624 7404
rect 35676 7352 35682 7404
rect 35894 7352 35900 7404
rect 35952 7392 35958 7404
rect 36998 7392 37004 7404
rect 35952 7364 37004 7392
rect 35952 7352 35958 7364
rect 36998 7352 37004 7364
rect 37056 7352 37062 7404
rect 37366 7352 37372 7404
rect 37424 7352 37430 7404
rect 37458 7352 37464 7404
rect 37516 7392 37522 7404
rect 37921 7395 37979 7401
rect 37921 7392 37933 7395
rect 37516 7364 37933 7392
rect 37516 7352 37522 7364
rect 37921 7361 37933 7364
rect 37967 7361 37979 7395
rect 37921 7355 37979 7361
rect 38194 7352 38200 7404
rect 38252 7392 38258 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 38252 7364 38577 7392
rect 38252 7352 38258 7364
rect 38565 7361 38577 7364
rect 38611 7361 38623 7395
rect 38565 7355 38623 7361
rect 38930 7352 38936 7404
rect 38988 7392 38994 7404
rect 39301 7395 39359 7401
rect 39301 7392 39313 7395
rect 38988 7364 39313 7392
rect 38988 7352 38994 7364
rect 39301 7361 39313 7364
rect 39347 7361 39359 7395
rect 39301 7355 39359 7361
rect 39390 7352 39396 7404
rect 39448 7392 39454 7404
rect 40037 7395 40095 7401
rect 40037 7392 40049 7395
rect 39448 7364 40049 7392
rect 39448 7352 39454 7364
rect 40037 7361 40049 7364
rect 40083 7361 40095 7395
rect 40037 7355 40095 7361
rect 20548 7265 20576 7352
rect 29178 7324 29184 7336
rect 22066 7296 25176 7324
rect 18647 7228 20484 7256
rect 20533 7259 20591 7265
rect 18647 7225 18659 7228
rect 18601 7219 18659 7225
rect 20533 7225 20545 7259
rect 20579 7225 20591 7259
rect 20533 7219 20591 7225
rect 21821 7259 21879 7265
rect 21821 7225 21833 7259
rect 21867 7256 21879 7259
rect 22066 7256 22094 7296
rect 25148 7268 25176 7296
rect 25240 7296 29184 7324
rect 21867 7228 22094 7256
rect 23017 7259 23075 7265
rect 21867 7225 21879 7228
rect 21821 7219 21879 7225
rect 23017 7225 23029 7259
rect 23063 7256 23075 7259
rect 23566 7256 23572 7268
rect 23063 7228 23572 7256
rect 23063 7225 23075 7228
rect 23017 7219 23075 7225
rect 23566 7216 23572 7228
rect 23624 7216 23630 7268
rect 25130 7216 25136 7268
rect 25188 7216 25194 7268
rect 25240 7265 25268 7296
rect 29178 7284 29184 7296
rect 29236 7284 29242 7336
rect 29270 7284 29276 7336
rect 29328 7324 29334 7336
rect 41386 7324 41414 7432
rect 42536 7401 42564 7432
rect 43073 7429 43085 7432
rect 43119 7429 43131 7463
rect 43073 7423 43131 7429
rect 41509 7395 41567 7401
rect 41509 7361 41521 7395
rect 41555 7361 41567 7395
rect 41509 7355 41567 7361
rect 42521 7395 42579 7401
rect 42521 7361 42533 7395
rect 42567 7361 42579 7395
rect 42521 7355 42579 7361
rect 29328 7296 41414 7324
rect 29328 7284 29334 7296
rect 25225 7259 25283 7265
rect 25225 7225 25237 7259
rect 25271 7225 25283 7259
rect 25225 7219 25283 7225
rect 25961 7259 26019 7265
rect 25961 7225 25973 7259
rect 26007 7256 26019 7259
rect 28994 7256 29000 7268
rect 26007 7228 29000 7256
rect 26007 7225 26019 7228
rect 25961 7219 26019 7225
rect 28994 7216 29000 7228
rect 29052 7216 29058 7268
rect 30392 7228 31432 7256
rect 19886 7188 19892 7200
rect 18156 7160 19892 7188
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 20073 7191 20131 7197
rect 20073 7157 20085 7191
rect 20119 7188 20131 7191
rect 20346 7188 20352 7200
rect 20119 7160 20352 7188
rect 20119 7157 20131 7160
rect 20073 7151 20131 7157
rect 20346 7148 20352 7160
rect 20404 7148 20410 7200
rect 20809 7191 20867 7197
rect 20809 7157 20821 7191
rect 20855 7188 20867 7191
rect 21082 7188 21088 7200
rect 20855 7160 21088 7188
rect 20855 7157 20867 7160
rect 20809 7151 20867 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 22278 7148 22284 7200
rect 22336 7148 22342 7200
rect 23750 7148 23756 7200
rect 23808 7148 23814 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 24854 7188 24860 7200
rect 24535 7160 24860 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 24854 7148 24860 7160
rect 24912 7148 24918 7200
rect 26973 7191 27031 7197
rect 26973 7157 26985 7191
rect 27019 7188 27031 7191
rect 27338 7188 27344 7200
rect 27019 7160 27344 7188
rect 27019 7157 27031 7160
rect 26973 7151 27031 7157
rect 27338 7148 27344 7160
rect 27396 7148 27402 7200
rect 27433 7191 27491 7197
rect 27433 7157 27445 7191
rect 27479 7188 27491 7191
rect 28166 7188 28172 7200
rect 27479 7160 28172 7188
rect 27479 7157 27491 7160
rect 27433 7151 27491 7157
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 28445 7191 28503 7197
rect 28445 7157 28457 7191
rect 28491 7188 28503 7191
rect 28718 7188 28724 7200
rect 28491 7160 28724 7188
rect 28491 7157 28503 7160
rect 28445 7151 28503 7157
rect 28718 7148 28724 7160
rect 28776 7148 28782 7200
rect 29638 7148 29644 7200
rect 29696 7148 29702 7200
rect 30392 7197 30420 7228
rect 30377 7191 30435 7197
rect 30377 7157 30389 7191
rect 30423 7157 30435 7191
rect 31404 7188 31432 7228
rect 31478 7216 31484 7268
rect 31536 7256 31542 7268
rect 31536 7228 39344 7256
rect 31536 7216 31542 7228
rect 31938 7188 31944 7200
rect 31404 7160 31944 7188
rect 30377 7151 30435 7157
rect 31938 7148 31944 7160
rect 31996 7148 32002 7200
rect 33042 7148 33048 7200
rect 33100 7188 33106 7200
rect 39206 7188 39212 7200
rect 33100 7160 39212 7188
rect 33100 7148 33106 7160
rect 39206 7148 39212 7160
rect 39264 7148 39270 7200
rect 39316 7188 39344 7228
rect 41524 7188 41552 7355
rect 42610 7352 42616 7404
rect 42668 7392 42674 7404
rect 43717 7395 43775 7401
rect 43717 7392 43729 7395
rect 42668 7364 43729 7392
rect 42668 7352 42674 7364
rect 43717 7361 43729 7364
rect 43763 7361 43775 7395
rect 43717 7355 43775 7361
rect 39316 7160 41552 7188
rect 1104 7098 44896 7120
rect 1104 7046 6423 7098
rect 6475 7046 6487 7098
rect 6539 7046 6551 7098
rect 6603 7046 6615 7098
rect 6667 7046 6679 7098
rect 6731 7046 17370 7098
rect 17422 7046 17434 7098
rect 17486 7046 17498 7098
rect 17550 7046 17562 7098
rect 17614 7046 17626 7098
rect 17678 7046 28317 7098
rect 28369 7046 28381 7098
rect 28433 7046 28445 7098
rect 28497 7046 28509 7098
rect 28561 7046 28573 7098
rect 28625 7046 39264 7098
rect 39316 7046 39328 7098
rect 39380 7046 39392 7098
rect 39444 7046 39456 7098
rect 39508 7046 39520 7098
rect 39572 7046 44896 7098
rect 1104 7024 44896 7046
rect 9122 6944 9128 6996
rect 9180 6984 9186 6996
rect 23658 6984 23664 6996
rect 9180 6956 23664 6984
rect 9180 6944 9186 6956
rect 23658 6944 23664 6956
rect 23716 6944 23722 6996
rect 25590 6944 25596 6996
rect 25648 6984 25654 6996
rect 33781 6987 33839 6993
rect 25648 6956 31754 6984
rect 25648 6944 25654 6956
rect 22554 6876 22560 6928
rect 22612 6916 22618 6928
rect 27154 6916 27160 6928
rect 22612 6888 27160 6916
rect 22612 6876 22618 6888
rect 27154 6876 27160 6888
rect 27212 6876 27218 6928
rect 31726 6916 31754 6956
rect 33781 6953 33793 6987
rect 33827 6984 33839 6987
rect 34146 6984 34152 6996
rect 33827 6956 34152 6984
rect 33827 6953 33839 6956
rect 33781 6947 33839 6953
rect 34146 6944 34152 6956
rect 34204 6944 34210 6996
rect 34422 6944 34428 6996
rect 34480 6944 34486 6996
rect 34701 6987 34759 6993
rect 34701 6953 34713 6987
rect 34747 6984 34759 6987
rect 34882 6984 34888 6996
rect 34747 6956 34888 6984
rect 34747 6953 34759 6956
rect 34701 6947 34759 6953
rect 34882 6944 34888 6956
rect 34940 6944 34946 6996
rect 35253 6987 35311 6993
rect 35253 6953 35265 6987
rect 35299 6984 35311 6987
rect 35618 6984 35624 6996
rect 35299 6956 35624 6984
rect 35299 6953 35311 6956
rect 35253 6947 35311 6953
rect 35618 6944 35624 6956
rect 35676 6944 35682 6996
rect 37093 6987 37151 6993
rect 37093 6953 37105 6987
rect 37139 6984 37151 6987
rect 37458 6984 37464 6996
rect 37139 6956 37464 6984
rect 37139 6953 37151 6956
rect 37093 6947 37151 6953
rect 37458 6944 37464 6956
rect 37516 6944 37522 6996
rect 37829 6987 37887 6993
rect 37829 6953 37841 6987
rect 37875 6984 37887 6987
rect 38194 6984 38200 6996
rect 37875 6956 38200 6984
rect 37875 6953 37887 6956
rect 37829 6947 37887 6953
rect 38194 6944 38200 6956
rect 38252 6944 38258 6996
rect 38565 6987 38623 6993
rect 38565 6953 38577 6987
rect 38611 6984 38623 6987
rect 38930 6984 38936 6996
rect 38611 6956 38936 6984
rect 38611 6953 38623 6956
rect 38565 6947 38623 6953
rect 38930 6944 38936 6956
rect 38988 6944 38994 6996
rect 44266 6944 44272 6996
rect 44324 6944 44330 6996
rect 34440 6916 34468 6944
rect 31726 6888 34468 6916
rect 35268 6888 36952 6916
rect 842 6808 848 6860
rect 900 6848 906 6860
rect 1765 6851 1823 6857
rect 1765 6848 1777 6851
rect 900 6820 1777 6848
rect 900 6808 906 6820
rect 1765 6817 1777 6820
rect 1811 6817 1823 6851
rect 1765 6811 1823 6817
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 15988 6820 35020 6848
rect 15988 6808 15994 6820
rect 17034 6740 17040 6792
rect 17092 6780 17098 6792
rect 33965 6783 34023 6789
rect 33965 6780 33977 6783
rect 17092 6752 17356 6780
rect 17092 6740 17098 6752
rect 1489 6715 1547 6721
rect 1489 6681 1501 6715
rect 1535 6712 1547 6715
rect 17218 6712 17224 6724
rect 1535 6684 17224 6712
rect 1535 6681 1547 6684
rect 1489 6675 1547 6681
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 17328 6712 17356 6752
rect 33152 6752 33977 6780
rect 33152 6724 33180 6752
rect 33965 6749 33977 6752
rect 34011 6749 34023 6783
rect 33965 6743 34023 6749
rect 17328 6684 31754 6712
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 26602 6644 26608 6656
rect 8352 6616 26608 6644
rect 8352 6604 8358 6616
rect 26602 6604 26608 6616
rect 26660 6604 26666 6656
rect 31726 6644 31754 6684
rect 33134 6672 33140 6724
rect 33192 6672 33198 6724
rect 33980 6712 34008 6743
rect 34606 6740 34612 6792
rect 34664 6780 34670 6792
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 34664 6752 34897 6780
rect 34664 6740 34670 6752
rect 34885 6749 34897 6752
rect 34931 6749 34943 6783
rect 34992 6780 35020 6820
rect 35268 6780 35296 6888
rect 35342 6808 35348 6860
rect 35400 6848 35406 6860
rect 36924 6848 36952 6888
rect 36998 6876 37004 6928
rect 37056 6916 37062 6928
rect 37056 6888 38148 6916
rect 37056 6876 37062 6888
rect 35400 6820 36584 6848
rect 36924 6820 38056 6848
rect 35400 6808 35406 6820
rect 36556 6789 36584 6820
rect 36541 6783 36599 6789
rect 34992 6756 35388 6780
rect 35437 6759 35495 6765
rect 35437 6756 35449 6759
rect 34992 6752 35449 6756
rect 34885 6743 34943 6749
rect 35360 6728 35449 6752
rect 35437 6725 35449 6728
rect 35483 6725 35495 6759
rect 36541 6749 36553 6783
rect 36587 6749 36599 6783
rect 37277 6783 37335 6789
rect 37277 6780 37289 6783
rect 36541 6743 36599 6749
rect 36740 6752 37289 6780
rect 35250 6712 35256 6724
rect 33980 6684 35256 6712
rect 35250 6672 35256 6684
rect 35308 6672 35314 6724
rect 35437 6719 35495 6725
rect 36740 6724 36768 6752
rect 37277 6749 37289 6752
rect 37323 6749 37335 6783
rect 37277 6743 37335 6749
rect 37366 6740 37372 6792
rect 37424 6740 37430 6792
rect 38028 6789 38056 6820
rect 38013 6783 38071 6789
rect 38013 6749 38025 6783
rect 38059 6749 38071 6783
rect 38120 6780 38148 6888
rect 43901 6851 43959 6857
rect 43901 6817 43913 6851
rect 43947 6848 43959 6851
rect 45094 6848 45100 6860
rect 43947 6820 45100 6848
rect 43947 6817 43959 6820
rect 43901 6811 43959 6817
rect 45094 6808 45100 6820
rect 45152 6808 45158 6860
rect 38749 6783 38807 6789
rect 38749 6780 38761 6783
rect 38120 6752 38761 6780
rect 38013 6743 38071 6749
rect 38749 6749 38761 6752
rect 38795 6749 38807 6783
rect 38749 6743 38807 6749
rect 38838 6740 38844 6792
rect 38896 6780 38902 6792
rect 44177 6783 44235 6789
rect 44177 6780 44189 6783
rect 38896 6752 44189 6780
rect 38896 6740 38902 6752
rect 44177 6749 44189 6752
rect 44223 6749 44235 6783
rect 44177 6743 44235 6749
rect 36722 6672 36728 6724
rect 36780 6672 36786 6724
rect 36262 6644 36268 6656
rect 31726 6616 36268 6644
rect 36262 6604 36268 6616
rect 36320 6604 36326 6656
rect 36357 6647 36415 6653
rect 36357 6613 36369 6647
rect 36403 6644 36415 6647
rect 37384 6644 37412 6740
rect 43622 6672 43628 6724
rect 43680 6672 43686 6724
rect 36403 6616 37412 6644
rect 36403 6613 36415 6616
rect 36357 6607 36415 6613
rect 1104 6554 45051 6576
rect 1104 6502 11896 6554
rect 11948 6502 11960 6554
rect 12012 6502 12024 6554
rect 12076 6502 12088 6554
rect 12140 6502 12152 6554
rect 12204 6502 22843 6554
rect 22895 6502 22907 6554
rect 22959 6502 22971 6554
rect 23023 6502 23035 6554
rect 23087 6502 23099 6554
rect 23151 6502 33790 6554
rect 33842 6502 33854 6554
rect 33906 6502 33918 6554
rect 33970 6502 33982 6554
rect 34034 6502 34046 6554
rect 34098 6502 44737 6554
rect 44789 6502 44801 6554
rect 44853 6502 44865 6554
rect 44917 6502 44929 6554
rect 44981 6502 44993 6554
rect 45045 6502 45051 6554
rect 1104 6480 45051 6502
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 34606 6440 34612 6452
rect 16724 6412 34612 6440
rect 16724 6400 16730 6412
rect 34606 6400 34612 6412
rect 34664 6400 34670 6452
rect 36262 6400 36268 6452
rect 36320 6440 36326 6452
rect 38838 6440 38844 6452
rect 36320 6412 38844 6440
rect 36320 6400 36326 6412
rect 38838 6400 38844 6412
rect 38896 6400 38902 6452
rect 18874 6332 18880 6384
rect 18932 6372 18938 6384
rect 33134 6372 33140 6384
rect 18932 6344 33140 6372
rect 18932 6332 18938 6344
rect 33134 6332 33140 6344
rect 33192 6332 33198 6384
rect 34624 6372 34652 6400
rect 36722 6372 36728 6384
rect 34624 6344 36728 6372
rect 36722 6332 36728 6344
rect 36780 6332 36786 6384
rect 6822 6264 6828 6316
rect 6880 6304 6886 6316
rect 25866 6304 25872 6316
rect 6880 6276 25872 6304
rect 6880 6264 6886 6276
rect 25866 6264 25872 6276
rect 25924 6264 25930 6316
rect 16850 6196 16856 6248
rect 16908 6236 16914 6248
rect 35894 6236 35900 6248
rect 16908 6208 35900 6236
rect 16908 6196 16914 6208
rect 35894 6196 35900 6208
rect 35952 6196 35958 6248
rect 3142 6128 3148 6180
rect 3200 6168 3206 6180
rect 27982 6168 27988 6180
rect 3200 6140 27988 6168
rect 3200 6128 3206 6140
rect 27982 6128 27988 6140
rect 28040 6128 28046 6180
rect 19702 6060 19708 6112
rect 19760 6100 19766 6112
rect 33042 6100 33048 6112
rect 19760 6072 33048 6100
rect 19760 6060 19766 6072
rect 33042 6060 33048 6072
rect 33100 6060 33106 6112
rect 1104 6010 44896 6032
rect 1104 5958 6423 6010
rect 6475 5958 6487 6010
rect 6539 5958 6551 6010
rect 6603 5958 6615 6010
rect 6667 5958 6679 6010
rect 6731 5958 17370 6010
rect 17422 5958 17434 6010
rect 17486 5958 17498 6010
rect 17550 5958 17562 6010
rect 17614 5958 17626 6010
rect 17678 5958 28317 6010
rect 28369 5958 28381 6010
rect 28433 5958 28445 6010
rect 28497 5958 28509 6010
rect 28561 5958 28573 6010
rect 28625 5958 39264 6010
rect 39316 5958 39328 6010
rect 39380 5958 39392 6010
rect 39444 5958 39456 6010
rect 39508 5958 39520 6010
rect 39572 5958 44896 6010
rect 1104 5936 44896 5958
rect 19334 5856 19340 5908
rect 19392 5896 19398 5908
rect 30374 5896 30380 5908
rect 19392 5868 30380 5896
rect 19392 5856 19398 5868
rect 30374 5856 30380 5868
rect 30432 5856 30438 5908
rect 43622 5896 43628 5908
rect 41386 5868 43628 5896
rect 25038 5788 25044 5840
rect 25096 5828 25102 5840
rect 37458 5828 37464 5840
rect 25096 5800 37464 5828
rect 25096 5788 25102 5800
rect 37458 5788 37464 5800
rect 37516 5788 37522 5840
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 41386 5760 41414 5868
rect 43622 5856 43628 5868
rect 43680 5856 43686 5908
rect 18104 5732 41414 5760
rect 18104 5720 18110 5732
rect 14458 5652 14464 5704
rect 14516 5692 14522 5704
rect 19242 5692 19248 5704
rect 14516 5664 19248 5692
rect 14516 5652 14522 5664
rect 19242 5652 19248 5664
rect 19300 5652 19306 5704
rect 1104 5466 45051 5488
rect 1104 5414 11896 5466
rect 11948 5414 11960 5466
rect 12012 5414 12024 5466
rect 12076 5414 12088 5466
rect 12140 5414 12152 5466
rect 12204 5414 22843 5466
rect 22895 5414 22907 5466
rect 22959 5414 22971 5466
rect 23023 5414 23035 5466
rect 23087 5414 23099 5466
rect 23151 5414 33790 5466
rect 33842 5414 33854 5466
rect 33906 5414 33918 5466
rect 33970 5414 33982 5466
rect 34034 5414 34046 5466
rect 34098 5414 44737 5466
rect 44789 5414 44801 5466
rect 44853 5414 44865 5466
rect 44917 5414 44929 5466
rect 44981 5414 44993 5466
rect 45045 5414 45051 5466
rect 1104 5392 45051 5414
rect 23290 5176 23296 5228
rect 23348 5216 23354 5228
rect 39022 5216 39028 5228
rect 23348 5188 39028 5216
rect 23348 5176 23354 5188
rect 39022 5176 39028 5188
rect 39080 5176 39086 5228
rect 17862 5108 17868 5160
rect 17920 5148 17926 5160
rect 33410 5148 33416 5160
rect 17920 5120 33416 5148
rect 17920 5108 17926 5120
rect 33410 5108 33416 5120
rect 33468 5108 33474 5160
rect 10870 5040 10876 5092
rect 10928 5080 10934 5092
rect 26970 5080 26976 5092
rect 10928 5052 26976 5080
rect 10928 5040 10934 5052
rect 26970 5040 26976 5052
rect 27028 5040 27034 5092
rect 8386 4972 8392 5024
rect 8444 5012 8450 5024
rect 27062 5012 27068 5024
rect 8444 4984 27068 5012
rect 8444 4972 8450 4984
rect 27062 4972 27068 4984
rect 27120 4972 27126 5024
rect 1104 4922 44896 4944
rect 1104 4870 6423 4922
rect 6475 4870 6487 4922
rect 6539 4870 6551 4922
rect 6603 4870 6615 4922
rect 6667 4870 6679 4922
rect 6731 4870 17370 4922
rect 17422 4870 17434 4922
rect 17486 4870 17498 4922
rect 17550 4870 17562 4922
rect 17614 4870 17626 4922
rect 17678 4870 28317 4922
rect 28369 4870 28381 4922
rect 28433 4870 28445 4922
rect 28497 4870 28509 4922
rect 28561 4870 28573 4922
rect 28625 4870 39264 4922
rect 39316 4870 39328 4922
rect 39380 4870 39392 4922
rect 39444 4870 39456 4922
rect 39508 4870 39520 4922
rect 39572 4870 44896 4922
rect 1104 4848 44896 4870
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 26510 4808 26516 4820
rect 7340 4780 26516 4808
rect 7340 4768 7346 4780
rect 26510 4768 26516 4780
rect 26568 4768 26574 4820
rect 27154 4768 27160 4820
rect 27212 4808 27218 4820
rect 39114 4808 39120 4820
rect 27212 4780 39120 4808
rect 27212 4768 27218 4780
rect 39114 4768 39120 4780
rect 39172 4768 39178 4820
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 21818 4604 21824 4616
rect 13780 4576 21824 4604
rect 13780 4564 13786 4576
rect 21818 4564 21824 4576
rect 21876 4564 21882 4616
rect 10318 4496 10324 4548
rect 10376 4536 10382 4548
rect 23290 4536 23296 4548
rect 10376 4508 23296 4536
rect 10376 4496 10382 4508
rect 23290 4496 23296 4508
rect 23348 4496 23354 4548
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 22646 4468 22652 4480
rect 10928 4440 22652 4468
rect 10928 4428 10934 4440
rect 22646 4428 22652 4440
rect 22704 4428 22710 4480
rect 1104 4378 45051 4400
rect 1104 4326 11896 4378
rect 11948 4326 11960 4378
rect 12012 4326 12024 4378
rect 12076 4326 12088 4378
rect 12140 4326 12152 4378
rect 12204 4326 22843 4378
rect 22895 4326 22907 4378
rect 22959 4326 22971 4378
rect 23023 4326 23035 4378
rect 23087 4326 23099 4378
rect 23151 4326 33790 4378
rect 33842 4326 33854 4378
rect 33906 4326 33918 4378
rect 33970 4326 33982 4378
rect 34034 4326 34046 4378
rect 34098 4326 44737 4378
rect 44789 4326 44801 4378
rect 44853 4326 44865 4378
rect 44917 4326 44929 4378
rect 44981 4326 44993 4378
rect 45045 4326 45051 4378
rect 1104 4304 45051 4326
rect 17218 4224 17224 4276
rect 17276 4264 17282 4276
rect 30742 4264 30748 4276
rect 17276 4236 30748 4264
rect 17276 4224 17282 4236
rect 30742 4224 30748 4236
rect 30800 4224 30806 4276
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 18782 4196 18788 4208
rect 11112 4168 18788 4196
rect 11112 4156 11118 4168
rect 18782 4156 18788 4168
rect 18840 4156 18846 4208
rect 18892 4168 19380 4196
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 18892 4128 18920 4168
rect 9732 4100 18920 4128
rect 9732 4088 9738 4100
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 19352 4128 19380 4168
rect 21284 4168 21772 4196
rect 21284 4128 21312 4168
rect 19352 4100 21312 4128
rect 21361 4131 21419 4137
rect 21361 4097 21373 4131
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 10686 4020 10692 4072
rect 10744 4060 10750 4072
rect 21376 4060 21404 4091
rect 21634 4088 21640 4140
rect 21692 4088 21698 4140
rect 21744 4128 21772 4168
rect 21818 4156 21824 4208
rect 21876 4196 21882 4208
rect 32030 4196 32036 4208
rect 21876 4168 32036 4196
rect 21876 4156 21882 4168
rect 32030 4156 32036 4168
rect 32088 4156 32094 4208
rect 22005 4131 22063 4137
rect 22005 4128 22017 4131
rect 21744 4100 22017 4128
rect 22005 4097 22017 4100
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 26329 4131 26387 4137
rect 26329 4097 26341 4131
rect 26375 4128 26387 4131
rect 26694 4128 26700 4140
rect 26375 4100 26700 4128
rect 26375 4097 26387 4100
rect 26329 4091 26387 4097
rect 26694 4088 26700 4100
rect 26752 4088 26758 4140
rect 26786 4088 26792 4140
rect 26844 4088 26850 4140
rect 32674 4088 32680 4140
rect 32732 4088 32738 4140
rect 31018 4060 31024 4072
rect 10744 4032 21404 4060
rect 23124 4032 31024 4060
rect 10744 4020 10750 4032
rect 23124 4004 23152 4032
rect 31018 4020 31024 4032
rect 31076 4020 31082 4072
rect 16758 3952 16764 4004
rect 16816 3992 16822 4004
rect 18874 3992 18880 4004
rect 16816 3964 18880 3992
rect 16816 3952 16822 3964
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 19058 3952 19064 4004
rect 19116 3952 19122 4004
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 21542 3992 21548 4004
rect 19484 3964 21548 3992
rect 19484 3952 19490 3964
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 23106 3952 23112 4004
rect 23164 3952 23170 4004
rect 23290 3952 23296 4004
rect 23348 3992 23354 4004
rect 24394 3992 24400 4004
rect 23348 3964 24400 3992
rect 23348 3952 23354 3964
rect 24394 3952 24400 3964
rect 24452 3952 24458 4004
rect 26510 3952 26516 4004
rect 26568 3952 26574 4004
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 18785 3927 18843 3933
rect 18785 3924 18797 3927
rect 18564 3896 18797 3924
rect 18564 3884 18570 3896
rect 18785 3893 18797 3896
rect 18831 3893 18843 3927
rect 18785 3887 18843 3893
rect 21174 3884 21180 3936
rect 21232 3884 21238 3936
rect 21450 3884 21456 3936
rect 21508 3884 21514 3936
rect 21821 3927 21879 3933
rect 21821 3893 21833 3927
rect 21867 3924 21879 3927
rect 22094 3924 22100 3936
rect 21867 3896 22100 3924
rect 21867 3893 21879 3896
rect 21821 3887 21879 3893
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 22370 3884 22376 3936
rect 22428 3924 22434 3936
rect 25406 3924 25412 3936
rect 22428 3896 25412 3924
rect 22428 3884 22434 3896
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 26605 3927 26663 3933
rect 26605 3893 26617 3927
rect 26651 3924 26663 3927
rect 27154 3924 27160 3936
rect 26651 3896 27160 3924
rect 26651 3893 26663 3896
rect 26605 3887 26663 3893
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 32493 3927 32551 3933
rect 32493 3893 32505 3927
rect 32539 3924 32551 3927
rect 33410 3924 33416 3936
rect 32539 3896 33416 3924
rect 32539 3893 32551 3896
rect 32493 3887 32551 3893
rect 33410 3884 33416 3896
rect 33468 3884 33474 3936
rect 1104 3834 44896 3856
rect 1104 3782 6423 3834
rect 6475 3782 6487 3834
rect 6539 3782 6551 3834
rect 6603 3782 6615 3834
rect 6667 3782 6679 3834
rect 6731 3782 17370 3834
rect 17422 3782 17434 3834
rect 17486 3782 17498 3834
rect 17550 3782 17562 3834
rect 17614 3782 17626 3834
rect 17678 3782 28317 3834
rect 28369 3782 28381 3834
rect 28433 3782 28445 3834
rect 28497 3782 28509 3834
rect 28561 3782 28573 3834
rect 28625 3782 39264 3834
rect 39316 3782 39328 3834
rect 39380 3782 39392 3834
rect 39444 3782 39456 3834
rect 39508 3782 39520 3834
rect 39572 3782 44896 3834
rect 1104 3760 44896 3782
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 18693 3723 18751 3729
rect 18693 3720 18705 3723
rect 11020 3692 18705 3720
rect 11020 3680 11026 3692
rect 18693 3689 18705 3692
rect 18739 3689 18751 3723
rect 18693 3683 18751 3689
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 19245 3723 19303 3729
rect 18840 3692 19196 3720
rect 18840 3680 18846 3692
rect 16574 3612 16580 3664
rect 16632 3652 16638 3664
rect 16632 3624 16712 3652
rect 16632 3612 16638 3624
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 16540 3488 16589 3516
rect 16540 3476 16546 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16684 3516 16712 3624
rect 16758 3612 16764 3664
rect 16816 3612 16822 3664
rect 16853 3655 16911 3661
rect 16853 3621 16865 3655
rect 16899 3621 16911 3655
rect 16853 3615 16911 3621
rect 17313 3655 17371 3661
rect 17313 3621 17325 3655
rect 17359 3652 17371 3655
rect 17862 3652 17868 3664
rect 17359 3624 17868 3652
rect 17359 3621 17371 3624
rect 17313 3615 17371 3621
rect 16868 3584 16896 3615
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 19168 3652 19196 3692
rect 19245 3689 19257 3723
rect 19291 3720 19303 3723
rect 19794 3720 19800 3732
rect 19291 3692 19800 3720
rect 19291 3689 19303 3692
rect 19245 3683 19303 3689
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 20254 3680 20260 3732
rect 20312 3680 20318 3732
rect 20990 3680 20996 3732
rect 21048 3680 21054 3732
rect 21542 3680 21548 3732
rect 21600 3680 21606 3732
rect 21637 3723 21695 3729
rect 21637 3689 21649 3723
rect 21683 3720 21695 3723
rect 28718 3720 28724 3732
rect 21683 3692 28724 3720
rect 21683 3689 21695 3692
rect 21637 3683 21695 3689
rect 28718 3680 28724 3692
rect 28776 3680 28782 3732
rect 29822 3680 29828 3732
rect 29880 3680 29886 3732
rect 30834 3680 30840 3732
rect 30892 3680 30898 3732
rect 32766 3680 32772 3732
rect 32824 3720 32830 3732
rect 33045 3723 33103 3729
rect 33045 3720 33057 3723
rect 32824 3692 33057 3720
rect 32824 3680 32830 3692
rect 33045 3689 33057 3692
rect 33091 3689 33103 3723
rect 33045 3683 33103 3689
rect 33134 3680 33140 3732
rect 33192 3680 33198 3732
rect 17972 3624 19104 3652
rect 19168 3624 21404 3652
rect 17972 3584 18000 3624
rect 16868 3556 17172 3584
rect 17144 3525 17172 3556
rect 17512 3556 18000 3584
rect 19076 3584 19104 3624
rect 19076 3556 20024 3584
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16684 3488 17049 3516
rect 16577 3479 16635 3485
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 16942 3408 16948 3460
rect 17000 3448 17006 3460
rect 17420 3448 17448 3479
rect 17000 3420 17448 3448
rect 17000 3408 17006 3420
rect 11238 3340 11244 3392
rect 11296 3380 11302 3392
rect 17512 3380 17540 3556
rect 17678 3516 17684 3528
rect 17604 3488 17684 3516
rect 17604 3389 17632 3488
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 17862 3476 17868 3528
rect 17920 3476 17926 3528
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 18156 3448 18184 3479
rect 18414 3476 18420 3528
rect 18472 3476 18478 3528
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 19061 3519 19119 3525
rect 19061 3485 19073 3519
rect 19107 3485 19119 3519
rect 19061 3479 19119 3485
rect 17880 3420 18184 3448
rect 18524 3448 18552 3479
rect 18782 3448 18788 3460
rect 18524 3420 18788 3448
rect 17880 3392 17908 3420
rect 18782 3408 18788 3420
rect 18840 3408 18846 3460
rect 19076 3392 19104 3479
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 19996 3525 20024 3556
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 19981 3519 20039 3525
rect 19981 3485 19993 3519
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 19720 3448 19748 3479
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20404 3488 20545 3516
rect 20404 3476 20410 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21140 3488 21281 3516
rect 21140 3476 21146 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21376 3516 21404 3624
rect 21560 3584 21588 3680
rect 22278 3612 22284 3664
rect 22336 3652 22342 3664
rect 23017 3655 23075 3661
rect 22336 3624 22600 3652
rect 22336 3612 22342 3624
rect 21560 3556 22416 3584
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 21376 3488 21465 3516
rect 21269 3479 21327 3485
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 21542 3476 21548 3528
rect 21600 3516 21606 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21600 3488 21925 3516
rect 21600 3476 21606 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22186 3476 22192 3528
rect 22244 3476 22250 3528
rect 22278 3476 22284 3528
rect 22336 3476 22342 3528
rect 22296 3448 22324 3476
rect 19720 3420 20024 3448
rect 19996 3392 20024 3420
rect 21100 3420 22324 3448
rect 22388 3448 22416 3556
rect 22462 3476 22468 3528
rect 22520 3476 22526 3528
rect 22572 3525 22600 3624
rect 23017 3621 23029 3655
rect 23063 3652 23075 3655
rect 23474 3652 23480 3664
rect 23063 3624 23480 3652
rect 23063 3621 23075 3624
rect 23017 3615 23075 3621
rect 23474 3612 23480 3624
rect 23532 3612 23538 3664
rect 23566 3612 23572 3664
rect 23624 3612 23630 3664
rect 23658 3612 23664 3664
rect 23716 3652 23722 3664
rect 23753 3655 23811 3661
rect 23753 3652 23765 3655
rect 23716 3624 23765 3652
rect 23716 3612 23722 3624
rect 23753 3621 23765 3624
rect 23799 3621 23811 3655
rect 23753 3615 23811 3621
rect 23845 3655 23903 3661
rect 23845 3621 23857 3655
rect 23891 3652 23903 3655
rect 24762 3652 24768 3664
rect 23891 3624 24768 3652
rect 23891 3621 23903 3624
rect 23845 3615 23903 3621
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 24854 3612 24860 3664
rect 24912 3612 24918 3664
rect 25866 3612 25872 3664
rect 25924 3612 25930 3664
rect 26602 3612 26608 3664
rect 26660 3612 26666 3664
rect 26970 3612 26976 3664
rect 27028 3612 27034 3664
rect 27062 3612 27068 3664
rect 27120 3652 27126 3664
rect 27341 3655 27399 3661
rect 27341 3652 27353 3655
rect 27120 3624 27353 3652
rect 27120 3612 27126 3624
rect 27341 3621 27353 3624
rect 27387 3621 27399 3655
rect 27341 3615 27399 3621
rect 27433 3655 27491 3661
rect 27433 3621 27445 3655
rect 27479 3652 27491 3655
rect 28353 3655 28411 3661
rect 27479 3624 28304 3652
rect 27479 3621 27491 3624
rect 27433 3615 27491 3621
rect 23584 3584 23612 3612
rect 23492 3556 23612 3584
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3485 22615 3519
rect 22557 3479 22615 3485
rect 23198 3476 23204 3528
rect 23256 3476 23262 3528
rect 23492 3525 23520 3556
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3516 23627 3519
rect 23615 3488 23980 3516
rect 23615 3485 23627 3488
rect 23569 3479 23627 3485
rect 23952 3448 23980 3488
rect 24026 3476 24032 3528
rect 24084 3476 24090 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 24360 3488 24685 3516
rect 24360 3476 24366 3488
rect 24673 3485 24685 3488
rect 24719 3485 24731 3519
rect 24872 3516 24900 3612
rect 25130 3544 25136 3596
rect 25188 3584 25194 3596
rect 27706 3584 27712 3596
rect 25188 3556 25544 3584
rect 25188 3544 25194 3556
rect 24949 3519 25007 3525
rect 24949 3516 24961 3519
rect 24872 3488 24961 3516
rect 24673 3479 24731 3485
rect 24949 3485 24961 3488
rect 24995 3485 25007 3519
rect 24949 3479 25007 3485
rect 25222 3476 25228 3528
rect 25280 3476 25286 3528
rect 25516 3525 25544 3556
rect 26436 3556 27712 3584
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3485 25559 3519
rect 25501 3479 25559 3485
rect 25682 3476 25688 3528
rect 25740 3476 25746 3528
rect 26145 3519 26203 3525
rect 26145 3485 26157 3519
rect 26191 3485 26203 3519
rect 26145 3479 26203 3485
rect 24118 3448 24124 3460
rect 22388 3420 23428 3448
rect 23952 3420 24124 3448
rect 11296 3352 17540 3380
rect 17589 3383 17647 3389
rect 11296 3340 11302 3352
rect 17589 3349 17601 3383
rect 17635 3349 17647 3383
rect 17589 3343 17647 3349
rect 17678 3340 17684 3392
rect 17736 3340 17742 3392
rect 17862 3340 17868 3392
rect 17920 3340 17926 3392
rect 17954 3340 17960 3392
rect 18012 3340 18018 3392
rect 18230 3340 18236 3392
rect 18288 3340 18294 3392
rect 18874 3340 18880 3392
rect 18932 3340 18938 3392
rect 19058 3340 19064 3392
rect 19116 3340 19122 3392
rect 19518 3340 19524 3392
rect 19576 3340 19582 3392
rect 19794 3340 19800 3392
rect 19852 3340 19858 3392
rect 19978 3340 19984 3392
rect 20036 3340 20042 3392
rect 20349 3383 20407 3389
rect 20349 3349 20361 3383
rect 20395 3380 20407 3383
rect 20898 3380 20904 3392
rect 20395 3352 20904 3380
rect 20395 3349 20407 3352
rect 20349 3343 20407 3349
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 21100 3389 21128 3420
rect 21085 3383 21143 3389
rect 21085 3349 21097 3383
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 21726 3340 21732 3392
rect 21784 3340 21790 3392
rect 22002 3340 22008 3392
rect 22060 3340 22066 3392
rect 22278 3340 22284 3392
rect 22336 3340 22342 3392
rect 22738 3340 22744 3392
rect 22796 3340 22802 3392
rect 23106 3340 23112 3392
rect 23164 3380 23170 3392
rect 23293 3383 23351 3389
rect 23293 3380 23305 3383
rect 23164 3352 23305 3380
rect 23164 3340 23170 3352
rect 23293 3349 23305 3352
rect 23339 3349 23351 3383
rect 23400 3380 23428 3420
rect 24118 3408 24124 3420
rect 24176 3408 24182 3460
rect 26160 3448 26188 3479
rect 26436 3457 26464 3556
rect 27706 3544 27712 3556
rect 27764 3544 27770 3596
rect 27798 3544 27804 3596
rect 27856 3544 27862 3596
rect 28276 3584 28304 3624
rect 28353 3621 28365 3655
rect 28399 3652 28411 3655
rect 29454 3652 29460 3664
rect 28399 3624 29460 3652
rect 28399 3621 28411 3624
rect 28353 3615 28411 3621
rect 29454 3612 29460 3624
rect 29512 3612 29518 3664
rect 31573 3655 31631 3661
rect 31573 3621 31585 3655
rect 31619 3652 31631 3655
rect 33152 3652 33180 3680
rect 31619 3624 33180 3652
rect 31619 3621 31631 3624
rect 31573 3615 31631 3621
rect 28276 3556 28948 3584
rect 27157 3519 27215 3525
rect 27157 3485 27169 3519
rect 27203 3516 27215 3519
rect 27522 3516 27528 3528
rect 27203 3488 27528 3516
rect 27203 3485 27215 3488
rect 27157 3479 27215 3485
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 27614 3476 27620 3528
rect 27672 3476 27678 3528
rect 27816 3516 27844 3544
rect 27893 3519 27951 3525
rect 27893 3516 27905 3519
rect 27816 3488 27905 3516
rect 27893 3485 27905 3488
rect 27939 3485 27951 3519
rect 27893 3479 27951 3485
rect 28000 3488 28212 3516
rect 24228 3420 26188 3448
rect 26421 3451 26479 3457
rect 24228 3380 24256 3420
rect 26421 3417 26433 3451
rect 26467 3417 26479 3451
rect 26421 3411 26479 3417
rect 26786 3408 26792 3460
rect 26844 3408 26850 3460
rect 27338 3408 27344 3460
rect 27396 3448 27402 3460
rect 28000 3448 28028 3488
rect 27396 3420 28028 3448
rect 28077 3451 28135 3457
rect 27396 3408 27402 3420
rect 28077 3417 28089 3451
rect 28123 3417 28135 3451
rect 28184 3448 28212 3488
rect 28258 3476 28264 3528
rect 28316 3516 28322 3528
rect 28537 3519 28595 3525
rect 28537 3516 28549 3519
rect 28316 3488 28549 3516
rect 28316 3476 28322 3488
rect 28537 3485 28549 3488
rect 28583 3485 28595 3519
rect 28537 3479 28595 3485
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3485 28871 3519
rect 28813 3479 28871 3485
rect 28828 3448 28856 3479
rect 28184 3420 28856 3448
rect 28920 3448 28948 3556
rect 28994 3544 29000 3596
rect 29052 3544 29058 3596
rect 29178 3544 29184 3596
rect 29236 3544 29242 3596
rect 30558 3584 30564 3596
rect 29564 3556 30564 3584
rect 29012 3516 29040 3544
rect 29089 3519 29147 3525
rect 29089 3516 29101 3519
rect 29012 3488 29101 3516
rect 29089 3485 29101 3488
rect 29135 3485 29147 3519
rect 29196 3516 29224 3544
rect 29365 3519 29423 3525
rect 29365 3516 29377 3519
rect 29196 3488 29377 3516
rect 29089 3479 29147 3485
rect 29365 3485 29377 3488
rect 29411 3485 29423 3519
rect 29365 3479 29423 3485
rect 29564 3448 29592 3556
rect 30558 3544 30564 3556
rect 30616 3544 30622 3596
rect 35434 3584 35440 3596
rect 30760 3556 35440 3584
rect 29638 3476 29644 3528
rect 29696 3516 29702 3528
rect 30193 3519 30251 3525
rect 30193 3516 30205 3519
rect 29696 3488 30205 3516
rect 29696 3476 29702 3488
rect 30193 3485 30205 3488
rect 30239 3485 30251 3519
rect 30193 3479 30251 3485
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 30760 3525 30788 3556
rect 35434 3544 35440 3556
rect 35492 3544 35498 3596
rect 30469 3519 30527 3525
rect 30469 3516 30481 3519
rect 30340 3488 30481 3516
rect 30340 3476 30346 3488
rect 30469 3485 30481 3488
rect 30515 3485 30527 3519
rect 30469 3479 30527 3485
rect 30745 3519 30803 3525
rect 30745 3485 30757 3519
rect 30791 3485 30803 3519
rect 30745 3479 30803 3485
rect 31202 3476 31208 3528
rect 31260 3476 31266 3528
rect 31478 3476 31484 3528
rect 31536 3476 31542 3528
rect 31754 3476 31760 3528
rect 31812 3476 31818 3528
rect 32030 3476 32036 3528
rect 32088 3476 32094 3528
rect 32306 3476 32312 3528
rect 32364 3476 32370 3528
rect 32582 3476 32588 3528
rect 32640 3476 32646 3528
rect 28920 3420 29592 3448
rect 29733 3451 29791 3457
rect 28077 3411 28135 3417
rect 29733 3417 29745 3451
rect 29779 3448 29791 3451
rect 30650 3448 30656 3460
rect 29779 3420 30656 3448
rect 29779 3417 29791 3420
rect 29733 3411 29791 3417
rect 23400 3352 24256 3380
rect 23293 3343 23351 3349
rect 24486 3340 24492 3392
rect 24544 3340 24550 3392
rect 24762 3340 24768 3392
rect 24820 3340 24826 3392
rect 25038 3340 25044 3392
rect 25096 3340 25102 3392
rect 25314 3340 25320 3392
rect 25372 3340 25378 3392
rect 25958 3340 25964 3392
rect 26016 3340 26022 3392
rect 27706 3340 27712 3392
rect 27764 3340 27770 3392
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 28092 3380 28120 3411
rect 30650 3408 30656 3420
rect 30708 3408 30714 3460
rect 32490 3448 32496 3460
rect 31036 3420 32496 3448
rect 28040 3352 28120 3380
rect 28040 3340 28046 3352
rect 28166 3340 28172 3392
rect 28224 3340 28230 3392
rect 28626 3340 28632 3392
rect 28684 3340 28690 3392
rect 28902 3340 28908 3392
rect 28960 3340 28966 3392
rect 29178 3340 29184 3392
rect 29236 3340 29242 3392
rect 30006 3340 30012 3392
rect 30064 3340 30070 3392
rect 30282 3340 30288 3392
rect 30340 3340 30346 3392
rect 31036 3389 31064 3420
rect 32490 3408 32496 3420
rect 32548 3408 32554 3460
rect 32950 3408 32956 3460
rect 33008 3408 33014 3460
rect 31021 3383 31079 3389
rect 31021 3349 31033 3383
rect 31067 3349 31079 3383
rect 31021 3343 31079 3349
rect 31294 3340 31300 3392
rect 31352 3340 31358 3392
rect 31846 3340 31852 3392
rect 31904 3340 31910 3392
rect 32122 3340 32128 3392
rect 32180 3340 32186 3392
rect 32401 3383 32459 3389
rect 32401 3349 32413 3383
rect 32447 3380 32459 3383
rect 32858 3380 32864 3392
rect 32447 3352 32864 3380
rect 32447 3349 32459 3352
rect 32401 3343 32459 3349
rect 32858 3340 32864 3352
rect 32916 3340 32922 3392
rect 1104 3290 45051 3312
rect 1104 3238 11896 3290
rect 11948 3238 11960 3290
rect 12012 3238 12024 3290
rect 12076 3238 12088 3290
rect 12140 3238 12152 3290
rect 12204 3238 22843 3290
rect 22895 3238 22907 3290
rect 22959 3238 22971 3290
rect 23023 3238 23035 3290
rect 23087 3238 23099 3290
rect 23151 3238 33790 3290
rect 33842 3238 33854 3290
rect 33906 3238 33918 3290
rect 33970 3238 33982 3290
rect 34034 3238 34046 3290
rect 34098 3238 44737 3290
rect 44789 3238 44801 3290
rect 44853 3238 44865 3290
rect 44917 3238 44929 3290
rect 44981 3238 44993 3290
rect 45045 3238 45051 3290
rect 1104 3216 45051 3238
rect 13722 3136 13728 3188
rect 13780 3136 13786 3188
rect 14550 3136 14556 3188
rect 14608 3136 14614 3188
rect 17126 3136 17132 3188
rect 17184 3136 17190 3188
rect 17218 3136 17224 3188
rect 17276 3136 17282 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 13538 3000 13544 3052
rect 13596 3000 13602 3052
rect 14366 3000 14372 3052
rect 14424 3000 14430 3052
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16850 3040 16856 3052
rect 15979 3012 16856 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 17144 3040 17172 3136
rect 17083 3012 17172 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 15654 2932 15660 2984
rect 15712 2932 15718 2984
rect 16960 2972 16988 3003
rect 17218 2972 17224 2984
rect 16960 2944 17224 2972
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 17328 2972 17356 3139
rect 17954 3136 17960 3188
rect 18012 3136 18018 3188
rect 18138 3136 18144 3188
rect 18196 3136 18202 3188
rect 18524 3148 18828 3176
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 17972 3108 18000 3136
rect 18049 3111 18107 3117
rect 18049 3108 18061 3111
rect 17736 3080 17781 3108
rect 17972 3080 18061 3108
rect 17736 3068 17742 3080
rect 18049 3077 18061 3080
rect 18095 3077 18107 3111
rect 18049 3071 18107 3077
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 18524 3108 18552 3148
rect 18800 3117 18828 3148
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 19576 3148 20208 3176
rect 19576 3136 19582 3148
rect 18288 3080 18552 3108
rect 18785 3111 18843 3117
rect 18288 3068 18294 3080
rect 18785 3077 18797 3111
rect 18831 3077 18843 3111
rect 18785 3071 18843 3077
rect 18874 3068 18880 3120
rect 18932 3108 18938 3120
rect 20180 3117 20208 3148
rect 21450 3136 21456 3188
rect 21508 3136 21514 3188
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 21784 3148 22094 3176
rect 21784 3136 21790 3148
rect 19705 3111 19763 3117
rect 19705 3108 19717 3111
rect 18932 3080 19717 3108
rect 18932 3068 18938 3080
rect 19705 3077 19717 3080
rect 19751 3077 19763 3111
rect 19705 3071 19763 3077
rect 20165 3111 20223 3117
rect 20165 3077 20177 3111
rect 20211 3077 20223 3111
rect 20165 3071 20223 3077
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 18138 3040 18144 3052
rect 17543 3012 18144 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 18417 3003 18475 3009
rect 18984 3012 19165 3040
rect 18432 2972 18460 3003
rect 17328 2944 18460 2972
rect 18506 2932 18512 2984
rect 18564 2932 18570 2984
rect 9309 2907 9367 2913
rect 9309 2873 9321 2907
rect 9355 2904 9367 2907
rect 17954 2904 17960 2916
rect 9355 2876 17960 2904
rect 9355 2873 9367 2876
rect 9309 2867 9367 2873
rect 17954 2864 17960 2876
rect 18012 2864 18018 2916
rect 18322 2864 18328 2916
rect 18380 2864 18386 2916
rect 18524 2904 18552 2932
rect 18984 2904 19012 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 20717 3043 20775 3049
rect 20717 3040 20729 3043
rect 19153 3003 19211 3009
rect 19260 3012 20729 3040
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19260 2972 19288 3012
rect 20717 3009 20729 3012
rect 20763 3009 20775 3043
rect 20717 3003 20775 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 19116 2944 19288 2972
rect 19337 2975 19395 2981
rect 19116 2932 19122 2944
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19610 2972 19616 2984
rect 19383 2944 19616 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 19702 2932 19708 2984
rect 19760 2972 19766 2984
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 19760 2944 19901 2972
rect 19760 2932 19766 2944
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 19978 2932 19984 2984
rect 20036 2972 20042 2984
rect 21284 2972 21312 3003
rect 20036 2944 21312 2972
rect 21468 2972 21496 3136
rect 22066 3108 22094 3148
rect 22278 3136 22284 3188
rect 22336 3176 22342 3188
rect 22336 3148 23336 3176
rect 22336 3136 22342 3148
rect 23308 3117 23336 3148
rect 23750 3136 23756 3188
rect 23808 3136 23814 3188
rect 24026 3136 24032 3188
rect 24084 3136 24090 3188
rect 24486 3136 24492 3188
rect 24544 3136 24550 3188
rect 25314 3136 25320 3188
rect 25372 3136 25378 3188
rect 25406 3136 25412 3188
rect 25464 3176 25470 3188
rect 25464 3148 25912 3176
rect 25464 3136 25470 3148
rect 22741 3111 22799 3117
rect 22741 3108 22753 3111
rect 22066 3080 22753 3108
rect 22741 3077 22753 3080
rect 22787 3077 22799 3111
rect 22741 3071 22799 3077
rect 23293 3111 23351 3117
rect 23293 3077 23305 3111
rect 23339 3077 23351 3111
rect 23768 3108 23796 3136
rect 24504 3108 24532 3136
rect 25225 3111 25283 3117
rect 25225 3108 25237 3111
rect 23768 3080 24256 3108
rect 24504 3080 25237 3108
rect 23293 3071 23351 3077
rect 22002 3000 22008 3052
rect 22060 3000 22066 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 22204 2972 22232 3003
rect 22462 3000 22468 3052
rect 22520 3000 22526 3052
rect 22646 3000 22652 3052
rect 22704 3040 22710 3052
rect 24228 3049 24256 3080
rect 25225 3077 25237 3080
rect 25271 3077 25283 3111
rect 25332 3108 25360 3136
rect 25777 3111 25835 3117
rect 25777 3108 25789 3111
rect 25332 3080 25789 3108
rect 25225 3071 25283 3077
rect 25777 3077 25789 3080
rect 25823 3077 25835 3111
rect 25884 3108 25912 3148
rect 25958 3136 25964 3188
rect 26016 3176 26022 3188
rect 26016 3148 27108 3176
rect 26016 3136 26022 3148
rect 27080 3117 27108 3148
rect 27154 3136 27160 3188
rect 27212 3136 27218 3188
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 28261 3179 28319 3185
rect 28261 3176 28273 3179
rect 27580 3148 28273 3176
rect 27580 3136 27586 3148
rect 28261 3145 28273 3148
rect 28307 3145 28319 3179
rect 28261 3139 28319 3145
rect 28626 3136 28632 3188
rect 28684 3136 28690 3188
rect 29178 3136 29184 3188
rect 29236 3136 29242 3188
rect 29730 3136 29736 3188
rect 29788 3176 29794 3188
rect 30469 3179 30527 3185
rect 30469 3176 30481 3179
rect 29788 3148 30481 3176
rect 29788 3136 29794 3148
rect 30469 3145 30481 3148
rect 30515 3145 30527 3179
rect 30469 3139 30527 3145
rect 30558 3136 30564 3188
rect 30616 3136 30622 3188
rect 31294 3136 31300 3188
rect 31352 3176 31358 3188
rect 31352 3148 31754 3176
rect 31352 3136 31358 3148
rect 26329 3111 26387 3117
rect 26329 3108 26341 3111
rect 25884 3080 26341 3108
rect 25777 3071 25835 3077
rect 26329 3077 26341 3080
rect 26375 3077 26387 3111
rect 26329 3071 26387 3077
rect 27065 3111 27123 3117
rect 27065 3077 27077 3111
rect 27111 3077 27123 3111
rect 27172 3108 27200 3136
rect 27617 3111 27675 3117
rect 27617 3108 27629 3111
rect 27172 3080 27629 3108
rect 27065 3071 27123 3077
rect 27617 3077 27629 3080
rect 27663 3077 27675 3111
rect 27617 3071 27675 3077
rect 27706 3068 27712 3120
rect 27764 3108 27770 3120
rect 28644 3108 28672 3136
rect 29196 3108 29224 3136
rect 29825 3111 29883 3117
rect 29825 3108 29837 3111
rect 27764 3080 28304 3108
rect 28644 3080 29040 3108
rect 29196 3080 29837 3108
rect 27764 3068 27770 3080
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 22704 3012 23949 3040
rect 22704 3000 22710 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 24394 3000 24400 3052
rect 24452 3040 24458 3052
rect 24489 3043 24547 3049
rect 24489 3040 24501 3043
rect 24452 3012 24501 3040
rect 24452 3000 24458 3012
rect 24489 3009 24501 3012
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 24673 3043 24731 3049
rect 24673 3009 24685 3043
rect 24719 3009 24731 3043
rect 24673 3003 24731 3009
rect 28169 3043 28227 3049
rect 28169 3009 28181 3043
rect 28215 3009 28227 3043
rect 28276 3040 28304 3080
rect 28721 3043 28779 3049
rect 28721 3040 28733 3043
rect 28276 3012 28733 3040
rect 28169 3003 28227 3009
rect 28721 3009 28733 3012
rect 28767 3009 28779 3043
rect 29012 3040 29040 3080
rect 29825 3077 29837 3080
rect 29871 3077 29883 3111
rect 29825 3071 29883 3077
rect 30006 3068 30012 3120
rect 30064 3068 30070 3120
rect 30374 3068 30380 3120
rect 30432 3068 30438 3120
rect 29273 3043 29331 3049
rect 29273 3040 29285 3043
rect 29012 3012 29285 3040
rect 28721 3003 28779 3009
rect 29273 3009 29285 3012
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 21468 2944 22232 2972
rect 20036 2932 20042 2944
rect 18524 2876 19012 2904
rect 19150 2864 19156 2916
rect 19208 2904 19214 2916
rect 22480 2904 22508 3000
rect 24688 2972 24716 3003
rect 23768 2944 24716 2972
rect 28184 2972 28212 3003
rect 30024 2972 30052 3068
rect 28184 2944 30052 2972
rect 30576 2972 30604 3136
rect 30650 3068 30656 3120
rect 30708 3108 30714 3120
rect 31386 3108 31392 3120
rect 30708 3080 31392 3108
rect 30708 3068 30714 3080
rect 31386 3068 31392 3080
rect 31444 3068 31450 3120
rect 31726 3108 31754 3148
rect 31846 3136 31852 3188
rect 31904 3176 31910 3188
rect 31904 3148 32812 3176
rect 31904 3136 31910 3148
rect 32217 3111 32275 3117
rect 32217 3108 32229 3111
rect 31726 3080 32229 3108
rect 32217 3077 32229 3080
rect 32263 3077 32275 3111
rect 32217 3071 32275 3077
rect 32490 3068 32496 3120
rect 32548 3108 32554 3120
rect 32674 3108 32680 3120
rect 32548 3080 32680 3108
rect 32548 3068 32554 3080
rect 32674 3068 32680 3080
rect 32732 3068 32738 3120
rect 32784 3117 32812 3148
rect 32858 3136 32864 3188
rect 32916 3136 32922 3188
rect 33594 3136 33600 3188
rect 33652 3176 33658 3188
rect 34517 3179 34575 3185
rect 34517 3176 34529 3179
rect 33652 3148 34529 3176
rect 33652 3136 33658 3148
rect 34517 3145 34529 3148
rect 34563 3145 34575 3179
rect 34517 3139 34575 3145
rect 35434 3136 35440 3188
rect 35492 3136 35498 3188
rect 39114 3136 39120 3188
rect 39172 3136 39178 3188
rect 32769 3111 32827 3117
rect 32769 3077 32781 3111
rect 32815 3077 32827 3111
rect 32876 3108 32904 3136
rect 34425 3111 34483 3117
rect 34425 3108 34437 3111
rect 32876 3080 34437 3108
rect 32769 3071 32827 3077
rect 34425 3077 34437 3080
rect 34471 3077 34483 3111
rect 34425 3071 34483 3077
rect 30742 3000 30748 3052
rect 30800 3040 30806 3052
rect 30929 3043 30987 3049
rect 30929 3040 30941 3043
rect 30800 3012 30941 3040
rect 30800 3000 30806 3012
rect 30929 3009 30941 3012
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 31018 3000 31024 3052
rect 31076 3040 31082 3052
rect 31481 3043 31539 3049
rect 31481 3040 31493 3043
rect 31076 3012 31493 3040
rect 31076 3000 31082 3012
rect 31481 3009 31493 3012
rect 31527 3009 31539 3043
rect 31481 3003 31539 3009
rect 32122 3000 32128 3052
rect 32180 3040 32186 3052
rect 32858 3040 32864 3052
rect 32180 3012 32864 3040
rect 32180 3000 32186 3012
rect 32858 3000 32864 3012
rect 32916 3000 32922 3052
rect 33321 3043 33379 3049
rect 33321 3009 33333 3043
rect 33367 3009 33379 3043
rect 33321 3003 33379 3009
rect 33336 2972 33364 3003
rect 33410 3000 33416 3052
rect 33468 3040 33474 3052
rect 33873 3043 33931 3049
rect 33873 3040 33885 3043
rect 33468 3012 33885 3040
rect 33468 3000 33474 3012
rect 33873 3009 33885 3012
rect 33919 3009 33931 3043
rect 33873 3003 33931 3009
rect 34330 3000 34336 3052
rect 34388 3040 34394 3052
rect 34977 3043 35035 3049
rect 34977 3040 34989 3043
rect 34388 3012 34989 3040
rect 34388 3000 34394 3012
rect 34977 3009 34989 3012
rect 35023 3009 35035 3043
rect 34977 3003 35035 3009
rect 35066 3000 35072 3052
rect 35124 3040 35130 3052
rect 35621 3043 35679 3049
rect 35621 3040 35633 3043
rect 35124 3012 35633 3040
rect 35124 3000 35130 3012
rect 35621 3009 35633 3012
rect 35667 3009 35679 3043
rect 35621 3003 35679 3009
rect 38930 3000 38936 3052
rect 38988 3000 38994 3052
rect 30576 2944 33364 2972
rect 19208 2876 22508 2904
rect 19208 2864 19214 2876
rect 22646 2864 22652 2916
rect 22704 2904 22710 2916
rect 23768 2913 23796 2944
rect 23753 2907 23811 2913
rect 22704 2876 23520 2904
rect 22704 2864 22710 2876
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 16390 2836 16396 2848
rect 14608 2808 16396 2836
rect 14608 2796 14614 2808
rect 16390 2796 16396 2808
rect 16448 2796 16454 2848
rect 16761 2839 16819 2845
rect 16761 2805 16773 2839
rect 16807 2836 16819 2839
rect 17126 2836 17132 2848
rect 16807 2808 17132 2836
rect 16807 2805 16819 2808
rect 16761 2799 16819 2805
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 17773 2839 17831 2845
rect 17773 2836 17785 2839
rect 17368 2808 17785 2836
rect 17368 2796 17374 2808
rect 17773 2805 17785 2808
rect 17819 2805 17831 2839
rect 18340 2836 18368 2864
rect 18509 2839 18567 2845
rect 18509 2836 18521 2839
rect 18340 2808 18521 2836
rect 17773 2799 17831 2805
rect 18509 2805 18521 2808
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 18877 2839 18935 2845
rect 18877 2836 18889 2839
rect 18748 2808 18889 2836
rect 18748 2796 18754 2808
rect 18877 2805 18889 2808
rect 18923 2805 18935 2839
rect 18877 2799 18935 2805
rect 20254 2796 20260 2848
rect 20312 2796 20318 2848
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 20809 2839 20867 2845
rect 20809 2836 20821 2839
rect 20680 2808 20821 2836
rect 20680 2796 20686 2808
rect 20809 2805 20821 2808
rect 20855 2805 20867 2839
rect 20809 2799 20867 2805
rect 21358 2796 21364 2848
rect 21416 2796 21422 2848
rect 21818 2796 21824 2848
rect 21876 2796 21882 2848
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 22281 2839 22339 2845
rect 22281 2836 22293 2839
rect 22060 2808 22293 2836
rect 22060 2796 22066 2808
rect 22281 2805 22293 2808
rect 22327 2805 22339 2839
rect 22281 2799 22339 2805
rect 22554 2796 22560 2848
rect 22612 2836 22618 2848
rect 22833 2839 22891 2845
rect 22833 2836 22845 2839
rect 22612 2808 22845 2836
rect 22612 2796 22618 2808
rect 22833 2805 22845 2808
rect 22879 2805 22891 2839
rect 22833 2799 22891 2805
rect 23382 2796 23388 2848
rect 23440 2796 23446 2848
rect 23492 2836 23520 2876
rect 23753 2873 23765 2907
rect 23799 2873 23811 2907
rect 25406 2904 25412 2916
rect 23753 2867 23811 2873
rect 24320 2876 25412 2904
rect 24210 2836 24216 2848
rect 23492 2808 24216 2836
rect 24210 2796 24216 2808
rect 24268 2796 24274 2848
rect 24320 2845 24348 2876
rect 25406 2864 25412 2876
rect 25464 2864 25470 2916
rect 26970 2864 26976 2916
rect 27028 2904 27034 2916
rect 27028 2876 27752 2904
rect 27028 2864 27034 2876
rect 24305 2839 24363 2845
rect 24305 2805 24317 2839
rect 24351 2805 24363 2839
rect 24305 2799 24363 2805
rect 24486 2796 24492 2848
rect 24544 2836 24550 2848
rect 24765 2839 24823 2845
rect 24765 2836 24777 2839
rect 24544 2808 24777 2836
rect 24544 2796 24550 2808
rect 24765 2805 24777 2808
rect 24811 2805 24823 2839
rect 24765 2799 24823 2805
rect 25038 2796 25044 2848
rect 25096 2836 25102 2848
rect 25317 2839 25375 2845
rect 25317 2836 25329 2839
rect 25096 2808 25329 2836
rect 25096 2796 25102 2808
rect 25317 2805 25329 2808
rect 25363 2805 25375 2839
rect 25317 2799 25375 2805
rect 25590 2796 25596 2848
rect 25648 2836 25654 2848
rect 25869 2839 25927 2845
rect 25869 2836 25881 2839
rect 25648 2808 25881 2836
rect 25648 2796 25654 2808
rect 25869 2805 25881 2808
rect 25915 2805 25927 2839
rect 25869 2799 25927 2805
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26421 2839 26479 2845
rect 26421 2836 26433 2839
rect 26108 2808 26433 2836
rect 26108 2796 26114 2808
rect 26421 2805 26433 2808
rect 26467 2805 26479 2839
rect 26421 2799 26479 2805
rect 26602 2796 26608 2848
rect 26660 2836 26666 2848
rect 27724 2845 27752 2876
rect 29178 2864 29184 2916
rect 29236 2904 29242 2916
rect 29236 2876 29960 2904
rect 29236 2864 29242 2876
rect 27157 2839 27215 2845
rect 27157 2836 27169 2839
rect 26660 2808 27169 2836
rect 26660 2796 26666 2808
rect 27157 2805 27169 2808
rect 27203 2805 27215 2839
rect 27157 2799 27215 2805
rect 27709 2839 27767 2845
rect 27709 2805 27721 2839
rect 27755 2805 27767 2839
rect 27709 2799 27767 2805
rect 28442 2796 28448 2848
rect 28500 2836 28506 2848
rect 28813 2839 28871 2845
rect 28813 2836 28825 2839
rect 28500 2808 28825 2836
rect 28500 2796 28506 2808
rect 28813 2805 28825 2808
rect 28859 2805 28871 2839
rect 28813 2799 28871 2805
rect 28902 2796 28908 2848
rect 28960 2836 28966 2848
rect 29932 2845 29960 2876
rect 30558 2864 30564 2916
rect 30616 2904 30622 2916
rect 30616 2876 31616 2904
rect 30616 2864 30622 2876
rect 29365 2839 29423 2845
rect 29365 2836 29377 2839
rect 28960 2808 29377 2836
rect 28960 2796 28966 2808
rect 29365 2805 29377 2808
rect 29411 2805 29423 2839
rect 29365 2799 29423 2805
rect 29917 2839 29975 2845
rect 29917 2805 29929 2839
rect 29963 2805 29975 2839
rect 29917 2799 29975 2805
rect 30190 2796 30196 2848
rect 30248 2836 30254 2848
rect 31588 2845 31616 2876
rect 32030 2864 32036 2916
rect 32088 2904 32094 2916
rect 32953 2907 33011 2913
rect 32953 2904 32965 2907
rect 32088 2876 32965 2904
rect 32088 2864 32094 2876
rect 32953 2873 32965 2876
rect 32999 2873 33011 2907
rect 32953 2867 33011 2873
rect 33042 2864 33048 2916
rect 33100 2904 33106 2916
rect 33100 2876 34008 2904
rect 33100 2864 33106 2876
rect 31021 2839 31079 2845
rect 31021 2836 31033 2839
rect 30248 2808 31033 2836
rect 30248 2796 30254 2808
rect 31021 2805 31033 2808
rect 31067 2805 31079 2839
rect 31021 2799 31079 2805
rect 31573 2839 31631 2845
rect 31573 2805 31585 2839
rect 31619 2805 31631 2839
rect 31573 2799 31631 2805
rect 31662 2796 31668 2848
rect 31720 2836 31726 2848
rect 32309 2839 32367 2845
rect 32309 2836 32321 2839
rect 31720 2808 32321 2836
rect 31720 2796 31726 2808
rect 32309 2805 32321 2808
rect 32355 2805 32367 2839
rect 32309 2799 32367 2805
rect 32490 2796 32496 2848
rect 32548 2836 32554 2848
rect 33980 2845 34008 2876
rect 33413 2839 33471 2845
rect 33413 2836 33425 2839
rect 32548 2808 33425 2836
rect 32548 2796 32554 2808
rect 33413 2805 33425 2808
rect 33459 2805 33471 2839
rect 33413 2799 33471 2805
rect 33965 2839 34023 2845
rect 33965 2805 33977 2839
rect 34011 2805 34023 2839
rect 33965 2799 34023 2805
rect 34146 2796 34152 2848
rect 34204 2836 34210 2848
rect 35069 2839 35127 2845
rect 35069 2836 35081 2839
rect 34204 2808 35081 2836
rect 34204 2796 34210 2808
rect 35069 2805 35081 2808
rect 35115 2805 35127 2839
rect 35069 2799 35127 2805
rect 1104 2746 44896 2768
rect 1104 2694 6423 2746
rect 6475 2694 6487 2746
rect 6539 2694 6551 2746
rect 6603 2694 6615 2746
rect 6667 2694 6679 2746
rect 6731 2694 17370 2746
rect 17422 2694 17434 2746
rect 17486 2694 17498 2746
rect 17550 2694 17562 2746
rect 17614 2694 17626 2746
rect 17678 2694 28317 2746
rect 28369 2694 28381 2746
rect 28433 2694 28445 2746
rect 28497 2694 28509 2746
rect 28561 2694 28573 2746
rect 28625 2694 39264 2746
rect 39316 2694 39328 2746
rect 39380 2694 39392 2746
rect 39444 2694 39456 2746
rect 39508 2694 39520 2746
rect 39572 2694 44896 2746
rect 1104 2672 44896 2694
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6730 2632 6736 2644
rect 6595 2604 6736 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 9582 2632 9588 2644
rect 6840 2604 9588 2632
rect 5905 2567 5963 2573
rect 5905 2533 5917 2567
rect 5951 2564 5963 2567
rect 6840 2564 6868 2604
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 9674 2592 9680 2644
rect 9732 2592 9738 2644
rect 9950 2592 9956 2644
rect 10008 2592 10014 2644
rect 12986 2632 12992 2644
rect 10336 2604 12992 2632
rect 5951 2536 6868 2564
rect 7101 2567 7159 2573
rect 5951 2533 5963 2536
rect 5905 2527 5963 2533
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 10226 2564 10232 2576
rect 7147 2536 10232 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10336 2573 10364 2604
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 13170 2592 13176 2644
rect 13228 2592 13234 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 15105 2635 15163 2641
rect 15105 2632 15117 2635
rect 13320 2604 15117 2632
rect 13320 2592 13326 2604
rect 15105 2601 15117 2604
rect 15151 2601 15163 2635
rect 15105 2595 15163 2601
rect 15381 2635 15439 2641
rect 15381 2601 15393 2635
rect 15427 2632 15439 2635
rect 16942 2632 16948 2644
rect 15427 2604 16948 2632
rect 15427 2601 15439 2604
rect 15381 2595 15439 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 18322 2592 18328 2644
rect 18380 2592 18386 2644
rect 18877 2635 18935 2641
rect 18877 2601 18889 2635
rect 18923 2632 18935 2635
rect 19978 2632 19984 2644
rect 18923 2604 19984 2632
rect 18923 2601 18935 2604
rect 18877 2595 18935 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 23198 2632 23204 2644
rect 20864 2604 23204 2632
rect 20864 2592 20870 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 24394 2592 24400 2644
rect 24452 2632 24458 2644
rect 25133 2635 25191 2641
rect 25133 2632 25145 2635
rect 24452 2604 25145 2632
rect 24452 2592 24458 2604
rect 25133 2601 25145 2604
rect 25179 2601 25191 2635
rect 25133 2595 25191 2601
rect 25498 2592 25504 2644
rect 25556 2632 25562 2644
rect 26237 2635 26295 2641
rect 26237 2632 26249 2635
rect 25556 2604 26249 2632
rect 25556 2592 25562 2604
rect 26237 2601 26249 2604
rect 26283 2601 26295 2635
rect 26237 2595 26295 2601
rect 26510 2592 26516 2644
rect 26568 2632 26574 2644
rect 26789 2635 26847 2641
rect 26789 2632 26801 2635
rect 26568 2604 26801 2632
rect 26568 2592 26574 2604
rect 26789 2601 26801 2604
rect 26835 2601 26847 2635
rect 26789 2595 26847 2601
rect 26878 2592 26884 2644
rect 26936 2632 26942 2644
rect 27709 2635 27767 2641
rect 27709 2632 27721 2635
rect 26936 2604 27721 2632
rect 26936 2592 26942 2604
rect 27709 2601 27721 2604
rect 27755 2601 27767 2635
rect 27709 2595 27767 2601
rect 28626 2592 28632 2644
rect 28684 2632 28690 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 28684 2604 29745 2632
rect 28684 2592 28690 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 29733 2595 29791 2601
rect 30837 2635 30895 2641
rect 30837 2601 30849 2635
rect 30883 2601 30895 2635
rect 30837 2595 30895 2601
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2533 10379 2567
rect 10321 2527 10379 2533
rect 11054 2524 11060 2576
rect 11112 2524 11118 2576
rect 11330 2524 11336 2576
rect 11388 2524 11394 2576
rect 11977 2567 12035 2573
rect 11977 2533 11989 2567
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 12253 2567 12311 2573
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 14458 2564 14464 2576
rect 12299 2536 14464 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 11238 2496 11244 2508
rect 6840 2468 11244 2496
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 5626 2428 5632 2440
rect 5491 2400 5632 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 5902 2428 5908 2440
rect 5767 2400 5908 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6270 2428 6276 2440
rect 6043 2400 6276 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 6840 2360 6868 2468
rect 11238 2456 11244 2468
rect 11296 2456 11302 2508
rect 11992 2496 12020 2527
rect 14458 2524 14464 2536
rect 14516 2524 14522 2576
rect 14553 2567 14611 2573
rect 14553 2533 14565 2567
rect 14599 2564 14611 2567
rect 14642 2564 14648 2576
rect 14599 2536 14648 2564
rect 14599 2533 14611 2536
rect 14553 2527 14611 2533
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 14752 2536 15424 2564
rect 14752 2496 14780 2536
rect 15396 2508 15424 2536
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 16448 2536 28028 2564
rect 16448 2524 16454 2536
rect 15102 2496 15108 2508
rect 11992 2468 14780 2496
rect 14936 2468 15108 2496
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7466 2388 7472 2440
rect 7524 2388 7530 2440
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 8018 2388 8024 2440
rect 8076 2388 8082 2440
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 8754 2388 8760 2440
rect 8812 2388 8818 2440
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9398 2428 9404 2440
rect 9263 2400 9404 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 6196 2332 6868 2360
rect 7668 2332 8432 2360
rect 5626 2252 5632 2304
rect 5684 2252 5690 2304
rect 6196 2301 6224 2332
rect 6181 2295 6239 2301
rect 6181 2261 6193 2295
rect 6227 2261 6239 2295
rect 6181 2255 6239 2261
rect 6825 2295 6883 2301
rect 6825 2261 6837 2295
rect 6871 2292 6883 2295
rect 7098 2292 7104 2304
rect 6871 2264 7104 2292
rect 6871 2261 6883 2264
rect 6825 2255 6883 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7374 2252 7380 2304
rect 7432 2252 7438 2304
rect 7668 2301 7696 2332
rect 8404 2304 8432 2332
rect 7653 2295 7711 2301
rect 7653 2261 7665 2295
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7926 2252 7932 2304
rect 7984 2252 7990 2304
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 8496 2301 8524 2388
rect 8772 2301 8800 2388
rect 8956 2360 8984 2391
rect 9398 2388 9404 2400
rect 9456 2388 9462 2440
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9674 2428 9680 2440
rect 9539 2400 9680 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10410 2428 10416 2440
rect 10091 2400 10416 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 9306 2360 9312 2372
rect 8956 2332 9312 2360
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 9784 2360 9812 2391
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10502 2388 10508 2440
rect 10560 2388 10566 2440
rect 10686 2388 10692 2440
rect 10744 2388 10750 2440
rect 10778 2388 10784 2440
rect 10836 2388 10842 2440
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11054 2428 11060 2440
rect 10919 2400 11060 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 11422 2428 11428 2440
rect 11195 2400 11428 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11514 2388 11520 2440
rect 11572 2388 11578 2440
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2428 11851 2431
rect 11974 2428 11980 2440
rect 11839 2400 11980 2428
rect 11839 2397 11851 2400
rect 11793 2391 11851 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 12526 2428 12532 2440
rect 12391 2400 12532 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 10134 2360 10140 2372
rect 9784 2332 10140 2360
rect 10134 2320 10140 2332
rect 10192 2320 10198 2372
rect 10704 2360 10732 2388
rect 10244 2332 10732 2360
rect 8481 2295 8539 2301
rect 8481 2261 8493 2295
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 8757 2295 8815 2301
rect 8757 2261 8769 2295
rect 8803 2261 8815 2295
rect 8757 2255 8815 2261
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 9214 2292 9220 2304
rect 9171 2264 9220 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9401 2295 9459 2301
rect 9401 2261 9413 2295
rect 9447 2292 9459 2295
rect 9490 2292 9496 2304
rect 9447 2264 9496 2292
rect 9447 2261 9459 2264
rect 9401 2255 9459 2261
rect 9490 2252 9496 2264
rect 9548 2252 9554 2304
rect 10244 2301 10272 2332
rect 11882 2320 11888 2372
rect 11940 2360 11946 2372
rect 12084 2360 12112 2391
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 12802 2428 12808 2440
rect 12667 2400 12808 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 12802 2388 12808 2400
rect 12860 2388 12866 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 13170 2428 13176 2440
rect 12943 2400 13176 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 13354 2388 13360 2440
rect 13412 2388 13418 2440
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 13630 2428 13636 2440
rect 13495 2400 13636 2428
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 13722 2388 13728 2440
rect 13780 2388 13786 2440
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2428 14519 2431
rect 14642 2428 14648 2440
rect 14507 2400 14648 2428
rect 14507 2397 14519 2400
rect 14461 2391 14519 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 14734 2388 14740 2440
rect 14792 2388 14798 2440
rect 13280 2360 13308 2388
rect 14550 2360 14556 2372
rect 11940 2332 12112 2360
rect 12820 2332 13308 2360
rect 13648 2332 14556 2360
rect 11940 2320 11946 2332
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2261 10287 2295
rect 10229 2255 10287 2261
rect 10594 2252 10600 2304
rect 10652 2252 10658 2304
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 12526 2252 12532 2304
rect 12584 2252 12590 2304
rect 12820 2301 12848 2332
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 13078 2252 13084 2304
rect 13136 2252 13142 2304
rect 13648 2301 13676 2332
rect 14550 2320 14556 2332
rect 14608 2320 14614 2372
rect 14936 2360 14964 2468
rect 15102 2456 15108 2468
rect 15160 2456 15166 2508
rect 15378 2456 15384 2508
rect 15436 2456 15442 2508
rect 15930 2456 15936 2508
rect 15988 2456 15994 2508
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 16945 2499 17003 2505
rect 16945 2496 16957 2499
rect 16908 2468 16957 2496
rect 16908 2456 16914 2468
rect 16945 2465 16957 2468
rect 16991 2465 17003 2499
rect 16945 2459 17003 2465
rect 17957 2499 18015 2505
rect 17957 2465 17969 2499
rect 18003 2496 18015 2499
rect 18046 2496 18052 2508
rect 18003 2468 18052 2496
rect 18003 2465 18015 2468
rect 17957 2459 18015 2465
rect 18046 2456 18052 2468
rect 18104 2456 18110 2508
rect 19702 2496 19708 2508
rect 18248 2468 19708 2496
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15194 2428 15200 2440
rect 15059 2400 15200 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2428 15715 2431
rect 15838 2428 15844 2440
rect 15703 2400 15844 2428
rect 15703 2397 15715 2400
rect 15657 2391 15715 2397
rect 14844 2332 14964 2360
rect 15580 2360 15608 2391
rect 15838 2388 15844 2400
rect 15896 2388 15902 2440
rect 16390 2388 16396 2440
rect 16448 2428 16454 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16448 2400 16681 2428
rect 16448 2388 16454 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17126 2388 17132 2440
rect 17184 2428 17190 2440
rect 18248 2437 18276 2468
rect 19702 2456 19708 2468
rect 19760 2456 19766 2508
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2496 19947 2499
rect 20346 2496 20352 2508
rect 19935 2468 20352 2496
rect 19935 2465 19947 2468
rect 19889 2459 19947 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 20441 2499 20499 2505
rect 20441 2465 20453 2499
rect 20487 2496 20499 2499
rect 20714 2496 20720 2508
rect 20487 2468 20720 2496
rect 20487 2465 20499 2468
rect 20441 2459 20499 2465
rect 20714 2456 20720 2468
rect 20772 2456 20778 2508
rect 21818 2456 21824 2508
rect 21876 2496 21882 2508
rect 21876 2468 23336 2496
rect 21876 2456 21882 2468
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17184 2400 17785 2428
rect 17184 2388 17190 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2397 18291 2431
rect 18233 2391 18291 2397
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 18656 2400 18797 2428
rect 18656 2388 18662 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 18874 2388 18880 2440
rect 18932 2428 18938 2440
rect 19061 2431 19119 2437
rect 19061 2428 19073 2431
rect 18932 2400 19073 2428
rect 18932 2388 18938 2400
rect 19061 2397 19073 2400
rect 19107 2397 19119 2431
rect 19061 2391 19119 2397
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19392 2400 19441 2428
rect 19392 2388 19398 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 19794 2428 19800 2440
rect 19659 2400 19800 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 19794 2388 19800 2400
rect 19852 2388 19858 2440
rect 21174 2388 21180 2440
rect 21232 2428 21238 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 21232 2400 21281 2428
rect 21232 2388 21238 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21542 2388 21548 2440
rect 21600 2428 21606 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21600 2400 22017 2428
rect 21600 2388 21606 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22094 2388 22100 2440
rect 22152 2428 22158 2440
rect 23308 2437 23336 2468
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 22152 2400 22201 2428
rect 22152 2388 22158 2400
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 23293 2431 23351 2437
rect 22189 2391 22247 2397
rect 22296 2400 22876 2428
rect 16850 2360 16856 2372
rect 15580 2332 16856 2360
rect 13633 2295 13691 2301
rect 13633 2261 13645 2295
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 14182 2292 14188 2304
rect 13955 2264 14188 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 14274 2252 14280 2304
rect 14332 2252 14338 2304
rect 14844 2301 14872 2332
rect 16850 2320 16856 2332
rect 16908 2320 16914 2372
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 18616 2332 20177 2360
rect 14829 2295 14887 2301
rect 14829 2261 14841 2295
rect 14875 2261 14887 2295
rect 14829 2255 14887 2261
rect 18046 2252 18052 2304
rect 18104 2252 18110 2304
rect 18616 2301 18644 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20165 2323 20223 2329
rect 20717 2363 20775 2369
rect 20717 2329 20729 2363
rect 20763 2329 20775 2363
rect 20717 2323 20775 2329
rect 21085 2363 21143 2369
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21450 2360 21456 2372
rect 21131 2332 21456 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2261 18659 2295
rect 18601 2255 18659 2261
rect 19245 2295 19303 2301
rect 19245 2261 19257 2295
rect 19291 2292 19303 2295
rect 20732 2292 20760 2323
rect 21450 2320 21456 2332
rect 21508 2320 21514 2372
rect 21634 2320 21640 2372
rect 21692 2320 21698 2372
rect 22296 2360 22324 2400
rect 21836 2332 22324 2360
rect 21836 2301 21864 2332
rect 22370 2320 22376 2372
rect 22428 2360 22434 2372
rect 22557 2363 22615 2369
rect 22557 2360 22569 2363
rect 22428 2332 22569 2360
rect 22428 2320 22434 2332
rect 22557 2329 22569 2332
rect 22603 2329 22615 2363
rect 22557 2323 22615 2329
rect 22741 2363 22799 2369
rect 22741 2329 22753 2363
rect 22787 2329 22799 2363
rect 22848 2360 22876 2400
rect 23293 2397 23305 2431
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 23566 2388 23572 2440
rect 23624 2428 23630 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23624 2400 23857 2428
rect 23624 2388 23630 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 24854 2388 24860 2440
rect 24912 2428 24918 2440
rect 25041 2431 25099 2437
rect 25041 2428 25053 2431
rect 24912 2400 25053 2428
rect 24912 2388 24918 2400
rect 25041 2397 25053 2400
rect 25087 2397 25099 2431
rect 25041 2391 25099 2397
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25593 2431 25651 2437
rect 25593 2428 25605 2431
rect 25464 2400 25605 2428
rect 25464 2388 25470 2400
rect 25593 2397 25605 2400
rect 25639 2397 25651 2431
rect 25593 2391 25651 2397
rect 26602 2388 26608 2440
rect 26660 2388 26666 2440
rect 27617 2431 27675 2437
rect 27617 2397 27629 2431
rect 27663 2428 27675 2431
rect 27890 2428 27896 2440
rect 27663 2400 27896 2428
rect 27663 2397 27675 2400
rect 27617 2391 27675 2397
rect 27890 2388 27896 2400
rect 27948 2388 27954 2440
rect 24489 2363 24547 2369
rect 24489 2360 24501 2363
rect 22848 2332 24501 2360
rect 22741 2323 22799 2329
rect 24489 2329 24501 2332
rect 24535 2329 24547 2363
rect 25240 2360 25268 2388
rect 26145 2363 26203 2369
rect 26145 2360 26157 2363
rect 25240 2332 26157 2360
rect 24489 2323 24547 2329
rect 26145 2329 26157 2332
rect 26191 2329 26203 2363
rect 26145 2323 26203 2329
rect 19291 2264 20760 2292
rect 21821 2295 21879 2301
rect 19291 2261 19303 2264
rect 19245 2255 19303 2261
rect 21821 2261 21833 2295
rect 21867 2261 21879 2295
rect 21821 2255 21879 2261
rect 21910 2252 21916 2304
rect 21968 2292 21974 2304
rect 22756 2292 22784 2323
rect 26326 2320 26332 2372
rect 26384 2360 26390 2372
rect 26384 2332 26924 2360
rect 26384 2320 26390 2332
rect 21968 2264 22784 2292
rect 21968 2252 21974 2264
rect 22830 2252 22836 2304
rect 22888 2252 22894 2304
rect 23566 2252 23572 2304
rect 23624 2252 23630 2304
rect 23658 2252 23664 2304
rect 23716 2292 23722 2304
rect 23937 2295 23995 2301
rect 23937 2292 23949 2295
rect 23716 2264 23949 2292
rect 23716 2252 23722 2264
rect 23937 2261 23949 2264
rect 23983 2261 23995 2295
rect 23937 2255 23995 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 24581 2295 24639 2301
rect 24581 2292 24593 2295
rect 24084 2264 24593 2292
rect 24084 2252 24090 2264
rect 24581 2261 24593 2264
rect 24627 2261 24639 2295
rect 24581 2255 24639 2261
rect 24946 2252 24952 2304
rect 25004 2292 25010 2304
rect 25685 2295 25743 2301
rect 25685 2292 25697 2295
rect 25004 2264 25697 2292
rect 25004 2252 25010 2264
rect 25685 2261 25697 2264
rect 25731 2261 25743 2295
rect 26896 2292 26924 2332
rect 27062 2320 27068 2372
rect 27120 2320 27126 2372
rect 27430 2320 27436 2372
rect 27488 2360 27494 2372
rect 28000 2360 28028 2536
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 30377 2567 30435 2573
rect 30377 2564 30389 2567
rect 28960 2536 30389 2564
rect 28960 2524 28966 2536
rect 30377 2533 30389 2536
rect 30423 2533 30435 2567
rect 30377 2527 30435 2533
rect 28074 2456 28080 2508
rect 28132 2496 28138 2508
rect 28997 2499 29055 2505
rect 28997 2496 29009 2499
rect 28132 2468 29009 2496
rect 28132 2456 28138 2468
rect 28997 2465 29009 2468
rect 29043 2465 29055 2499
rect 28997 2459 29055 2465
rect 29546 2456 29552 2508
rect 29604 2496 29610 2508
rect 30852 2496 30880 2595
rect 31110 2592 31116 2644
rect 31168 2632 31174 2644
rect 32309 2635 32367 2641
rect 32309 2632 32321 2635
rect 31168 2604 32321 2632
rect 31168 2592 31174 2604
rect 32309 2601 32321 2604
rect 32355 2601 32367 2635
rect 32309 2595 32367 2601
rect 32950 2592 32956 2644
rect 33008 2592 33014 2644
rect 33502 2592 33508 2644
rect 33560 2632 33566 2644
rect 34885 2635 34943 2641
rect 34885 2632 34897 2635
rect 33560 2604 34897 2632
rect 33560 2592 33566 2604
rect 34885 2601 34897 2604
rect 34931 2601 34943 2635
rect 34885 2595 34943 2601
rect 35894 2592 35900 2644
rect 35952 2632 35958 2644
rect 36081 2635 36139 2641
rect 36081 2632 36093 2635
rect 35952 2604 36093 2632
rect 35952 2592 35958 2604
rect 36081 2601 36093 2604
rect 36127 2601 36139 2635
rect 36081 2595 36139 2601
rect 36630 2592 36636 2644
rect 36688 2592 36694 2644
rect 37090 2592 37096 2644
rect 37148 2592 37154 2644
rect 37458 2592 37464 2644
rect 37516 2592 37522 2644
rect 37826 2592 37832 2644
rect 37884 2632 37890 2644
rect 38013 2635 38071 2641
rect 38013 2632 38025 2635
rect 37884 2604 38025 2632
rect 37884 2592 37890 2604
rect 38013 2601 38025 2604
rect 38059 2601 38071 2635
rect 38013 2595 38071 2601
rect 39022 2592 39028 2644
rect 39080 2632 39086 2644
rect 39117 2635 39175 2641
rect 39117 2632 39129 2635
rect 39080 2604 39129 2632
rect 39080 2592 39086 2604
rect 39117 2601 39129 2604
rect 39163 2601 39175 2635
rect 39117 2595 39175 2601
rect 31757 2567 31815 2573
rect 31757 2564 31769 2567
rect 29604 2468 30880 2496
rect 30944 2536 31769 2564
rect 29604 2456 29610 2468
rect 28169 2431 28227 2437
rect 28169 2397 28181 2431
rect 28215 2428 28227 2431
rect 28534 2428 28540 2440
rect 28215 2400 28540 2428
rect 28215 2397 28227 2400
rect 28169 2391 28227 2397
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 28718 2388 28724 2440
rect 28776 2388 28782 2440
rect 29086 2388 29092 2440
rect 29144 2388 29150 2440
rect 29362 2388 29368 2440
rect 29420 2388 29426 2440
rect 29454 2388 29460 2440
rect 29512 2428 29518 2440
rect 29641 2431 29699 2437
rect 29641 2428 29653 2431
rect 29512 2400 29653 2428
rect 29512 2388 29518 2400
rect 29641 2397 29653 2400
rect 29687 2397 29699 2431
rect 29641 2391 29699 2397
rect 30742 2388 30748 2440
rect 30800 2388 30806 2440
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 30944 2428 30972 2536
rect 31757 2533 31769 2536
rect 31803 2533 31815 2567
rect 32968 2564 32996 2592
rect 34333 2567 34391 2573
rect 34333 2564 34345 2567
rect 32968 2536 34345 2564
rect 31757 2527 31815 2533
rect 34333 2533 34345 2536
rect 34379 2533 34391 2567
rect 34333 2527 34391 2533
rect 34422 2524 34428 2576
rect 34480 2564 34486 2576
rect 35989 2567 36047 2573
rect 35989 2564 36001 2567
rect 34480 2536 36001 2564
rect 34480 2524 34486 2536
rect 35989 2533 36001 2536
rect 36035 2533 36047 2567
rect 35989 2527 36047 2533
rect 36998 2524 37004 2576
rect 37056 2564 37062 2576
rect 37056 2536 37872 2564
rect 37056 2524 37062 2536
rect 31662 2456 31668 2508
rect 31720 2496 31726 2508
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 31720 2468 33609 2496
rect 31720 2456 31726 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 33597 2459 33655 2465
rect 35250 2456 35256 2508
rect 35308 2496 35314 2508
rect 35308 2468 36308 2496
rect 35308 2456 35314 2468
rect 30892 2400 30972 2428
rect 30892 2388 30898 2400
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 31444 2400 31754 2428
rect 31444 2388 31450 2400
rect 28994 2360 29000 2372
rect 27488 2332 27844 2360
rect 28000 2332 29000 2360
rect 27488 2320 27494 2332
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26896 2264 27169 2292
rect 25685 2255 25743 2261
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27816 2292 27844 2332
rect 28994 2320 29000 2332
rect 29052 2320 29058 2372
rect 29104 2360 29132 2388
rect 30193 2363 30251 2369
rect 30193 2360 30205 2363
rect 29104 2332 30205 2360
rect 30193 2329 30205 2332
rect 30239 2329 30251 2363
rect 30193 2323 30251 2329
rect 30374 2320 30380 2372
rect 30432 2360 30438 2372
rect 31297 2363 31355 2369
rect 31297 2360 31309 2363
rect 30432 2332 31309 2360
rect 30432 2320 30438 2332
rect 31297 2329 31309 2332
rect 31343 2329 31355 2363
rect 31726 2360 31754 2400
rect 31938 2388 31944 2440
rect 31996 2388 32002 2440
rect 32140 2400 32352 2428
rect 32140 2360 32168 2400
rect 31726 2332 32168 2360
rect 31297 2323 31355 2329
rect 32214 2320 32220 2372
rect 32272 2320 32278 2372
rect 32324 2360 32352 2400
rect 32674 2388 32680 2440
rect 32732 2428 32738 2440
rect 32769 2431 32827 2437
rect 32769 2428 32781 2431
rect 32732 2400 32781 2428
rect 32732 2388 32738 2400
rect 32769 2397 32781 2400
rect 32815 2397 32827 2431
rect 32769 2391 32827 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32916 2400 33088 2428
rect 32916 2388 32922 2400
rect 33060 2360 33088 2400
rect 33134 2388 33140 2440
rect 33192 2428 33198 2440
rect 33321 2431 33379 2437
rect 33321 2428 33333 2431
rect 33192 2400 33333 2428
rect 33192 2388 33198 2400
rect 33321 2397 33333 2400
rect 33367 2397 33379 2431
rect 33321 2391 33379 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 36280 2437 36308 2468
rect 36538 2456 36544 2508
rect 36596 2496 36602 2508
rect 36596 2468 37320 2496
rect 36596 2456 36602 2468
rect 34517 2431 34575 2437
rect 34517 2428 34529 2431
rect 33468 2400 34529 2428
rect 33468 2388 33474 2400
rect 34517 2397 34529 2400
rect 34563 2397 34575 2431
rect 35805 2431 35863 2437
rect 35805 2428 35817 2431
rect 34517 2391 34575 2397
rect 34624 2400 35817 2428
rect 33873 2363 33931 2369
rect 33873 2360 33885 2363
rect 32324 2332 32904 2360
rect 33060 2332 33885 2360
rect 28261 2295 28319 2301
rect 28261 2292 28273 2295
rect 27816 2264 28273 2292
rect 27157 2255 27215 2261
rect 28261 2261 28273 2264
rect 28307 2261 28319 2295
rect 28261 2255 28319 2261
rect 29181 2295 29239 2301
rect 29181 2261 29193 2295
rect 29227 2292 29239 2295
rect 29638 2292 29644 2304
rect 29227 2264 29644 2292
rect 29227 2261 29239 2264
rect 29181 2255 29239 2261
rect 29638 2252 29644 2264
rect 29696 2252 29702 2304
rect 30098 2252 30104 2304
rect 30156 2292 30162 2304
rect 32876 2301 32904 2332
rect 33873 2329 33885 2332
rect 33919 2329 33931 2363
rect 33873 2323 33931 2329
rect 34330 2320 34336 2372
rect 34388 2360 34394 2372
rect 34624 2360 34652 2400
rect 35805 2397 35817 2400
rect 35851 2397 35863 2431
rect 35805 2391 35863 2397
rect 36265 2431 36323 2437
rect 36265 2397 36277 2431
rect 36311 2397 36323 2431
rect 36265 2391 36323 2397
rect 36357 2431 36415 2437
rect 36357 2397 36369 2431
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 34388 2332 34652 2360
rect 34388 2320 34394 2332
rect 34790 2320 34796 2372
rect 34848 2320 34854 2372
rect 35342 2320 35348 2372
rect 35400 2320 35406 2372
rect 35894 2320 35900 2372
rect 35952 2360 35958 2372
rect 36372 2360 36400 2391
rect 36814 2388 36820 2440
rect 36872 2388 36878 2440
rect 37292 2437 37320 2468
rect 37844 2437 37872 2536
rect 38102 2524 38108 2576
rect 38160 2564 38166 2576
rect 38289 2567 38347 2573
rect 38289 2564 38301 2567
rect 38160 2536 38301 2564
rect 38160 2524 38166 2536
rect 38289 2533 38301 2536
rect 38335 2533 38347 2567
rect 38289 2527 38347 2533
rect 38838 2524 38844 2576
rect 38896 2564 38902 2576
rect 38896 2536 39344 2564
rect 38896 2524 38902 2536
rect 37918 2456 37924 2508
rect 37976 2496 37982 2508
rect 37976 2468 38424 2496
rect 37976 2456 37982 2468
rect 38396 2437 38424 2468
rect 38470 2456 38476 2508
rect 38528 2496 38534 2508
rect 38528 2468 38976 2496
rect 38528 2456 38534 2468
rect 38948 2437 38976 2468
rect 36909 2431 36967 2437
rect 36909 2397 36921 2431
rect 36955 2397 36967 2431
rect 36909 2391 36967 2397
rect 37277 2431 37335 2437
rect 37277 2397 37289 2431
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 37829 2431 37887 2437
rect 37829 2397 37841 2431
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 38105 2431 38163 2437
rect 38105 2397 38117 2431
rect 38151 2397 38163 2431
rect 38105 2391 38163 2397
rect 38381 2431 38439 2437
rect 38381 2397 38393 2431
rect 38427 2397 38439 2431
rect 38381 2391 38439 2397
rect 38657 2431 38715 2437
rect 38657 2397 38669 2431
rect 38703 2397 38715 2431
rect 38657 2391 38715 2397
rect 38933 2431 38991 2437
rect 38933 2397 38945 2431
rect 38979 2397 38991 2431
rect 39209 2431 39267 2437
rect 39209 2428 39221 2431
rect 38933 2391 38991 2397
rect 39040 2400 39221 2428
rect 36924 2360 36952 2391
rect 37568 2360 37596 2391
rect 35952 2332 36400 2360
rect 36464 2332 36952 2360
rect 37292 2332 37596 2360
rect 35952 2320 35958 2332
rect 31389 2295 31447 2301
rect 31389 2292 31401 2295
rect 30156 2264 31401 2292
rect 30156 2252 30162 2264
rect 31389 2261 31401 2264
rect 31435 2261 31447 2295
rect 31389 2255 31447 2261
rect 32861 2295 32919 2301
rect 32861 2261 32873 2295
rect 32907 2261 32919 2295
rect 32861 2255 32919 2261
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 33965 2295 34023 2301
rect 33965 2292 33977 2295
rect 33192 2264 33977 2292
rect 33192 2252 33198 2264
rect 33965 2261 33977 2264
rect 34011 2261 34023 2295
rect 33965 2255 34023 2261
rect 35434 2252 35440 2304
rect 35492 2252 35498 2304
rect 36078 2252 36084 2304
rect 36136 2292 36142 2304
rect 36464 2292 36492 2332
rect 36136 2264 36492 2292
rect 36136 2252 36142 2264
rect 36538 2252 36544 2304
rect 36596 2252 36602 2304
rect 36630 2252 36636 2304
rect 36688 2292 36694 2304
rect 37292 2292 37320 2332
rect 37642 2320 37648 2372
rect 37700 2360 37706 2372
rect 38120 2360 38148 2391
rect 37700 2332 38148 2360
rect 37700 2320 37706 2332
rect 38194 2320 38200 2372
rect 38252 2360 38258 2372
rect 38672 2360 38700 2391
rect 38252 2332 38700 2360
rect 38252 2320 38258 2332
rect 38746 2320 38752 2372
rect 38804 2360 38810 2372
rect 39040 2360 39068 2400
rect 39209 2397 39221 2400
rect 39255 2397 39267 2431
rect 39316 2428 39344 2536
rect 39390 2456 39396 2508
rect 39448 2496 39454 2508
rect 39448 2468 39988 2496
rect 39448 2456 39454 2468
rect 39485 2431 39543 2437
rect 39485 2428 39497 2431
rect 39316 2400 39497 2428
rect 39209 2391 39267 2397
rect 39485 2397 39497 2400
rect 39531 2397 39543 2431
rect 39485 2391 39543 2397
rect 39853 2431 39911 2437
rect 39853 2397 39865 2431
rect 39899 2397 39911 2431
rect 39960 2428 39988 2468
rect 40034 2456 40040 2508
rect 40092 2496 40098 2508
rect 40092 2468 40724 2496
rect 40092 2456 40098 2468
rect 40129 2431 40187 2437
rect 40129 2428 40141 2431
rect 39960 2400 40141 2428
rect 39853 2391 39911 2397
rect 40129 2397 40141 2400
rect 40175 2397 40187 2431
rect 40129 2391 40187 2397
rect 38804 2332 39068 2360
rect 38804 2320 38810 2332
rect 39114 2320 39120 2372
rect 39172 2360 39178 2372
rect 39868 2360 39896 2391
rect 40402 2388 40408 2440
rect 40460 2388 40466 2440
rect 40696 2437 40724 2468
rect 40681 2431 40739 2437
rect 40681 2397 40693 2431
rect 40727 2397 40739 2431
rect 40681 2391 40739 2397
rect 40957 2431 41015 2437
rect 40957 2397 40969 2431
rect 41003 2397 41015 2431
rect 40957 2391 41015 2397
rect 39172 2332 39896 2360
rect 39172 2320 39178 2332
rect 40218 2320 40224 2372
rect 40276 2360 40282 2372
rect 40972 2360 41000 2391
rect 40276 2332 41000 2360
rect 40276 2320 40282 2332
rect 36688 2264 37320 2292
rect 36688 2252 36694 2264
rect 37734 2252 37740 2304
rect 37792 2252 37798 2304
rect 38378 2252 38384 2304
rect 38436 2292 38442 2304
rect 38565 2295 38623 2301
rect 38565 2292 38577 2295
rect 38436 2264 38577 2292
rect 38436 2252 38442 2264
rect 38565 2261 38577 2264
rect 38611 2261 38623 2295
rect 38565 2255 38623 2261
rect 38841 2295 38899 2301
rect 38841 2261 38853 2295
rect 38887 2292 38899 2295
rect 39022 2292 39028 2304
rect 38887 2264 39028 2292
rect 38887 2261 38899 2264
rect 38841 2255 38899 2261
rect 39022 2252 39028 2264
rect 39080 2252 39086 2304
rect 39298 2252 39304 2304
rect 39356 2292 39362 2304
rect 39393 2295 39451 2301
rect 39393 2292 39405 2295
rect 39356 2264 39405 2292
rect 39356 2252 39362 2264
rect 39393 2261 39405 2264
rect 39439 2261 39451 2295
rect 39393 2255 39451 2261
rect 39666 2252 39672 2304
rect 39724 2252 39730 2304
rect 40034 2252 40040 2304
rect 40092 2252 40098 2304
rect 40310 2252 40316 2304
rect 40368 2252 40374 2304
rect 40589 2295 40647 2301
rect 40589 2261 40601 2295
rect 40635 2292 40647 2295
rect 40678 2292 40684 2304
rect 40635 2264 40684 2292
rect 40635 2261 40647 2264
rect 40589 2255 40647 2261
rect 40678 2252 40684 2264
rect 40736 2252 40742 2304
rect 40862 2252 40868 2304
rect 40920 2252 40926 2304
rect 41138 2252 41144 2304
rect 41196 2252 41202 2304
rect 1104 2202 45051 2224
rect 1104 2150 11896 2202
rect 11948 2150 11960 2202
rect 12012 2150 12024 2202
rect 12076 2150 12088 2202
rect 12140 2150 12152 2202
rect 12204 2150 22843 2202
rect 22895 2150 22907 2202
rect 22959 2150 22971 2202
rect 23023 2150 23035 2202
rect 23087 2150 23099 2202
rect 23151 2150 33790 2202
rect 33842 2150 33854 2202
rect 33906 2150 33918 2202
rect 33970 2150 33982 2202
rect 34034 2150 34046 2202
rect 34098 2150 44737 2202
rect 44789 2150 44801 2202
rect 44853 2150 44865 2202
rect 44917 2150 44929 2202
rect 44981 2150 44993 2202
rect 45045 2150 45051 2202
rect 1104 2128 45051 2150
rect 8202 2048 8208 2100
rect 8260 2048 8266 2100
rect 8386 2048 8392 2100
rect 8444 2088 8450 2100
rect 10870 2088 10876 2100
rect 8444 2060 10876 2088
rect 8444 2048 8450 2060
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 14458 2048 14464 2100
rect 14516 2048 14522 2100
rect 15286 2048 15292 2100
rect 15344 2048 15350 2100
rect 15378 2048 15384 2100
rect 15436 2088 15442 2100
rect 15436 2060 27292 2088
rect 15436 2048 15442 2060
rect 8220 1748 8248 2048
rect 14476 1952 14504 2048
rect 15304 2020 15332 2048
rect 27154 2020 27160 2032
rect 15304 1992 27160 2020
rect 27154 1980 27160 1992
rect 27212 1980 27218 2032
rect 19150 1952 19156 1964
rect 14476 1924 19156 1952
rect 19150 1912 19156 1924
rect 19208 1912 19214 1964
rect 19886 1912 19892 1964
rect 19944 1912 19950 1964
rect 20990 1912 20996 1964
rect 21048 1952 21054 1964
rect 27062 1952 27068 1964
rect 21048 1924 27068 1952
rect 21048 1912 21054 1924
rect 27062 1912 27068 1924
rect 27120 1912 27126 1964
rect 27264 1952 27292 2060
rect 28534 2048 28540 2100
rect 28592 2088 28598 2100
rect 28592 2060 29592 2088
rect 28592 2048 28598 2060
rect 27338 1980 27344 2032
rect 27396 2020 27402 2032
rect 28994 2020 29000 2032
rect 27396 1992 29000 2020
rect 27396 1980 27402 1992
rect 28994 1980 29000 1992
rect 29052 1980 29058 2032
rect 29362 1980 29368 2032
rect 29420 1980 29426 2032
rect 29564 2020 29592 2060
rect 29638 2048 29644 2100
rect 29696 2088 29702 2100
rect 34790 2088 34796 2100
rect 29696 2060 34796 2088
rect 29696 2048 29702 2060
rect 34790 2048 34796 2060
rect 34848 2048 34854 2100
rect 35342 2048 35348 2100
rect 35400 2048 35406 2100
rect 39022 2048 39028 2100
rect 39080 2048 39086 2100
rect 30834 2020 30840 2032
rect 29564 1992 30840 2020
rect 30834 1980 30840 1992
rect 30892 1980 30898 2032
rect 35360 2020 35388 2048
rect 30944 1992 35388 2020
rect 29380 1952 29408 1980
rect 27264 1924 29408 1952
rect 30282 1912 30288 1964
rect 30340 1952 30346 1964
rect 30944 1952 30972 1992
rect 30340 1924 30972 1952
rect 31588 1924 31800 1952
rect 30340 1912 30346 1924
rect 14642 1844 14648 1896
rect 14700 1884 14706 1896
rect 14700 1856 16574 1884
rect 14700 1844 14706 1856
rect 9214 1776 9220 1828
rect 9272 1816 9278 1828
rect 15562 1816 15568 1828
rect 9272 1788 15568 1816
rect 9272 1776 9278 1788
rect 15562 1776 15568 1788
rect 15620 1776 15626 1828
rect 16546 1816 16574 1856
rect 18046 1844 18052 1896
rect 18104 1884 18110 1896
rect 19904 1884 19932 1912
rect 18104 1856 19932 1884
rect 18104 1844 18110 1856
rect 23198 1844 23204 1896
rect 23256 1884 23262 1896
rect 31588 1884 31616 1924
rect 23256 1856 31616 1884
rect 31772 1884 31800 1924
rect 32122 1912 32128 1964
rect 32180 1952 32186 1964
rect 32180 1924 38654 1952
rect 32180 1912 32186 1924
rect 38626 1884 38654 1924
rect 39040 1884 39068 2048
rect 39298 1912 39304 1964
rect 39356 1912 39362 1964
rect 31772 1856 35296 1884
rect 38626 1856 39068 1884
rect 23256 1844 23262 1856
rect 35268 1816 35296 1856
rect 39316 1816 39344 1912
rect 16546 1788 31524 1816
rect 35268 1788 39344 1816
rect 8220 1720 11652 1748
rect 5626 1640 5632 1692
rect 5684 1680 5690 1692
rect 5684 1652 6914 1680
rect 5684 1640 5690 1652
rect 6886 1408 6914 1652
rect 7374 1640 7380 1692
rect 7432 1680 7438 1692
rect 10318 1680 10324 1692
rect 7432 1652 10324 1680
rect 7432 1640 7438 1652
rect 10318 1640 10324 1652
rect 10376 1640 10382 1692
rect 10594 1640 10600 1692
rect 10652 1640 10658 1692
rect 10612 1476 10640 1640
rect 11624 1544 11652 1720
rect 12526 1708 12532 1760
rect 12584 1748 12590 1760
rect 31202 1748 31208 1760
rect 12584 1720 31208 1748
rect 12584 1708 12590 1720
rect 31202 1708 31208 1720
rect 31260 1708 31266 1760
rect 13354 1640 13360 1692
rect 13412 1680 13418 1692
rect 13412 1652 16574 1680
rect 13412 1640 13418 1652
rect 11698 1572 11704 1624
rect 11756 1612 11762 1624
rect 15194 1612 15200 1624
rect 11756 1584 15200 1612
rect 11756 1572 11762 1584
rect 15194 1572 15200 1584
rect 15252 1572 15258 1624
rect 16546 1612 16574 1652
rect 18782 1640 18788 1692
rect 18840 1680 18846 1692
rect 18840 1652 24164 1680
rect 18840 1640 18846 1652
rect 16546 1584 22140 1612
rect 13906 1544 13912 1556
rect 11624 1516 13912 1544
rect 13906 1504 13912 1516
rect 13964 1504 13970 1556
rect 18874 1544 18880 1556
rect 18708 1516 18880 1544
rect 18708 1476 18736 1516
rect 18874 1504 18880 1516
rect 18932 1504 18938 1556
rect 10612 1448 18736 1476
rect 22112 1476 22140 1584
rect 24136 1544 24164 1652
rect 26602 1640 26608 1692
rect 26660 1680 26666 1692
rect 31386 1680 31392 1692
rect 26660 1652 31392 1680
rect 26660 1640 26666 1652
rect 31386 1640 31392 1652
rect 31444 1640 31450 1692
rect 27154 1572 27160 1624
rect 27212 1612 27218 1624
rect 31202 1612 31208 1624
rect 27212 1584 31208 1612
rect 27212 1572 27218 1584
rect 31202 1572 31208 1584
rect 31260 1572 31266 1624
rect 31496 1612 31524 1788
rect 40678 1708 40684 1760
rect 40736 1708 40742 1760
rect 40696 1612 40724 1708
rect 31496 1584 40724 1612
rect 39666 1544 39672 1556
rect 24136 1516 39672 1544
rect 39666 1504 39672 1516
rect 39724 1504 39730 1556
rect 40310 1504 40316 1556
rect 40368 1504 40374 1556
rect 40328 1476 40356 1504
rect 22112 1448 40356 1476
rect 18598 1408 18604 1420
rect 6886 1380 18604 1408
rect 18598 1368 18604 1380
rect 18656 1368 18662 1420
rect 24118 1368 24124 1420
rect 24176 1408 24182 1420
rect 27154 1408 27160 1420
rect 24176 1380 27160 1408
rect 24176 1368 24182 1380
rect 27154 1368 27160 1380
rect 27212 1368 27218 1420
rect 31202 1368 31208 1420
rect 31260 1408 31266 1420
rect 32122 1408 32128 1420
rect 31260 1380 32128 1408
rect 31260 1368 31266 1380
rect 32122 1368 32128 1380
rect 32180 1368 32186 1420
rect 32398 1368 32404 1420
rect 32456 1408 32462 1420
rect 33134 1408 33140 1420
rect 32456 1380 33140 1408
rect 32456 1368 32462 1380
rect 33134 1368 33140 1380
rect 33192 1368 33198 1420
rect 34054 1368 34060 1420
rect 34112 1408 34118 1420
rect 35434 1408 35440 1420
rect 34112 1380 35440 1408
rect 34112 1368 34118 1380
rect 35434 1368 35440 1380
rect 35492 1368 35498 1420
rect 35894 1368 35900 1420
rect 35952 1408 35958 1420
rect 36814 1408 36820 1420
rect 35952 1380 36820 1408
rect 35952 1368 35958 1380
rect 36814 1368 36820 1380
rect 36872 1368 36878 1420
rect 39850 1368 39856 1420
rect 39908 1408 39914 1420
rect 40402 1408 40408 1420
rect 39908 1380 40408 1408
rect 39908 1368 39914 1380
rect 40402 1368 40408 1380
rect 40460 1368 40466 1420
rect 14734 1300 14740 1352
rect 14792 1340 14798 1352
rect 40862 1340 40868 1352
rect 14792 1312 40868 1340
rect 14792 1300 14798 1312
rect 40862 1300 40868 1312
rect 40920 1300 40926 1352
rect 15102 1232 15108 1284
rect 15160 1272 15166 1284
rect 41138 1272 41144 1284
rect 15160 1244 41144 1272
rect 15160 1232 15166 1244
rect 41138 1232 41144 1244
rect 41196 1232 41202 1284
rect 13906 1164 13912 1216
rect 13964 1204 13970 1216
rect 21542 1204 21548 1216
rect 13964 1176 21548 1204
rect 13964 1164 13970 1176
rect 21542 1164 21548 1176
rect 21600 1164 21606 1216
rect 38378 1164 38384 1216
rect 38436 1164 38442 1216
rect 31386 1096 31392 1148
rect 31444 1136 31450 1148
rect 38396 1136 38424 1164
rect 31444 1108 38424 1136
rect 31444 1096 31450 1108
<< via1 >>
rect 20536 8168 20588 8220
rect 30748 8168 30800 8220
rect 18328 8100 18380 8152
rect 10784 8032 10836 8084
rect 20996 8032 21048 8084
rect 23480 7964 23532 8016
rect 19524 7896 19576 7948
rect 17224 7828 17276 7880
rect 25688 7828 25740 7880
rect 31484 7828 31536 7880
rect 42708 7828 42760 7880
rect 19800 7760 19852 7812
rect 36912 7760 36964 7812
rect 9864 7692 9916 7744
rect 18604 7692 18656 7744
rect 29276 7692 29328 7744
rect 11896 7590 11948 7642
rect 11960 7590 12012 7642
rect 12024 7590 12076 7642
rect 12088 7590 12140 7642
rect 12152 7590 12204 7642
rect 22843 7590 22895 7642
rect 22907 7590 22959 7642
rect 22971 7590 23023 7642
rect 23035 7590 23087 7642
rect 23099 7590 23151 7642
rect 33790 7590 33842 7642
rect 33854 7590 33906 7642
rect 33918 7590 33970 7642
rect 33982 7590 34034 7642
rect 34046 7590 34098 7642
rect 44737 7590 44789 7642
rect 44801 7590 44853 7642
rect 44865 7590 44917 7642
rect 44929 7590 44981 7642
rect 44993 7590 45045 7642
rect 1584 7488 1636 7540
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 3056 7488 3108 7540
rect 3976 7488 4028 7540
rect 4528 7488 4580 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 5908 7531 5960 7540
rect 5908 7497 5917 7531
rect 5917 7497 5951 7531
rect 5951 7497 5960 7531
rect 5908 7488 5960 7497
rect 6828 7488 6880 7540
rect 7380 7531 7432 7540
rect 7380 7497 7389 7531
rect 7389 7497 7423 7531
rect 7423 7497 7432 7531
rect 7380 7488 7432 7497
rect 8944 7488 8996 7540
rect 9680 7488 9732 7540
rect 10508 7531 10560 7540
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 11888 7488 11940 7540
rect 12624 7488 12676 7540
rect 13820 7531 13872 7540
rect 13820 7497 13829 7531
rect 13829 7497 13863 7531
rect 13863 7497 13872 7531
rect 13820 7488 13872 7497
rect 14096 7488 14148 7540
rect 15016 7488 15068 7540
rect 15568 7488 15620 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 3148 7352 3200 7404
rect 4620 7352 4672 7404
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 8300 7463 8352 7472
rect 8300 7429 8309 7463
rect 8309 7429 8343 7463
rect 8343 7429 8352 7463
rect 8300 7420 8352 7429
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 11704 7420 11756 7472
rect 19156 7488 19208 7540
rect 19248 7488 19300 7540
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 19340 7488 19392 7497
rect 19800 7531 19852 7540
rect 19800 7497 19809 7531
rect 19809 7497 19843 7531
rect 19843 7497 19852 7531
rect 19800 7488 19852 7497
rect 19892 7488 19944 7540
rect 23480 7531 23532 7540
rect 23480 7497 23489 7531
rect 23489 7497 23523 7531
rect 23523 7497 23532 7531
rect 23480 7488 23532 7497
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 25688 7531 25740 7540
rect 25688 7497 25697 7531
rect 25697 7497 25731 7531
rect 25731 7497 25740 7531
rect 25688 7488 25740 7497
rect 27896 7488 27948 7540
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 10784 7352 10836 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 10876 7284 10928 7336
rect 8300 7216 8352 7268
rect 13268 7352 13320 7404
rect 13176 7284 13228 7336
rect 14280 7395 14332 7404
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 14648 7352 14700 7404
rect 15108 7352 15160 7404
rect 16488 7395 16540 7404
rect 16488 7361 16497 7395
rect 16497 7361 16531 7395
rect 16531 7361 16540 7395
rect 16488 7352 16540 7361
rect 17040 7352 17092 7404
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18512 7352 18564 7404
rect 19064 7284 19116 7336
rect 19984 7352 20036 7404
rect 19800 7284 19852 7336
rect 8392 7148 8444 7200
rect 8668 7148 8720 7200
rect 14464 7148 14516 7200
rect 17132 7191 17184 7200
rect 17132 7157 17141 7191
rect 17141 7157 17175 7191
rect 17175 7157 17184 7191
rect 17132 7148 17184 7157
rect 18052 7191 18104 7200
rect 18052 7157 18061 7191
rect 18061 7157 18095 7191
rect 18095 7157 18104 7191
rect 18052 7148 18104 7157
rect 20536 7352 20588 7404
rect 20720 7352 20772 7404
rect 21456 7352 21508 7404
rect 22192 7352 22244 7404
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 23204 7395 23256 7404
rect 23204 7361 23213 7395
rect 23213 7361 23247 7395
rect 23247 7361 23256 7395
rect 23204 7352 23256 7361
rect 23296 7395 23348 7404
rect 23296 7361 23305 7395
rect 23305 7361 23339 7395
rect 23339 7361 23348 7395
rect 23296 7352 23348 7361
rect 23664 7352 23716 7404
rect 24400 7352 24452 7404
rect 25044 7352 25096 7404
rect 25136 7352 25188 7404
rect 25596 7395 25648 7404
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 25872 7352 25924 7404
rect 27804 7420 27856 7472
rect 26608 7352 26660 7404
rect 27344 7352 27396 7404
rect 28080 7352 28132 7404
rect 29000 7420 29052 7472
rect 29092 7395 29144 7404
rect 29092 7361 29101 7395
rect 29101 7361 29135 7395
rect 29135 7361 29144 7395
rect 29092 7352 29144 7361
rect 29552 7352 29604 7404
rect 30380 7352 30432 7404
rect 31024 7488 31076 7540
rect 31760 7488 31812 7540
rect 32496 7488 32548 7540
rect 33232 7488 33284 7540
rect 34244 7531 34296 7540
rect 34244 7497 34253 7531
rect 34253 7497 34287 7531
rect 34287 7497 34296 7531
rect 34244 7488 34296 7497
rect 34704 7488 34756 7540
rect 35900 7531 35952 7540
rect 35900 7497 35909 7531
rect 35909 7497 35943 7531
rect 35943 7497 35952 7531
rect 35900 7488 35952 7497
rect 36176 7488 36228 7540
rect 30748 7420 30800 7472
rect 36912 7488 36964 7540
rect 37188 7488 37240 7540
rect 37648 7488 37700 7540
rect 38660 7531 38712 7540
rect 38660 7497 38669 7531
rect 38669 7497 38703 7531
rect 38703 7497 38712 7531
rect 38660 7488 38712 7497
rect 39120 7488 39172 7540
rect 39856 7488 39908 7540
rect 40592 7488 40644 7540
rect 41328 7488 41380 7540
rect 42616 7531 42668 7540
rect 42616 7497 42625 7531
rect 42625 7497 42659 7531
rect 42659 7497 42668 7531
rect 42616 7488 42668 7497
rect 42708 7488 42760 7540
rect 42800 7488 42852 7540
rect 43536 7488 43588 7540
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 33416 7395 33468 7404
rect 33416 7361 33425 7395
rect 33425 7361 33459 7395
rect 33459 7361 33468 7395
rect 33416 7352 33468 7361
rect 34152 7395 34204 7404
rect 34152 7361 34161 7395
rect 34161 7361 34195 7395
rect 34195 7361 34204 7395
rect 34152 7352 34204 7361
rect 34888 7395 34940 7404
rect 34888 7361 34897 7395
rect 34897 7361 34931 7395
rect 34931 7361 34940 7395
rect 34888 7352 34940 7361
rect 35624 7395 35676 7404
rect 35624 7361 35633 7395
rect 35633 7361 35667 7395
rect 35667 7361 35676 7395
rect 35624 7352 35676 7361
rect 35900 7352 35952 7404
rect 37004 7395 37056 7404
rect 37004 7361 37013 7395
rect 37013 7361 37047 7395
rect 37047 7361 37056 7395
rect 37004 7352 37056 7361
rect 37372 7395 37424 7404
rect 37372 7361 37381 7395
rect 37381 7361 37415 7395
rect 37415 7361 37424 7395
rect 37372 7352 37424 7361
rect 37464 7352 37516 7404
rect 38200 7352 38252 7404
rect 38936 7352 38988 7404
rect 39396 7352 39448 7404
rect 23572 7216 23624 7268
rect 25136 7216 25188 7268
rect 29184 7284 29236 7336
rect 29276 7284 29328 7336
rect 29000 7216 29052 7268
rect 19892 7148 19944 7200
rect 20352 7148 20404 7200
rect 21088 7148 21140 7200
rect 22284 7191 22336 7200
rect 22284 7157 22293 7191
rect 22293 7157 22327 7191
rect 22327 7157 22336 7191
rect 22284 7148 22336 7157
rect 23756 7191 23808 7200
rect 23756 7157 23765 7191
rect 23765 7157 23799 7191
rect 23799 7157 23808 7191
rect 23756 7148 23808 7157
rect 24860 7148 24912 7200
rect 27344 7148 27396 7200
rect 28172 7148 28224 7200
rect 28724 7148 28776 7200
rect 29644 7191 29696 7200
rect 29644 7157 29653 7191
rect 29653 7157 29687 7191
rect 29687 7157 29696 7191
rect 29644 7148 29696 7157
rect 31484 7216 31536 7268
rect 31944 7148 31996 7200
rect 33048 7148 33100 7200
rect 39212 7148 39264 7200
rect 42616 7352 42668 7404
rect 6423 7046 6475 7098
rect 6487 7046 6539 7098
rect 6551 7046 6603 7098
rect 6615 7046 6667 7098
rect 6679 7046 6731 7098
rect 17370 7046 17422 7098
rect 17434 7046 17486 7098
rect 17498 7046 17550 7098
rect 17562 7046 17614 7098
rect 17626 7046 17678 7098
rect 28317 7046 28369 7098
rect 28381 7046 28433 7098
rect 28445 7046 28497 7098
rect 28509 7046 28561 7098
rect 28573 7046 28625 7098
rect 39264 7046 39316 7098
rect 39328 7046 39380 7098
rect 39392 7046 39444 7098
rect 39456 7046 39508 7098
rect 39520 7046 39572 7098
rect 9128 6944 9180 6996
rect 23664 6944 23716 6996
rect 25596 6944 25648 6996
rect 22560 6876 22612 6928
rect 27160 6876 27212 6928
rect 34152 6944 34204 6996
rect 34428 6944 34480 6996
rect 34888 6944 34940 6996
rect 35624 6944 35676 6996
rect 37464 6944 37516 6996
rect 38200 6944 38252 6996
rect 38936 6944 38988 6996
rect 44272 6987 44324 6996
rect 44272 6953 44281 6987
rect 44281 6953 44315 6987
rect 44315 6953 44324 6987
rect 44272 6944 44324 6953
rect 848 6808 900 6860
rect 15936 6808 15988 6860
rect 17040 6740 17092 6792
rect 17224 6672 17276 6724
rect 8300 6604 8352 6656
rect 26608 6604 26660 6656
rect 33140 6672 33192 6724
rect 34612 6740 34664 6792
rect 35348 6808 35400 6860
rect 37004 6876 37056 6928
rect 35256 6672 35308 6724
rect 37372 6740 37424 6792
rect 45100 6808 45152 6860
rect 38844 6740 38896 6792
rect 36728 6672 36780 6724
rect 36268 6604 36320 6656
rect 43628 6715 43680 6724
rect 43628 6681 43637 6715
rect 43637 6681 43671 6715
rect 43671 6681 43680 6715
rect 43628 6672 43680 6681
rect 11896 6502 11948 6554
rect 11960 6502 12012 6554
rect 12024 6502 12076 6554
rect 12088 6502 12140 6554
rect 12152 6502 12204 6554
rect 22843 6502 22895 6554
rect 22907 6502 22959 6554
rect 22971 6502 23023 6554
rect 23035 6502 23087 6554
rect 23099 6502 23151 6554
rect 33790 6502 33842 6554
rect 33854 6502 33906 6554
rect 33918 6502 33970 6554
rect 33982 6502 34034 6554
rect 34046 6502 34098 6554
rect 44737 6502 44789 6554
rect 44801 6502 44853 6554
rect 44865 6502 44917 6554
rect 44929 6502 44981 6554
rect 44993 6502 45045 6554
rect 16672 6400 16724 6452
rect 34612 6400 34664 6452
rect 36268 6400 36320 6452
rect 38844 6400 38896 6452
rect 18880 6332 18932 6384
rect 33140 6332 33192 6384
rect 36728 6332 36780 6384
rect 6828 6264 6880 6316
rect 25872 6264 25924 6316
rect 16856 6196 16908 6248
rect 35900 6196 35952 6248
rect 3148 6128 3200 6180
rect 27988 6128 28040 6180
rect 19708 6060 19760 6112
rect 33048 6060 33100 6112
rect 6423 5958 6475 6010
rect 6487 5958 6539 6010
rect 6551 5958 6603 6010
rect 6615 5958 6667 6010
rect 6679 5958 6731 6010
rect 17370 5958 17422 6010
rect 17434 5958 17486 6010
rect 17498 5958 17550 6010
rect 17562 5958 17614 6010
rect 17626 5958 17678 6010
rect 28317 5958 28369 6010
rect 28381 5958 28433 6010
rect 28445 5958 28497 6010
rect 28509 5958 28561 6010
rect 28573 5958 28625 6010
rect 39264 5958 39316 6010
rect 39328 5958 39380 6010
rect 39392 5958 39444 6010
rect 39456 5958 39508 6010
rect 39520 5958 39572 6010
rect 19340 5856 19392 5908
rect 30380 5856 30432 5908
rect 25044 5788 25096 5840
rect 37464 5788 37516 5840
rect 18052 5720 18104 5772
rect 43628 5856 43680 5908
rect 14464 5652 14516 5704
rect 19248 5652 19300 5704
rect 11896 5414 11948 5466
rect 11960 5414 12012 5466
rect 12024 5414 12076 5466
rect 12088 5414 12140 5466
rect 12152 5414 12204 5466
rect 22843 5414 22895 5466
rect 22907 5414 22959 5466
rect 22971 5414 23023 5466
rect 23035 5414 23087 5466
rect 23099 5414 23151 5466
rect 33790 5414 33842 5466
rect 33854 5414 33906 5466
rect 33918 5414 33970 5466
rect 33982 5414 34034 5466
rect 34046 5414 34098 5466
rect 44737 5414 44789 5466
rect 44801 5414 44853 5466
rect 44865 5414 44917 5466
rect 44929 5414 44981 5466
rect 44993 5414 45045 5466
rect 23296 5176 23348 5228
rect 39028 5176 39080 5228
rect 17868 5108 17920 5160
rect 33416 5108 33468 5160
rect 10876 5040 10928 5092
rect 26976 5040 27028 5092
rect 8392 4972 8444 5024
rect 27068 4972 27120 5024
rect 6423 4870 6475 4922
rect 6487 4870 6539 4922
rect 6551 4870 6603 4922
rect 6615 4870 6667 4922
rect 6679 4870 6731 4922
rect 17370 4870 17422 4922
rect 17434 4870 17486 4922
rect 17498 4870 17550 4922
rect 17562 4870 17614 4922
rect 17626 4870 17678 4922
rect 28317 4870 28369 4922
rect 28381 4870 28433 4922
rect 28445 4870 28497 4922
rect 28509 4870 28561 4922
rect 28573 4870 28625 4922
rect 39264 4870 39316 4922
rect 39328 4870 39380 4922
rect 39392 4870 39444 4922
rect 39456 4870 39508 4922
rect 39520 4870 39572 4922
rect 7288 4768 7340 4820
rect 26516 4768 26568 4820
rect 27160 4768 27212 4820
rect 39120 4768 39172 4820
rect 13728 4564 13780 4616
rect 21824 4564 21876 4616
rect 10324 4496 10376 4548
rect 23296 4496 23348 4548
rect 10876 4428 10928 4480
rect 22652 4428 22704 4480
rect 11896 4326 11948 4378
rect 11960 4326 12012 4378
rect 12024 4326 12076 4378
rect 12088 4326 12140 4378
rect 12152 4326 12204 4378
rect 22843 4326 22895 4378
rect 22907 4326 22959 4378
rect 22971 4326 23023 4378
rect 23035 4326 23087 4378
rect 23099 4326 23151 4378
rect 33790 4326 33842 4378
rect 33854 4326 33906 4378
rect 33918 4326 33970 4378
rect 33982 4326 34034 4378
rect 34046 4326 34098 4378
rect 44737 4326 44789 4378
rect 44801 4326 44853 4378
rect 44865 4326 44917 4378
rect 44929 4326 44981 4378
rect 44993 4326 45045 4378
rect 17224 4224 17276 4276
rect 30748 4224 30800 4276
rect 11060 4156 11112 4208
rect 18788 4156 18840 4208
rect 9680 4088 9732 4140
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 10692 4020 10744 4072
rect 21640 4131 21692 4140
rect 21640 4097 21649 4131
rect 21649 4097 21683 4131
rect 21683 4097 21692 4131
rect 21640 4088 21692 4097
rect 21824 4156 21876 4208
rect 32036 4156 32088 4208
rect 26700 4088 26752 4140
rect 26792 4131 26844 4140
rect 26792 4097 26801 4131
rect 26801 4097 26835 4131
rect 26835 4097 26844 4131
rect 26792 4088 26844 4097
rect 32680 4131 32732 4140
rect 32680 4097 32689 4131
rect 32689 4097 32723 4131
rect 32723 4097 32732 4131
rect 32680 4088 32732 4097
rect 31024 4020 31076 4072
rect 16764 3952 16816 4004
rect 18880 3952 18932 4004
rect 19064 3995 19116 4004
rect 19064 3961 19073 3995
rect 19073 3961 19107 3995
rect 19107 3961 19116 3995
rect 19064 3952 19116 3961
rect 19432 3952 19484 4004
rect 21548 3952 21600 4004
rect 23112 3952 23164 4004
rect 23296 3952 23348 4004
rect 24400 3952 24452 4004
rect 26516 3995 26568 4004
rect 26516 3961 26525 3995
rect 26525 3961 26559 3995
rect 26559 3961 26568 3995
rect 26516 3952 26568 3961
rect 18512 3884 18564 3936
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 21180 3884 21232 3893
rect 21456 3927 21508 3936
rect 21456 3893 21465 3927
rect 21465 3893 21499 3927
rect 21499 3893 21508 3927
rect 21456 3884 21508 3893
rect 22100 3884 22152 3936
rect 22376 3884 22428 3936
rect 25412 3884 25464 3936
rect 27160 3884 27212 3936
rect 33416 3884 33468 3936
rect 6423 3782 6475 3834
rect 6487 3782 6539 3834
rect 6551 3782 6603 3834
rect 6615 3782 6667 3834
rect 6679 3782 6731 3834
rect 17370 3782 17422 3834
rect 17434 3782 17486 3834
rect 17498 3782 17550 3834
rect 17562 3782 17614 3834
rect 17626 3782 17678 3834
rect 28317 3782 28369 3834
rect 28381 3782 28433 3834
rect 28445 3782 28497 3834
rect 28509 3782 28561 3834
rect 28573 3782 28625 3834
rect 39264 3782 39316 3834
rect 39328 3782 39380 3834
rect 39392 3782 39444 3834
rect 39456 3782 39508 3834
rect 39520 3782 39572 3834
rect 10968 3680 11020 3732
rect 18788 3680 18840 3732
rect 16580 3612 16632 3664
rect 16488 3476 16540 3528
rect 16764 3655 16816 3664
rect 16764 3621 16773 3655
rect 16773 3621 16807 3655
rect 16807 3621 16816 3655
rect 16764 3612 16816 3621
rect 17868 3612 17920 3664
rect 19800 3680 19852 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 20996 3723 21048 3732
rect 20996 3689 21005 3723
rect 21005 3689 21039 3723
rect 21039 3689 21048 3723
rect 20996 3680 21048 3689
rect 21548 3680 21600 3732
rect 28724 3680 28776 3732
rect 29828 3723 29880 3732
rect 29828 3689 29837 3723
rect 29837 3689 29871 3723
rect 29871 3689 29880 3723
rect 29828 3680 29880 3689
rect 30840 3723 30892 3732
rect 30840 3689 30849 3723
rect 30849 3689 30883 3723
rect 30883 3689 30892 3723
rect 30840 3680 30892 3689
rect 32772 3680 32824 3732
rect 33140 3680 33192 3732
rect 16948 3408 17000 3460
rect 11244 3340 11296 3392
rect 17684 3476 17736 3528
rect 17868 3519 17920 3528
rect 17868 3485 17877 3519
rect 17877 3485 17911 3519
rect 17911 3485 17920 3519
rect 17868 3476 17920 3485
rect 18420 3519 18472 3528
rect 18420 3485 18429 3519
rect 18429 3485 18463 3519
rect 18463 3485 18472 3519
rect 18420 3476 18472 3485
rect 18788 3408 18840 3460
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 20352 3476 20404 3528
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 21088 3476 21140 3528
rect 22284 3612 22336 3664
rect 21548 3476 21600 3528
rect 22192 3519 22244 3528
rect 22192 3485 22201 3519
rect 22201 3485 22235 3519
rect 22235 3485 22244 3519
rect 22192 3476 22244 3485
rect 22284 3476 22336 3528
rect 22468 3519 22520 3528
rect 22468 3485 22477 3519
rect 22477 3485 22511 3519
rect 22511 3485 22520 3519
rect 22468 3476 22520 3485
rect 23480 3612 23532 3664
rect 23572 3612 23624 3664
rect 23664 3612 23716 3664
rect 24768 3612 24820 3664
rect 24860 3612 24912 3664
rect 25872 3655 25924 3664
rect 25872 3621 25881 3655
rect 25881 3621 25915 3655
rect 25915 3621 25924 3655
rect 25872 3612 25924 3621
rect 26608 3655 26660 3664
rect 26608 3621 26617 3655
rect 26617 3621 26651 3655
rect 26651 3621 26660 3655
rect 26608 3612 26660 3621
rect 26976 3655 27028 3664
rect 26976 3621 26985 3655
rect 26985 3621 27019 3655
rect 27019 3621 27028 3655
rect 26976 3612 27028 3621
rect 27068 3612 27120 3664
rect 23204 3519 23256 3528
rect 23204 3485 23213 3519
rect 23213 3485 23247 3519
rect 23247 3485 23256 3519
rect 23204 3476 23256 3485
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 24308 3476 24360 3528
rect 25136 3544 25188 3596
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 25688 3519 25740 3528
rect 25688 3485 25697 3519
rect 25697 3485 25731 3519
rect 25731 3485 25740 3519
rect 25688 3476 25740 3485
rect 17684 3383 17736 3392
rect 17684 3349 17693 3383
rect 17693 3349 17727 3383
rect 17727 3349 17736 3383
rect 17684 3340 17736 3349
rect 17868 3340 17920 3392
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 18236 3383 18288 3392
rect 18236 3349 18245 3383
rect 18245 3349 18279 3383
rect 18279 3349 18288 3383
rect 18236 3340 18288 3349
rect 18880 3383 18932 3392
rect 18880 3349 18889 3383
rect 18889 3349 18923 3383
rect 18923 3349 18932 3383
rect 18880 3340 18932 3349
rect 19064 3340 19116 3392
rect 19524 3383 19576 3392
rect 19524 3349 19533 3383
rect 19533 3349 19567 3383
rect 19567 3349 19576 3383
rect 19524 3340 19576 3349
rect 19800 3383 19852 3392
rect 19800 3349 19809 3383
rect 19809 3349 19843 3383
rect 19843 3349 19852 3383
rect 19800 3340 19852 3349
rect 19984 3340 20036 3392
rect 20904 3340 20956 3392
rect 21732 3383 21784 3392
rect 21732 3349 21741 3383
rect 21741 3349 21775 3383
rect 21775 3349 21784 3383
rect 21732 3340 21784 3349
rect 22008 3383 22060 3392
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 22284 3383 22336 3392
rect 22284 3349 22293 3383
rect 22293 3349 22327 3383
rect 22327 3349 22336 3383
rect 22284 3340 22336 3349
rect 22744 3383 22796 3392
rect 22744 3349 22753 3383
rect 22753 3349 22787 3383
rect 22787 3349 22796 3383
rect 22744 3340 22796 3349
rect 23112 3340 23164 3392
rect 24124 3408 24176 3460
rect 27712 3544 27764 3596
rect 27804 3544 27856 3596
rect 29460 3612 29512 3664
rect 27528 3476 27580 3528
rect 27620 3519 27672 3528
rect 27620 3485 27629 3519
rect 27629 3485 27663 3519
rect 27663 3485 27672 3519
rect 27620 3476 27672 3485
rect 26792 3451 26844 3460
rect 26792 3417 26801 3451
rect 26801 3417 26835 3451
rect 26835 3417 26844 3451
rect 26792 3408 26844 3417
rect 27344 3408 27396 3460
rect 28264 3476 28316 3528
rect 29000 3544 29052 3596
rect 29184 3544 29236 3596
rect 30564 3544 30616 3596
rect 29644 3476 29696 3528
rect 30288 3476 30340 3528
rect 35440 3544 35492 3596
rect 31208 3519 31260 3528
rect 31208 3485 31217 3519
rect 31217 3485 31251 3519
rect 31251 3485 31260 3519
rect 31208 3476 31260 3485
rect 31484 3519 31536 3528
rect 31484 3485 31493 3519
rect 31493 3485 31527 3519
rect 31527 3485 31536 3519
rect 31484 3476 31536 3485
rect 31760 3519 31812 3528
rect 31760 3485 31769 3519
rect 31769 3485 31803 3519
rect 31803 3485 31812 3519
rect 31760 3476 31812 3485
rect 32036 3519 32088 3528
rect 32036 3485 32045 3519
rect 32045 3485 32079 3519
rect 32079 3485 32088 3519
rect 32036 3476 32088 3485
rect 32312 3519 32364 3528
rect 32312 3485 32321 3519
rect 32321 3485 32355 3519
rect 32355 3485 32364 3519
rect 32312 3476 32364 3485
rect 32588 3519 32640 3528
rect 32588 3485 32597 3519
rect 32597 3485 32631 3519
rect 32631 3485 32640 3519
rect 32588 3476 32640 3485
rect 24492 3383 24544 3392
rect 24492 3349 24501 3383
rect 24501 3349 24535 3383
rect 24535 3349 24544 3383
rect 24492 3340 24544 3349
rect 24768 3383 24820 3392
rect 24768 3349 24777 3383
rect 24777 3349 24811 3383
rect 24811 3349 24820 3383
rect 24768 3340 24820 3349
rect 25044 3383 25096 3392
rect 25044 3349 25053 3383
rect 25053 3349 25087 3383
rect 25087 3349 25096 3383
rect 25044 3340 25096 3349
rect 25320 3383 25372 3392
rect 25320 3349 25329 3383
rect 25329 3349 25363 3383
rect 25363 3349 25372 3383
rect 25320 3340 25372 3349
rect 25964 3383 26016 3392
rect 25964 3349 25973 3383
rect 25973 3349 26007 3383
rect 26007 3349 26016 3383
rect 25964 3340 26016 3349
rect 27712 3383 27764 3392
rect 27712 3349 27721 3383
rect 27721 3349 27755 3383
rect 27755 3349 27764 3383
rect 27712 3340 27764 3349
rect 27988 3340 28040 3392
rect 30656 3408 30708 3460
rect 28172 3383 28224 3392
rect 28172 3349 28181 3383
rect 28181 3349 28215 3383
rect 28215 3349 28224 3383
rect 28172 3340 28224 3349
rect 28632 3383 28684 3392
rect 28632 3349 28641 3383
rect 28641 3349 28675 3383
rect 28675 3349 28684 3383
rect 28632 3340 28684 3349
rect 28908 3383 28960 3392
rect 28908 3349 28917 3383
rect 28917 3349 28951 3383
rect 28951 3349 28960 3383
rect 28908 3340 28960 3349
rect 29184 3383 29236 3392
rect 29184 3349 29193 3383
rect 29193 3349 29227 3383
rect 29227 3349 29236 3383
rect 29184 3340 29236 3349
rect 30012 3383 30064 3392
rect 30012 3349 30021 3383
rect 30021 3349 30055 3383
rect 30055 3349 30064 3383
rect 30012 3340 30064 3349
rect 30288 3383 30340 3392
rect 30288 3349 30297 3383
rect 30297 3349 30331 3383
rect 30331 3349 30340 3383
rect 30288 3340 30340 3349
rect 32496 3408 32548 3460
rect 32956 3451 33008 3460
rect 32956 3417 32965 3451
rect 32965 3417 32999 3451
rect 32999 3417 33008 3451
rect 32956 3408 33008 3417
rect 31300 3383 31352 3392
rect 31300 3349 31309 3383
rect 31309 3349 31343 3383
rect 31343 3349 31352 3383
rect 31300 3340 31352 3349
rect 31852 3383 31904 3392
rect 31852 3349 31861 3383
rect 31861 3349 31895 3383
rect 31895 3349 31904 3383
rect 31852 3340 31904 3349
rect 32128 3383 32180 3392
rect 32128 3349 32137 3383
rect 32137 3349 32171 3383
rect 32171 3349 32180 3383
rect 32128 3340 32180 3349
rect 32864 3340 32916 3392
rect 11896 3238 11948 3290
rect 11960 3238 12012 3290
rect 12024 3238 12076 3290
rect 12088 3238 12140 3290
rect 12152 3238 12204 3290
rect 22843 3238 22895 3290
rect 22907 3238 22959 3290
rect 22971 3238 23023 3290
rect 23035 3238 23087 3290
rect 23099 3238 23151 3290
rect 33790 3238 33842 3290
rect 33854 3238 33906 3290
rect 33918 3238 33970 3290
rect 33982 3238 34034 3290
rect 34046 3238 34098 3290
rect 44737 3238 44789 3290
rect 44801 3238 44853 3290
rect 44865 3238 44917 3290
rect 44929 3238 44981 3290
rect 44993 3238 45045 3290
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 17132 3136 17184 3188
rect 17224 3179 17276 3188
rect 17224 3145 17233 3179
rect 17233 3145 17267 3179
rect 17267 3145 17276 3179
rect 17224 3136 17276 3145
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 14372 3000 14424 3009
rect 16856 3000 16908 3052
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 17224 2932 17276 2984
rect 17960 3136 18012 3188
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 17684 3111 17736 3120
rect 17684 3077 17695 3111
rect 17695 3077 17729 3111
rect 17729 3077 17736 3111
rect 17684 3068 17736 3077
rect 18236 3068 18288 3120
rect 19524 3136 19576 3188
rect 18880 3068 18932 3120
rect 21456 3136 21508 3188
rect 21732 3136 21784 3188
rect 18144 3000 18196 3052
rect 18512 2932 18564 2984
rect 17960 2864 18012 2916
rect 18328 2864 18380 2916
rect 19064 2932 19116 2984
rect 19616 2932 19668 2984
rect 19708 2932 19760 2984
rect 19984 2932 20036 2984
rect 22284 3136 22336 3188
rect 23756 3136 23808 3188
rect 24032 3179 24084 3188
rect 24032 3145 24041 3179
rect 24041 3145 24075 3179
rect 24075 3145 24084 3179
rect 24032 3136 24084 3145
rect 24492 3136 24544 3188
rect 25320 3136 25372 3188
rect 25412 3136 25464 3188
rect 22008 3043 22060 3052
rect 22008 3009 22017 3043
rect 22017 3009 22051 3043
rect 22051 3009 22060 3043
rect 22008 3000 22060 3009
rect 22468 3000 22520 3052
rect 22652 3000 22704 3052
rect 25964 3136 26016 3188
rect 27160 3136 27212 3188
rect 27528 3136 27580 3188
rect 28632 3136 28684 3188
rect 29184 3136 29236 3188
rect 29736 3136 29788 3188
rect 30564 3136 30616 3188
rect 31300 3136 31352 3188
rect 27712 3068 27764 3120
rect 24400 3000 24452 3052
rect 30012 3068 30064 3120
rect 30380 3111 30432 3120
rect 30380 3077 30389 3111
rect 30389 3077 30423 3111
rect 30423 3077 30432 3111
rect 30380 3068 30432 3077
rect 19156 2864 19208 2916
rect 30656 3068 30708 3120
rect 31392 3068 31444 3120
rect 31852 3136 31904 3188
rect 32496 3068 32548 3120
rect 32680 3068 32732 3120
rect 32864 3136 32916 3188
rect 33600 3136 33652 3188
rect 35440 3179 35492 3188
rect 35440 3145 35449 3179
rect 35449 3145 35483 3179
rect 35483 3145 35492 3179
rect 35440 3136 35492 3145
rect 39120 3179 39172 3188
rect 39120 3145 39129 3179
rect 39129 3145 39163 3179
rect 39163 3145 39172 3179
rect 39120 3136 39172 3145
rect 30748 3000 30800 3052
rect 31024 3000 31076 3052
rect 32128 3000 32180 3052
rect 32864 3000 32916 3052
rect 33416 3000 33468 3052
rect 34336 3000 34388 3052
rect 35072 3000 35124 3052
rect 38936 3043 38988 3052
rect 38936 3009 38945 3043
rect 38945 3009 38979 3043
rect 38979 3009 38988 3043
rect 38936 3000 38988 3009
rect 22652 2864 22704 2916
rect 14556 2796 14608 2848
rect 16396 2796 16448 2848
rect 17132 2796 17184 2848
rect 17316 2796 17368 2848
rect 18696 2796 18748 2848
rect 20260 2839 20312 2848
rect 20260 2805 20269 2839
rect 20269 2805 20303 2839
rect 20303 2805 20312 2839
rect 20260 2796 20312 2805
rect 20628 2796 20680 2848
rect 21364 2839 21416 2848
rect 21364 2805 21373 2839
rect 21373 2805 21407 2839
rect 21407 2805 21416 2839
rect 21364 2796 21416 2805
rect 21824 2839 21876 2848
rect 21824 2805 21833 2839
rect 21833 2805 21867 2839
rect 21867 2805 21876 2839
rect 21824 2796 21876 2805
rect 22008 2796 22060 2848
rect 22560 2796 22612 2848
rect 23388 2839 23440 2848
rect 23388 2805 23397 2839
rect 23397 2805 23431 2839
rect 23431 2805 23440 2839
rect 23388 2796 23440 2805
rect 24216 2796 24268 2848
rect 25412 2864 25464 2916
rect 26976 2864 27028 2916
rect 24492 2796 24544 2848
rect 25044 2796 25096 2848
rect 25596 2796 25648 2848
rect 26056 2796 26108 2848
rect 26608 2796 26660 2848
rect 29184 2864 29236 2916
rect 28448 2796 28500 2848
rect 28908 2796 28960 2848
rect 30564 2864 30616 2916
rect 30196 2796 30248 2848
rect 32036 2864 32088 2916
rect 33048 2864 33100 2916
rect 31668 2796 31720 2848
rect 32496 2796 32548 2848
rect 34152 2796 34204 2848
rect 6423 2694 6475 2746
rect 6487 2694 6539 2746
rect 6551 2694 6603 2746
rect 6615 2694 6667 2746
rect 6679 2694 6731 2746
rect 17370 2694 17422 2746
rect 17434 2694 17486 2746
rect 17498 2694 17550 2746
rect 17562 2694 17614 2746
rect 17626 2694 17678 2746
rect 28317 2694 28369 2746
rect 28381 2694 28433 2746
rect 28445 2694 28497 2746
rect 28509 2694 28561 2746
rect 28573 2694 28625 2746
rect 39264 2694 39316 2746
rect 39328 2694 39380 2746
rect 39392 2694 39444 2746
rect 39456 2694 39508 2746
rect 39520 2694 39572 2746
rect 6736 2592 6788 2644
rect 9588 2592 9640 2644
rect 9680 2635 9732 2644
rect 9680 2601 9689 2635
rect 9689 2601 9723 2635
rect 9723 2601 9732 2635
rect 9680 2592 9732 2601
rect 9956 2635 10008 2644
rect 9956 2601 9965 2635
rect 9965 2601 9999 2635
rect 9999 2601 10008 2635
rect 9956 2592 10008 2601
rect 10232 2524 10284 2576
rect 12992 2592 13044 2644
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 13268 2592 13320 2644
rect 16948 2592 17000 2644
rect 18328 2635 18380 2644
rect 18328 2601 18337 2635
rect 18337 2601 18371 2635
rect 18371 2601 18380 2635
rect 18328 2592 18380 2601
rect 19984 2592 20036 2644
rect 20812 2592 20864 2644
rect 23204 2592 23256 2644
rect 24400 2592 24452 2644
rect 25504 2592 25556 2644
rect 26516 2592 26568 2644
rect 26884 2592 26936 2644
rect 28632 2592 28684 2644
rect 11060 2567 11112 2576
rect 11060 2533 11069 2567
rect 11069 2533 11103 2567
rect 11103 2533 11112 2567
rect 11060 2524 11112 2533
rect 11336 2567 11388 2576
rect 11336 2533 11345 2567
rect 11345 2533 11379 2567
rect 11379 2533 11388 2567
rect 11336 2524 11388 2533
rect 5632 2388 5684 2440
rect 5908 2388 5960 2440
rect 6276 2388 6328 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 11244 2456 11296 2508
rect 14464 2524 14516 2576
rect 14648 2524 14700 2576
rect 16396 2524 16448 2576
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7472 2431 7524 2440
rect 7472 2397 7481 2431
rect 7481 2397 7515 2431
rect 7515 2397 7524 2431
rect 7472 2388 7524 2397
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 8484 2388 8536 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 8760 2388 8812 2440
rect 5632 2295 5684 2304
rect 5632 2261 5641 2295
rect 5641 2261 5675 2295
rect 5675 2261 5684 2295
rect 5632 2252 5684 2261
rect 7104 2252 7156 2304
rect 7380 2295 7432 2304
rect 7380 2261 7389 2295
rect 7389 2261 7423 2295
rect 7423 2261 7432 2295
rect 7380 2252 7432 2261
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8208 2295 8260 2304
rect 8208 2261 8217 2295
rect 8217 2261 8251 2295
rect 8251 2261 8260 2295
rect 8208 2252 8260 2261
rect 8392 2252 8444 2304
rect 9404 2388 9456 2440
rect 9680 2388 9732 2440
rect 9312 2320 9364 2372
rect 10416 2388 10468 2440
rect 10508 2431 10560 2440
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 10692 2388 10744 2440
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11060 2388 11112 2440
rect 11428 2388 11480 2440
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 11980 2388 12032 2440
rect 10140 2320 10192 2372
rect 9220 2252 9272 2304
rect 9496 2252 9548 2304
rect 11888 2320 11940 2372
rect 12532 2388 12584 2440
rect 12808 2388 12860 2440
rect 13176 2388 13228 2440
rect 13268 2388 13320 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 13636 2388 13688 2440
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 14648 2388 14700 2440
rect 14740 2431 14792 2440
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10600 2252 10652 2261
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 12532 2295 12584 2304
rect 12532 2261 12541 2295
rect 12541 2261 12575 2295
rect 12575 2261 12584 2295
rect 12532 2252 12584 2261
rect 13084 2295 13136 2304
rect 13084 2261 13093 2295
rect 13093 2261 13127 2295
rect 13127 2261 13136 2295
rect 13084 2252 13136 2261
rect 14556 2320 14608 2372
rect 15108 2456 15160 2508
rect 15384 2456 15436 2508
rect 15936 2499 15988 2508
rect 15936 2465 15945 2499
rect 15945 2465 15979 2499
rect 15979 2465 15988 2499
rect 15936 2456 15988 2465
rect 16856 2456 16908 2508
rect 18052 2456 18104 2508
rect 15200 2388 15252 2440
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 15844 2388 15896 2440
rect 16396 2388 16448 2440
rect 17132 2388 17184 2440
rect 19708 2456 19760 2508
rect 20352 2456 20404 2508
rect 20720 2456 20772 2508
rect 21824 2456 21876 2508
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 18604 2388 18656 2440
rect 18880 2388 18932 2440
rect 19340 2388 19392 2440
rect 19800 2388 19852 2440
rect 21180 2388 21232 2440
rect 21548 2388 21600 2440
rect 22100 2388 22152 2440
rect 14188 2252 14240 2304
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 16856 2320 16908 2372
rect 18052 2295 18104 2304
rect 18052 2261 18061 2295
rect 18061 2261 18095 2295
rect 18095 2261 18104 2295
rect 18052 2252 18104 2261
rect 21456 2320 21508 2372
rect 21640 2363 21692 2372
rect 21640 2329 21649 2363
rect 21649 2329 21683 2363
rect 21683 2329 21692 2363
rect 21640 2320 21692 2329
rect 22376 2320 22428 2372
rect 23572 2388 23624 2440
rect 24860 2388 24912 2440
rect 25228 2388 25280 2440
rect 25412 2388 25464 2440
rect 26608 2431 26660 2440
rect 26608 2397 26617 2431
rect 26617 2397 26651 2431
rect 26651 2397 26660 2431
rect 26608 2388 26660 2397
rect 27896 2388 27948 2440
rect 21916 2252 21968 2304
rect 26332 2320 26384 2372
rect 22836 2295 22888 2304
rect 22836 2261 22845 2295
rect 22845 2261 22879 2295
rect 22879 2261 22888 2295
rect 22836 2252 22888 2261
rect 23572 2295 23624 2304
rect 23572 2261 23581 2295
rect 23581 2261 23615 2295
rect 23615 2261 23624 2295
rect 23572 2252 23624 2261
rect 23664 2252 23716 2304
rect 24032 2252 24084 2304
rect 24952 2252 25004 2304
rect 27068 2363 27120 2372
rect 27068 2329 27077 2363
rect 27077 2329 27111 2363
rect 27111 2329 27120 2363
rect 27068 2320 27120 2329
rect 27436 2320 27488 2372
rect 28908 2524 28960 2576
rect 28080 2456 28132 2508
rect 29552 2456 29604 2508
rect 31116 2592 31168 2644
rect 32956 2592 33008 2644
rect 33508 2592 33560 2644
rect 35900 2592 35952 2644
rect 36636 2635 36688 2644
rect 36636 2601 36645 2635
rect 36645 2601 36679 2635
rect 36679 2601 36688 2635
rect 36636 2592 36688 2601
rect 37096 2635 37148 2644
rect 37096 2601 37105 2635
rect 37105 2601 37139 2635
rect 37139 2601 37148 2635
rect 37096 2592 37148 2601
rect 37464 2635 37516 2644
rect 37464 2601 37473 2635
rect 37473 2601 37507 2635
rect 37507 2601 37516 2635
rect 37464 2592 37516 2601
rect 37832 2592 37884 2644
rect 39028 2592 39080 2644
rect 28540 2388 28592 2440
rect 28724 2431 28776 2440
rect 28724 2397 28733 2431
rect 28733 2397 28767 2431
rect 28767 2397 28776 2431
rect 28724 2388 28776 2397
rect 29092 2388 29144 2440
rect 29368 2431 29420 2440
rect 29368 2397 29377 2431
rect 29377 2397 29411 2431
rect 29411 2397 29420 2431
rect 29368 2388 29420 2397
rect 29460 2388 29512 2440
rect 30748 2431 30800 2440
rect 30748 2397 30757 2431
rect 30757 2397 30791 2431
rect 30791 2397 30800 2431
rect 30748 2388 30800 2397
rect 30840 2388 30892 2440
rect 34428 2524 34480 2576
rect 37004 2524 37056 2576
rect 31668 2456 31720 2508
rect 35256 2456 35308 2508
rect 31392 2388 31444 2440
rect 29000 2320 29052 2372
rect 30380 2320 30432 2372
rect 31944 2431 31996 2440
rect 31944 2397 31953 2431
rect 31953 2397 31987 2431
rect 31987 2397 31996 2431
rect 31944 2388 31996 2397
rect 32220 2363 32272 2372
rect 32220 2329 32229 2363
rect 32229 2329 32263 2363
rect 32263 2329 32272 2363
rect 32220 2320 32272 2329
rect 32680 2388 32732 2440
rect 32864 2388 32916 2440
rect 33140 2388 33192 2440
rect 33416 2388 33468 2440
rect 36544 2456 36596 2508
rect 29644 2252 29696 2304
rect 30104 2252 30156 2304
rect 34336 2320 34388 2372
rect 34796 2363 34848 2372
rect 34796 2329 34805 2363
rect 34805 2329 34839 2363
rect 34839 2329 34848 2363
rect 34796 2320 34848 2329
rect 35348 2363 35400 2372
rect 35348 2329 35357 2363
rect 35357 2329 35391 2363
rect 35391 2329 35400 2363
rect 35348 2320 35400 2329
rect 35900 2320 35952 2372
rect 36820 2431 36872 2440
rect 36820 2397 36829 2431
rect 36829 2397 36863 2431
rect 36863 2397 36872 2431
rect 36820 2388 36872 2397
rect 38108 2524 38160 2576
rect 38844 2524 38896 2576
rect 37924 2456 37976 2508
rect 38476 2456 38528 2508
rect 33140 2252 33192 2304
rect 35440 2295 35492 2304
rect 35440 2261 35449 2295
rect 35449 2261 35483 2295
rect 35483 2261 35492 2295
rect 35440 2252 35492 2261
rect 36084 2252 36136 2304
rect 36544 2295 36596 2304
rect 36544 2261 36553 2295
rect 36553 2261 36587 2295
rect 36587 2261 36596 2295
rect 36544 2252 36596 2261
rect 36636 2252 36688 2304
rect 37648 2320 37700 2372
rect 38200 2320 38252 2372
rect 38752 2320 38804 2372
rect 39396 2456 39448 2508
rect 40040 2456 40092 2508
rect 39120 2320 39172 2372
rect 40408 2431 40460 2440
rect 40408 2397 40417 2431
rect 40417 2397 40451 2431
rect 40451 2397 40460 2431
rect 40408 2388 40460 2397
rect 40224 2320 40276 2372
rect 37740 2295 37792 2304
rect 37740 2261 37749 2295
rect 37749 2261 37783 2295
rect 37783 2261 37792 2295
rect 37740 2252 37792 2261
rect 38384 2252 38436 2304
rect 39028 2252 39080 2304
rect 39304 2252 39356 2304
rect 39672 2295 39724 2304
rect 39672 2261 39681 2295
rect 39681 2261 39715 2295
rect 39715 2261 39724 2295
rect 39672 2252 39724 2261
rect 40040 2295 40092 2304
rect 40040 2261 40049 2295
rect 40049 2261 40083 2295
rect 40083 2261 40092 2295
rect 40040 2252 40092 2261
rect 40316 2295 40368 2304
rect 40316 2261 40325 2295
rect 40325 2261 40359 2295
rect 40359 2261 40368 2295
rect 40316 2252 40368 2261
rect 40684 2252 40736 2304
rect 40868 2295 40920 2304
rect 40868 2261 40877 2295
rect 40877 2261 40911 2295
rect 40911 2261 40920 2295
rect 40868 2252 40920 2261
rect 41144 2295 41196 2304
rect 41144 2261 41153 2295
rect 41153 2261 41187 2295
rect 41187 2261 41196 2295
rect 41144 2252 41196 2261
rect 11896 2150 11948 2202
rect 11960 2150 12012 2202
rect 12024 2150 12076 2202
rect 12088 2150 12140 2202
rect 12152 2150 12204 2202
rect 22843 2150 22895 2202
rect 22907 2150 22959 2202
rect 22971 2150 23023 2202
rect 23035 2150 23087 2202
rect 23099 2150 23151 2202
rect 33790 2150 33842 2202
rect 33854 2150 33906 2202
rect 33918 2150 33970 2202
rect 33982 2150 34034 2202
rect 34046 2150 34098 2202
rect 44737 2150 44789 2202
rect 44801 2150 44853 2202
rect 44865 2150 44917 2202
rect 44929 2150 44981 2202
rect 44993 2150 45045 2202
rect 8208 2048 8260 2100
rect 8392 2048 8444 2100
rect 10876 2048 10928 2100
rect 14464 2048 14516 2100
rect 15292 2048 15344 2100
rect 15384 2048 15436 2100
rect 27160 1980 27212 2032
rect 19156 1912 19208 1964
rect 19892 1912 19944 1964
rect 20996 1912 21048 1964
rect 27068 1912 27120 1964
rect 28540 2048 28592 2100
rect 27344 1980 27396 2032
rect 29000 1980 29052 2032
rect 29368 1980 29420 2032
rect 29644 2048 29696 2100
rect 34796 2048 34848 2100
rect 35348 2048 35400 2100
rect 39028 2048 39080 2100
rect 30840 1980 30892 2032
rect 30288 1912 30340 1964
rect 14648 1844 14700 1896
rect 9220 1776 9272 1828
rect 15568 1776 15620 1828
rect 18052 1844 18104 1896
rect 23204 1844 23256 1896
rect 32128 1912 32180 1964
rect 39304 1912 39356 1964
rect 5632 1640 5684 1692
rect 7380 1640 7432 1692
rect 10324 1640 10376 1692
rect 10600 1640 10652 1692
rect 12532 1708 12584 1760
rect 31208 1708 31260 1760
rect 13360 1640 13412 1692
rect 11704 1572 11756 1624
rect 15200 1572 15252 1624
rect 18788 1640 18840 1692
rect 13912 1504 13964 1556
rect 18880 1504 18932 1556
rect 26608 1640 26660 1692
rect 31392 1640 31444 1692
rect 27160 1572 27212 1624
rect 31208 1572 31260 1624
rect 40684 1708 40736 1760
rect 39672 1504 39724 1556
rect 40316 1504 40368 1556
rect 18604 1368 18656 1420
rect 24124 1368 24176 1420
rect 27160 1368 27212 1420
rect 31208 1368 31260 1420
rect 32128 1368 32180 1420
rect 32404 1368 32456 1420
rect 33140 1368 33192 1420
rect 34060 1368 34112 1420
rect 35440 1368 35492 1420
rect 35900 1368 35952 1420
rect 36820 1368 36872 1420
rect 39856 1368 39908 1420
rect 40408 1368 40460 1420
rect 14740 1300 14792 1352
rect 40868 1300 40920 1352
rect 15108 1232 15160 1284
rect 41144 1232 41196 1284
rect 13912 1164 13964 1216
rect 21548 1164 21600 1216
rect 38384 1164 38436 1216
rect 31392 1096 31444 1148
<< metal2 >>
rect 846 9840 902 10000
rect 1582 9840 1638 10000
rect 2318 9840 2374 10000
rect 2424 9846 2728 9874
rect 860 6866 888 9840
rect 1596 7546 1624 9840
rect 2332 9738 2360 9840
rect 2424 9738 2452 9846
rect 2332 9710 2452 9738
rect 2700 8242 2728 9846
rect 3054 9840 3110 10000
rect 3790 9840 3846 10000
rect 4526 9840 4582 10000
rect 5262 9840 5318 10000
rect 5998 9840 6054 10000
rect 6734 9840 6790 10000
rect 7470 9840 7526 10000
rect 8206 9840 8262 10000
rect 8942 9840 8998 10000
rect 9678 9840 9734 10000
rect 10414 9840 10470 10000
rect 11150 9840 11206 10000
rect 11886 9840 11942 10000
rect 12622 9840 12678 10000
rect 13358 9840 13414 10000
rect 13464 9846 13768 9874
rect 2700 8214 2820 8242
rect 2792 7546 2820 8214
rect 3068 7546 3096 9840
rect 3804 8514 3832 9840
rect 3804 8486 4016 8514
rect 3988 7546 4016 8486
rect 4540 7546 4568 9840
rect 5276 8242 5304 9840
rect 6012 8514 6040 9840
rect 6748 8650 6776 9840
rect 6748 8622 6868 8650
rect 5920 8486 6040 8514
rect 5276 8214 5580 8242
rect 5552 7546 5580 8214
rect 5920 7546 5948 8486
rect 6840 7546 6868 8622
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 7380 7540 7432 7546
rect 7484 7528 7512 9840
rect 8220 8242 8248 9840
rect 8220 8214 8340 8242
rect 7432 7500 7512 7528
rect 7380 7482 7432 7488
rect 8312 7478 8340 8214
rect 8956 7546 8984 9840
rect 9692 7546 9720 9840
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 8300 7472 8352 7478
rect 1766 7440 1822 7449
rect 8300 7414 8352 7420
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 1766 7375 1768 7384
rect 1820 7375 1822 7384
rect 3148 7404 3200 7410
rect 1768 7346 1820 7352
rect 3148 7346 3200 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 6736 7404 6788 7410
rect 7288 7404 7340 7410
rect 6788 7364 6868 7392
rect 6736 7346 6788 7352
rect 848 6860 900 6866
rect 848 6802 900 6808
rect 3160 6186 3188 7346
rect 4632 6225 4660 7346
rect 6423 7100 6731 7109
rect 6423 7098 6429 7100
rect 6485 7098 6509 7100
rect 6565 7098 6589 7100
rect 6645 7098 6669 7100
rect 6725 7098 6731 7100
rect 6485 7046 6487 7098
rect 6667 7046 6669 7098
rect 6423 7044 6429 7046
rect 6485 7044 6509 7046
rect 6565 7044 6589 7046
rect 6645 7044 6669 7046
rect 6725 7044 6731 7046
rect 6423 7035 6731 7044
rect 6840 6322 6868 7364
rect 7288 7346 7340 7352
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 4618 6216 4674 6225
rect 3148 6180 3200 6186
rect 4618 6151 4674 6160
rect 3148 6122 3200 6128
rect 6423 6012 6731 6021
rect 6423 6010 6429 6012
rect 6485 6010 6509 6012
rect 6565 6010 6589 6012
rect 6645 6010 6669 6012
rect 6725 6010 6731 6012
rect 6485 5958 6487 6010
rect 6667 5958 6669 6010
rect 6423 5956 6429 5958
rect 6485 5956 6509 5958
rect 6565 5956 6589 5958
rect 6645 5956 6669 5958
rect 6725 5956 6731 5958
rect 6423 5947 6731 5956
rect 6423 4924 6731 4933
rect 6423 4922 6429 4924
rect 6485 4922 6509 4924
rect 6565 4922 6589 4924
rect 6645 4922 6669 4924
rect 6725 4922 6731 4924
rect 6485 4870 6487 4922
rect 6667 4870 6669 4922
rect 6423 4868 6429 4870
rect 6485 4868 6509 4870
rect 6565 4868 6589 4870
rect 6645 4868 6669 4870
rect 6725 4868 6731 4870
rect 6423 4859 6731 4868
rect 7300 4826 7328 7346
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8312 6662 8340 7210
rect 8680 7206 8708 7414
rect 9876 7410 9904 7686
rect 10428 7528 10456 9840
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10508 7540 10560 7546
rect 10428 7500 10508 7528
rect 10508 7482 10560 7488
rect 10796 7410 10824 8026
rect 11060 7540 11112 7546
rect 11164 7528 11192 9840
rect 11900 8514 11928 9840
rect 11808 8486 11928 8514
rect 11702 7848 11758 7857
rect 11702 7783 11758 7792
rect 11112 7500 11192 7528
rect 11060 7482 11112 7488
rect 11716 7478 11744 7783
rect 11808 7528 11836 8486
rect 11896 7644 12204 7653
rect 11896 7642 11902 7644
rect 11958 7642 11982 7644
rect 12038 7642 12062 7644
rect 12118 7642 12142 7644
rect 12198 7642 12204 7644
rect 11958 7590 11960 7642
rect 12140 7590 12142 7642
rect 11896 7588 11902 7590
rect 11958 7588 11982 7590
rect 12038 7588 12062 7590
rect 12118 7588 12142 7590
rect 12198 7588 12204 7590
rect 11896 7579 12204 7588
rect 12636 7546 12664 9840
rect 13372 9738 13400 9840
rect 13464 9738 13492 9846
rect 13372 9710 13492 9738
rect 13740 8242 13768 9846
rect 14094 9840 14150 10000
rect 14830 9840 14886 10000
rect 15566 9840 15622 10000
rect 16302 9840 16358 10000
rect 17038 9840 17094 10000
rect 17774 9840 17830 10000
rect 18510 9840 18566 10000
rect 19246 9840 19302 10000
rect 19982 9840 20038 10000
rect 20718 9840 20774 10000
rect 21454 9840 21510 10000
rect 22190 9840 22246 10000
rect 22926 9840 22982 10000
rect 23032 9846 23244 9874
rect 13740 8214 13860 8242
rect 13832 7546 13860 8214
rect 14108 7546 14136 9840
rect 14844 8514 14872 9840
rect 14844 8486 15056 8514
rect 15028 7546 15056 8486
rect 15580 7546 15608 9840
rect 11888 7540 11940 7546
rect 11808 7500 11888 7528
rect 11888 7482 11940 7488
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 15108 7404 15160 7410
rect 16316 7392 16344 9840
rect 17052 7410 17080 9840
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 16488 7404 16540 7410
rect 16316 7364 16488 7392
rect 15108 7346 15160 7352
rect 16488 7346 16540 7352
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8404 5030 8432 7142
rect 9140 7002 9168 7346
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 10888 5098 10916 7278
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7930 4584 7986 4593
rect 7930 4519 7986 4528
rect 10324 4548 10376 4554
rect 6423 3836 6731 3845
rect 6423 3834 6429 3836
rect 6485 3834 6509 3836
rect 6565 3834 6589 3836
rect 6645 3834 6669 3836
rect 6725 3834 6731 3836
rect 6485 3782 6487 3834
rect 6667 3782 6669 3834
rect 6423 3780 6429 3782
rect 6485 3780 6509 3782
rect 6565 3780 6589 3782
rect 6645 3780 6669 3782
rect 6725 3780 6731 3782
rect 6423 3771 6731 3780
rect 6826 2816 6882 2825
rect 6423 2748 6731 2757
rect 6826 2751 6882 2760
rect 6423 2746 6429 2748
rect 6485 2746 6509 2748
rect 6565 2746 6589 2748
rect 6645 2746 6669 2748
rect 6725 2746 6731 2748
rect 6485 2694 6487 2746
rect 6667 2694 6669 2746
rect 6423 2692 6429 2694
rect 6485 2692 6509 2694
rect 6565 2692 6589 2694
rect 6645 2692 6669 2694
rect 6725 2692 6731 2694
rect 6423 2683 6731 2692
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6748 2530 6776 2586
rect 6840 2530 6868 2751
rect 6748 2502 6868 2530
rect 5632 2440 5684 2446
rect 5908 2440 5960 2446
rect 5684 2400 5764 2428
rect 5632 2382 5684 2388
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5644 1698 5672 2246
rect 5632 1692 5684 1698
rect 5632 1634 5684 1640
rect 5736 160 5764 2400
rect 6276 2440 6328 2446
rect 5960 2400 6040 2428
rect 5908 2382 5960 2388
rect 6012 160 6040 2400
rect 6276 2382 6328 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 6288 160 6316 2382
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6380 82 6408 2382
rect 6550 82 6606 160
rect 6380 54 6606 82
rect 6656 82 6684 2382
rect 6826 82 6882 160
rect 6656 54 6882 82
rect 6932 82 6960 2382
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1057 7144 2246
rect 7102 1048 7158 1057
rect 7102 983 7158 992
rect 7102 82 7158 160
rect 6932 54 7158 82
rect 7208 82 7236 2382
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7392 1698 7420 2246
rect 7380 1692 7432 1698
rect 7380 1634 7432 1640
rect 7378 82 7434 160
rect 7208 54 7434 82
rect 7484 82 7512 2382
rect 7654 82 7710 160
rect 7484 54 7710 82
rect 7760 82 7788 2382
rect 7944 2310 7972 4519
rect 10324 4490 10376 4496
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 8482 3496 8538 3505
rect 8482 3431 8538 3440
rect 8496 2446 8524 3431
rect 8758 3088 8814 3097
rect 8758 3023 8814 3032
rect 9128 3052 9180 3058
rect 8772 2446 8800 3023
rect 9128 2994 9180 3000
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7930 82 7986 160
rect 7760 54 7986 82
rect 8036 82 8064 2382
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8220 2106 8248 2246
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 8206 82 8262 160
rect 8036 54 8262 82
rect 8312 82 8340 2382
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 2106 8432 2246
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8482 82 8538 160
rect 8312 54 8538 82
rect 8588 82 8616 2382
rect 8758 82 8814 160
rect 8588 54 8814 82
rect 6550 0 6606 54
rect 6826 0 6882 54
rect 7102 0 7158 54
rect 7378 0 7434 54
rect 7654 0 7710 54
rect 7930 0 7986 54
rect 8206 0 8262 54
rect 8482 0 8538 54
rect 8758 0 8814 54
rect 9034 82 9090 160
rect 9140 82 9168 2994
rect 9402 2952 9458 2961
rect 9402 2887 9458 2896
rect 9416 2530 9444 2887
rect 9692 2650 9720 4082
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 9416 2502 9536 2530
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1834 9260 2246
rect 9220 1828 9272 1834
rect 9220 1770 9272 1776
rect 9324 160 9352 2314
rect 9034 54 9168 82
rect 9034 0 9090 54
rect 9310 0 9366 160
rect 9416 82 9444 2382
rect 9508 2310 9536 2502
rect 9600 2417 9628 2586
rect 9968 2553 9996 2586
rect 10232 2576 10284 2582
rect 9954 2544 10010 2553
rect 10232 2518 10284 2524
rect 9954 2479 10010 2488
rect 9680 2440 9732 2446
rect 9586 2408 9642 2417
rect 9680 2382 9732 2388
rect 9586 2343 9642 2352
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9586 82 9642 160
rect 9416 54 9642 82
rect 9692 82 9720 2382
rect 10140 2372 10192 2378
rect 10140 2314 10192 2320
rect 10152 160 10180 2314
rect 10244 1737 10272 2518
rect 10230 1728 10286 1737
rect 10336 1698 10364 4490
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10704 2446 10732 4014
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 10230 1663 10286 1672
rect 10324 1692 10376 1698
rect 10324 1634 10376 1640
rect 10428 160 10456 2382
rect 9862 82 9918 160
rect 9692 54 9918 82
rect 9586 0 9642 54
rect 9862 0 9918 54
rect 10138 0 10194 160
rect 10414 0 10470 160
rect 10520 82 10548 2382
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10612 1698 10640 2246
rect 10600 1692 10652 1698
rect 10600 1634 10652 1640
rect 10690 82 10746 160
rect 10520 54 10746 82
rect 10796 82 10824 2382
rect 10888 2106 10916 4422
rect 10980 3738 11008 7346
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 11896 6556 12204 6565
rect 11896 6554 11902 6556
rect 11958 6554 11982 6556
rect 12038 6554 12062 6556
rect 12118 6554 12142 6556
rect 12198 6554 12204 6556
rect 11958 6502 11960 6554
rect 12140 6502 12142 6554
rect 11896 6500 11902 6502
rect 11958 6500 11982 6502
rect 12038 6500 12062 6502
rect 12118 6500 12142 6502
rect 12198 6500 12204 6502
rect 11896 6491 12204 6500
rect 11896 5468 12204 5477
rect 11896 5466 11902 5468
rect 11958 5466 11982 5468
rect 12038 5466 12062 5468
rect 12118 5466 12142 5468
rect 12198 5466 12204 5468
rect 11958 5414 11960 5466
rect 12140 5414 12142 5466
rect 11896 5412 11902 5414
rect 11958 5412 11982 5414
rect 12038 5412 12062 5414
rect 12118 5412 12142 5414
rect 12198 5412 12204 5414
rect 11896 5403 12204 5412
rect 11896 4380 12204 4389
rect 11896 4378 11902 4380
rect 11958 4378 11982 4380
rect 12038 4378 12062 4380
rect 12118 4378 12142 4380
rect 12198 4378 12204 4380
rect 11958 4326 11960 4378
rect 12140 4326 12142 4378
rect 11896 4324 11902 4326
rect 11958 4324 11982 4326
rect 12038 4324 12062 4326
rect 12118 4324 12142 4326
rect 12198 4324 12204 4326
rect 11896 4315 12204 4324
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11072 2582 11100 4150
rect 11334 4040 11390 4049
rect 11334 3975 11390 3984
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 11256 2514 11284 3334
rect 11348 2582 11376 3975
rect 11896 3292 12204 3301
rect 11896 3290 11902 3292
rect 11958 3290 11982 3292
rect 12038 3290 12062 3292
rect 12118 3290 12142 3292
rect 12198 3290 12204 3292
rect 11958 3238 11960 3290
rect 12140 3238 12142 3290
rect 11896 3236 11902 3238
rect 11958 3236 11982 3238
rect 12038 3236 12062 3238
rect 12118 3236 12142 3238
rect 12198 3236 12204 3238
rect 11896 3227 12204 3236
rect 13188 2650 13216 7278
rect 13280 2650 13308 7346
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13358 3632 13414 3641
rect 13358 3567 13414 3576
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11900 2502 12388 2530
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11520 2440 11572 2446
rect 11572 2400 11836 2428
rect 11520 2382 11572 2388
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10966 82 11022 160
rect 10796 54 11022 82
rect 11072 82 11100 2382
rect 11440 1306 11468 2382
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11716 1630 11744 2246
rect 11704 1624 11756 1630
rect 11704 1566 11756 1572
rect 11440 1278 11560 1306
rect 11532 160 11560 1278
rect 11808 160 11836 2400
rect 11900 2378 11928 2502
rect 11980 2440 12032 2446
rect 12032 2400 12296 2428
rect 11980 2382 12032 2388
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11896 2204 12204 2213
rect 11896 2202 11902 2204
rect 11958 2202 11982 2204
rect 12038 2202 12062 2204
rect 12118 2202 12142 2204
rect 12198 2202 12204 2204
rect 11958 2150 11960 2202
rect 12140 2150 12142 2202
rect 11896 2148 11902 2150
rect 11958 2148 11982 2150
rect 12038 2148 12062 2150
rect 12118 2148 12142 2150
rect 12198 2148 12204 2150
rect 11896 2139 12204 2148
rect 12268 1306 12296 2400
rect 12084 1278 12296 1306
rect 12084 160 12112 1278
rect 12360 160 12388 2502
rect 12532 2440 12584 2446
rect 12808 2440 12860 2446
rect 12584 2400 12664 2428
rect 12532 2382 12584 2388
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12544 1766 12572 2246
rect 12532 1760 12584 1766
rect 12532 1702 12584 1708
rect 12636 160 12664 2400
rect 12860 2400 12940 2428
rect 12808 2382 12860 2388
rect 12912 160 12940 2400
rect 13004 2281 13032 2586
rect 13372 2530 13400 3567
rect 13740 3194 13768 4558
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13556 2774 13584 2994
rect 13280 2502 13400 2530
rect 13464 2746 13584 2774
rect 13280 2446 13308 2502
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13084 2304 13136 2310
rect 12990 2272 13046 2281
rect 13084 2246 13136 2252
rect 12990 2207 13046 2216
rect 13096 1873 13124 2246
rect 13082 1864 13138 1873
rect 13082 1799 13138 1808
rect 13188 160 13216 2382
rect 13372 1698 13400 2382
rect 13360 1692 13412 1698
rect 13360 1634 13412 1640
rect 13464 160 13492 2746
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13728 2440 13780 2446
rect 13780 2400 13860 2428
rect 13728 2382 13780 2388
rect 13648 1306 13676 2382
rect 13648 1278 13768 1306
rect 13740 160 13768 1278
rect 11242 82 11298 160
rect 11072 54 11298 82
rect 10690 0 10746 54
rect 10966 0 11022 54
rect 11242 0 11298 54
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 13832 82 13860 2400
rect 14292 2310 14320 7346
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 5710 14504 7142
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14554 4176 14610 4185
rect 14554 4111 14610 4120
rect 14462 3224 14518 3233
rect 14568 3194 14596 4111
rect 14462 3159 14518 3168
rect 14556 3188 14608 3194
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14200 2009 14228 2246
rect 14186 2000 14242 2009
rect 14186 1935 14242 1944
rect 13912 1556 13964 1562
rect 13912 1498 13964 1504
rect 13924 1222 13952 1498
rect 13912 1216 13964 1222
rect 13912 1158 13964 1164
rect 14002 82 14058 160
rect 13832 54 14058 82
rect 14002 0 14058 54
rect 14278 82 14334 160
rect 14384 82 14412 2994
rect 14476 2825 14504 3159
rect 14556 3130 14608 3136
rect 14556 2848 14608 2854
rect 14462 2816 14518 2825
rect 14556 2790 14608 2796
rect 14462 2751 14518 2760
rect 14464 2576 14516 2582
rect 14464 2518 14516 2524
rect 14476 2106 14504 2518
rect 14568 2378 14596 2790
rect 14660 2582 14688 7346
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 15120 2514 15148 7346
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15566 3360 15622 3369
rect 15566 3295 15622 3304
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14660 1902 14688 2382
rect 14648 1896 14700 1902
rect 14648 1838 14700 1844
rect 14752 1358 14780 2382
rect 15212 2258 15240 2382
rect 15120 2230 15240 2258
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 15120 1290 15148 2230
rect 15304 2106 15332 2382
rect 15396 2106 15424 2450
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15580 1834 15608 3295
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15568 1828 15620 1834
rect 15568 1770 15620 1776
rect 15200 1624 15252 1630
rect 15200 1566 15252 1572
rect 15108 1284 15160 1290
rect 15108 1226 15160 1232
rect 15212 1193 15240 1566
rect 15198 1184 15254 1193
rect 15198 1119 15254 1128
rect 15672 160 15700 2926
rect 15948 2514 15976 6802
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16408 2582 16436 2790
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 15936 2508 15988 2514
rect 15936 2450 15988 2456
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 16396 2440 16448 2446
rect 16396 2382 16448 2388
rect 14278 54 14412 82
rect 14278 0 14334 54
rect 14554 0 14610 160
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15856 82 15884 2382
rect 15934 82 15990 160
rect 15856 54 15990 82
rect 15934 0 15990 54
rect 16210 82 16266 160
rect 16408 82 16436 2382
rect 16500 160 16528 3470
rect 16592 2774 16620 3606
rect 16684 2938 16712 6394
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16776 3670 16804 3946
rect 16764 3664 16816 3670
rect 16764 3606 16816 3612
rect 16868 3058 16896 6190
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16684 2910 16896 2938
rect 16592 2746 16804 2774
rect 16776 160 16804 2746
rect 16868 2514 16896 2910
rect 16960 2650 16988 3402
rect 17052 3074 17080 6734
rect 17144 3194 17172 7142
rect 17236 6730 17264 7822
rect 17788 7392 17816 9840
rect 18328 8152 18380 8158
rect 18328 8094 18380 8100
rect 17868 7404 17920 7410
rect 17788 7364 17868 7392
rect 17868 7346 17920 7352
rect 17866 7304 17922 7313
rect 17788 7262 17866 7290
rect 17370 7100 17678 7109
rect 17370 7098 17376 7100
rect 17432 7098 17456 7100
rect 17512 7098 17536 7100
rect 17592 7098 17616 7100
rect 17672 7098 17678 7100
rect 17432 7046 17434 7098
rect 17614 7046 17616 7098
rect 17370 7044 17376 7046
rect 17432 7044 17456 7046
rect 17512 7044 17536 7046
rect 17592 7044 17616 7046
rect 17672 7044 17678 7046
rect 17370 7035 17678 7044
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17370 6012 17678 6021
rect 17370 6010 17376 6012
rect 17432 6010 17456 6012
rect 17512 6010 17536 6012
rect 17592 6010 17616 6012
rect 17672 6010 17678 6012
rect 17432 5958 17434 6010
rect 17614 5958 17616 6010
rect 17370 5956 17376 5958
rect 17432 5956 17456 5958
rect 17512 5956 17536 5958
rect 17592 5956 17616 5958
rect 17672 5956 17678 5958
rect 17370 5947 17678 5956
rect 17370 4924 17678 4933
rect 17370 4922 17376 4924
rect 17432 4922 17456 4924
rect 17512 4922 17536 4924
rect 17592 4922 17616 4924
rect 17672 4922 17678 4924
rect 17432 4870 17434 4922
rect 17614 4870 17616 4922
rect 17370 4868 17376 4870
rect 17432 4868 17456 4870
rect 17512 4868 17536 4870
rect 17592 4868 17616 4870
rect 17672 4868 17678 4870
rect 17370 4859 17678 4868
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17236 3194 17264 4218
rect 17370 3836 17678 3845
rect 17370 3834 17376 3836
rect 17432 3834 17456 3836
rect 17512 3834 17536 3836
rect 17592 3834 17616 3836
rect 17672 3834 17678 3836
rect 17432 3782 17434 3834
rect 17614 3782 17616 3834
rect 17370 3780 17376 3782
rect 17432 3780 17456 3782
rect 17512 3780 17536 3782
rect 17592 3780 17616 3782
rect 17672 3780 17678 3782
rect 17370 3771 17678 3780
rect 17788 3618 17816 7262
rect 17866 7239 17922 7248
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 18064 6361 18092 7142
rect 18050 6352 18106 6361
rect 18050 6287 18106 6296
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17880 3670 17908 5102
rect 18064 4026 18092 5714
rect 18234 5128 18290 5137
rect 17972 3998 18092 4026
rect 18156 5086 18234 5114
rect 17696 3590 17816 3618
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17696 3534 17724 3590
rect 17684 3528 17736 3534
rect 17868 3528 17920 3534
rect 17684 3470 17736 3476
rect 17788 3488 17868 3516
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 17696 3126 17724 3334
rect 17684 3120 17736 3126
rect 17052 3046 17356 3074
rect 17684 3062 17736 3068
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17144 2446 17172 2790
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 16856 2372 16908 2378
rect 16908 2332 17080 2360
rect 16856 2314 16908 2320
rect 17052 160 17080 2332
rect 17236 1578 17264 2926
rect 17328 2854 17356 3046
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17370 2748 17678 2757
rect 17370 2746 17376 2748
rect 17432 2746 17456 2748
rect 17512 2746 17536 2748
rect 17592 2746 17616 2748
rect 17672 2746 17678 2748
rect 17432 2694 17434 2746
rect 17614 2694 17616 2746
rect 17370 2692 17376 2694
rect 17432 2692 17456 2694
rect 17512 2692 17536 2694
rect 17592 2692 17616 2694
rect 17672 2692 17678 2694
rect 17370 2683 17678 2692
rect 17236 1550 17356 1578
rect 17328 160 17356 1550
rect 16210 54 16436 82
rect 16210 0 16266 54
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 82 17646 160
rect 17788 82 17816 3488
rect 17868 3470 17920 3476
rect 17972 3482 18000 3998
rect 17972 3454 18092 3482
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17880 160 17908 3334
rect 17972 3194 18000 3334
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17972 2825 18000 2858
rect 17958 2816 18014 2825
rect 17958 2751 18014 2760
rect 18064 2514 18092 3454
rect 18156 3194 18184 5086
rect 18234 5063 18290 5072
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18248 3126 18276 3334
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 1902 18092 2246
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 18156 160 18184 2994
rect 18340 2922 18368 8094
rect 18524 7410 18552 9840
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18432 2836 18460 3470
rect 18524 2990 18552 3878
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18616 2836 18644 7686
rect 19260 7546 19288 9840
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19352 7546 19472 7562
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 19340 7540 19472 7546
rect 19392 7534 19472 7540
rect 19340 7482 19392 7488
rect 19168 7426 19196 7482
rect 19168 7398 19380 7426
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18788 4208 18840 4214
rect 18788 4150 18840 4156
rect 18800 3738 18828 4150
rect 18892 4010 18920 6326
rect 18970 4312 19026 4321
rect 18970 4247 19026 4256
rect 18984 4146 19012 4247
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19076 4010 19104 7278
rect 19352 5914 19380 7398
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 19260 4298 19288 5646
rect 19260 4270 19380 4298
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 19064 4004 19116 4010
rect 19064 3946 19116 3952
rect 19260 3913 19288 4082
rect 19246 3904 19302 3913
rect 19246 3839 19302 3848
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18696 2848 18748 2854
rect 18432 2808 18552 2836
rect 18616 2808 18696 2836
rect 18326 2680 18382 2689
rect 18326 2615 18328 2624
rect 18380 2615 18382 2624
rect 18328 2586 18380 2592
rect 18524 2530 18552 2808
rect 18696 2790 18748 2796
rect 18432 2502 18552 2530
rect 18432 160 18460 2502
rect 18512 2440 18564 2446
rect 18510 2408 18512 2417
rect 18604 2440 18656 2446
rect 18564 2408 18566 2417
rect 18604 2382 18656 2388
rect 18510 2343 18566 2352
rect 18616 1426 18644 2382
rect 18800 1698 18828 3402
rect 18880 3392 18932 3398
rect 19064 3392 19116 3398
rect 18880 3334 18932 3340
rect 18984 3352 19064 3380
rect 18892 3126 18920 3334
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18880 2440 18932 2446
rect 18880 2382 18932 2388
rect 18788 1692 18840 1698
rect 18788 1634 18840 1640
rect 18892 1562 18920 2382
rect 18984 2122 19012 3352
rect 19064 3334 19116 3340
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19076 2689 19104 2926
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 19168 2825 19196 2858
rect 19154 2816 19210 2825
rect 19154 2751 19210 2760
rect 19352 2689 19380 4270
rect 19444 4010 19472 7534
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19536 3482 19564 7890
rect 19800 7812 19852 7818
rect 19800 7754 19852 7760
rect 19812 7546 19840 7754
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19062 2680 19118 2689
rect 19062 2615 19118 2624
rect 19338 2680 19394 2689
rect 19338 2615 19394 2624
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19352 2281 19380 2382
rect 19338 2272 19394 2281
rect 19338 2207 19394 2216
rect 18984 2094 19288 2122
rect 19156 1964 19208 1970
rect 19156 1906 19208 1912
rect 18880 1556 18932 1562
rect 18880 1498 18932 1504
rect 18604 1420 18656 1426
rect 18604 1362 18656 1368
rect 19168 1329 19196 1906
rect 19154 1320 19210 1329
rect 19154 1255 19210 1264
rect 18984 190 19104 218
rect 18984 160 19012 190
rect 17590 54 17816 82
rect 17590 0 17646 54
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 82 18750 160
rect 18786 96 18842 105
rect 18694 54 18786 82
rect 18694 0 18750 54
rect 18786 31 18842 40
rect 18970 0 19026 160
rect 19076 105 19104 190
rect 19260 160 19288 2094
rect 19062 96 19118 105
rect 19062 31 19118 40
rect 19246 0 19302 160
rect 19444 82 19472 3470
rect 19536 3454 19656 3482
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19536 3194 19564 3334
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19628 2990 19656 3454
rect 19720 2990 19748 6054
rect 19812 3738 19840 7278
rect 19904 7206 19932 7482
rect 19996 7410 20024 9840
rect 20536 8220 20588 8226
rect 20536 8162 20588 8168
rect 20258 7984 20314 7993
rect 20258 7919 20314 7928
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 20272 3738 20300 7919
rect 20548 7410 20576 8162
rect 20732 7410 20760 9840
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20364 3534 20392 7142
rect 21008 3738 21036 8026
rect 21468 7410 21496 9840
rect 22204 7410 22232 9840
rect 22940 9738 22968 9840
rect 23032 9738 23060 9846
rect 22940 9710 23060 9738
rect 22843 7644 23151 7653
rect 22843 7642 22849 7644
rect 22905 7642 22929 7644
rect 22985 7642 23009 7644
rect 23065 7642 23089 7644
rect 23145 7642 23151 7644
rect 22905 7590 22907 7642
rect 23087 7590 23089 7642
rect 22843 7588 22849 7590
rect 22905 7588 22929 7590
rect 22985 7588 23009 7590
rect 23065 7588 23089 7590
rect 23145 7588 23151 7590
rect 22843 7579 23151 7588
rect 23216 7410 23244 9846
rect 23662 9840 23718 10000
rect 24398 9840 24454 10000
rect 25134 9840 25190 10000
rect 25870 9840 25926 10000
rect 26606 9840 26662 10000
rect 27342 9840 27398 10000
rect 28078 9840 28134 10000
rect 28814 9840 28870 10000
rect 29550 9840 29606 10000
rect 30286 9840 30342 10000
rect 31022 9840 31078 10000
rect 31758 9840 31814 10000
rect 32494 9840 32550 10000
rect 33230 9840 33286 10000
rect 33966 9840 34022 10000
rect 34072 9846 34284 9874
rect 23480 8016 23532 8022
rect 23480 7958 23532 7964
rect 23492 7546 23520 7958
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23676 7410 23704 9840
rect 24412 7410 24440 9840
rect 24950 7848 25006 7857
rect 24950 7783 25006 7792
rect 24964 7546 24992 7783
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25148 7410 25176 9840
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25700 7546 25728 7822
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25884 7410 25912 9840
rect 26620 7410 26648 9840
rect 27356 7410 27384 9840
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27804 7472 27856 7478
rect 27804 7414 27856 7420
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 22284 7200 22336 7206
rect 22284 7142 22336 7148
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 21100 3534 21128 7142
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21836 4214 21864 4558
rect 21824 4208 21876 4214
rect 21824 4150 21876 4156
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 20076 3528 20128 3534
rect 19904 3488 20076 3516
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19720 1306 19748 2450
rect 19812 2446 19840 3334
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19904 1970 19932 3488
rect 20076 3470 20128 3476
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19996 3233 20024 3334
rect 19982 3224 20038 3233
rect 19982 3159 20038 3168
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19996 2650 20024 2926
rect 20260 2848 20312 2854
rect 20088 2796 20260 2802
rect 20088 2790 20312 2796
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20088 2774 20300 2790
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19892 1964 19944 1970
rect 19892 1906 19944 1912
rect 19720 1278 19840 1306
rect 19812 160 19840 1278
rect 20088 160 20116 2774
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20364 160 20392 2450
rect 20640 160 20668 2790
rect 20824 2650 20852 3470
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20916 2774 20944 3334
rect 20916 2746 21036 2774
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 19522 82 19578 160
rect 19444 54 19578 82
rect 19522 0 19578 54
rect 19798 0 19854 160
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20732 82 20760 2450
rect 21008 1970 21036 2746
rect 21192 2446 21220 3878
rect 21468 3194 21496 3878
rect 21560 3738 21588 3946
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21456 3188 21508 3194
rect 21456 3130 21508 3136
rect 21560 2961 21588 3470
rect 21546 2952 21602 2961
rect 21546 2887 21602 2896
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 20996 1964 21048 1970
rect 20996 1906 21048 1912
rect 20902 82 20958 160
rect 20732 54 20958 82
rect 20902 0 20958 54
rect 21178 82 21234 160
rect 21376 82 21404 2790
rect 21652 2553 21680 4082
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 21732 3392 21784 3398
rect 22008 3392 22060 3398
rect 21732 3334 21784 3340
rect 21928 3352 22008 3380
rect 21744 3194 21772 3334
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21638 2544 21694 2553
rect 21836 2514 21864 2790
rect 21638 2479 21694 2488
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 21548 2440 21600 2446
rect 21548 2382 21600 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 21468 160 21496 2314
rect 21560 1222 21588 2382
rect 21640 2372 21692 2378
rect 21640 2314 21692 2320
rect 21548 1216 21600 1222
rect 21548 1158 21600 1164
rect 21178 54 21404 82
rect 21178 0 21234 54
rect 21454 0 21510 160
rect 21652 82 21680 2314
rect 21928 2310 21956 3352
rect 22008 3334 22060 3340
rect 22006 3088 22062 3097
rect 22006 3023 22008 3032
rect 22060 3023 22062 3032
rect 22008 2994 22060 3000
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22020 160 22048 2790
rect 22112 2446 22140 3878
rect 22296 3670 22324 7142
rect 22572 6934 22600 7346
rect 22560 6928 22612 6934
rect 22560 6870 22612 6876
rect 22843 6556 23151 6565
rect 22843 6554 22849 6556
rect 22905 6554 22929 6556
rect 22985 6554 23009 6556
rect 23065 6554 23089 6556
rect 23145 6554 23151 6556
rect 22905 6502 22907 6554
rect 23087 6502 23089 6554
rect 22843 6500 22849 6502
rect 22905 6500 22929 6502
rect 22985 6500 23009 6502
rect 23065 6500 23089 6502
rect 23145 6500 23151 6502
rect 22843 6491 23151 6500
rect 22843 5468 23151 5477
rect 22843 5466 22849 5468
rect 22905 5466 22929 5468
rect 22985 5466 23009 5468
rect 23065 5466 23089 5468
rect 23145 5466 23151 5468
rect 22905 5414 22907 5466
rect 23087 5414 23089 5466
rect 22843 5412 22849 5414
rect 22905 5412 22929 5414
rect 22985 5412 23009 5414
rect 23065 5412 23089 5414
rect 23145 5412 23151 5414
rect 22843 5403 23151 5412
rect 23308 5234 23336 7346
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22376 3936 22428 3942
rect 22376 3878 22428 3884
rect 22284 3664 22336 3670
rect 22284 3606 22336 3612
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22284 3528 22336 3534
rect 22388 3516 22416 3878
rect 22336 3488 22416 3516
rect 22468 3528 22520 3534
rect 22284 3470 22336 3476
rect 22468 3470 22520 3476
rect 22204 3369 22232 3470
rect 22284 3392 22336 3398
rect 22190 3360 22246 3369
rect 22284 3334 22336 3340
rect 22190 3295 22246 3304
rect 22296 3194 22324 3334
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22480 3058 22508 3470
rect 22664 3058 22692 4422
rect 22843 4380 23151 4389
rect 22843 4378 22849 4380
rect 22905 4378 22929 4380
rect 22985 4378 23009 4380
rect 23065 4378 23089 4380
rect 23145 4378 23151 4380
rect 22905 4326 22907 4378
rect 23087 4326 23089 4378
rect 22843 4324 22849 4326
rect 22905 4324 22929 4326
rect 22985 4324 23009 4326
rect 23065 4324 23089 4326
rect 23145 4324 23151 4326
rect 22843 4315 23151 4324
rect 23308 4010 23336 4490
rect 23112 4004 23164 4010
rect 23112 3946 23164 3952
rect 23296 4004 23348 4010
rect 23296 3946 23348 3952
rect 23124 3398 23152 3946
rect 23584 3670 23612 7210
rect 23756 7200 23808 7206
rect 23756 7142 23808 7148
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23676 3670 23704 6938
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23204 3528 23256 3534
rect 23202 3496 23204 3505
rect 23256 3496 23258 3505
rect 23202 3431 23258 3440
rect 22744 3392 22796 3398
rect 22744 3334 22796 3340
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22480 2922 22692 2938
rect 22480 2916 22704 2922
rect 22480 2910 22652 2916
rect 22100 2440 22152 2446
rect 22100 2382 22152 2388
rect 22376 2372 22428 2378
rect 22376 2314 22428 2320
rect 21730 82 21786 160
rect 21652 54 21786 82
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22282 82 22338 160
rect 22388 82 22416 2314
rect 22480 1737 22508 2910
rect 22652 2858 22704 2864
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22466 1728 22522 1737
rect 22466 1663 22522 1672
rect 22572 160 22600 2790
rect 22756 2774 22784 3334
rect 22843 3292 23151 3301
rect 22843 3290 22849 3292
rect 22905 3290 22929 3292
rect 22985 3290 23009 3292
rect 23065 3290 23089 3292
rect 23145 3290 23151 3292
rect 22905 3238 22907 3290
rect 23087 3238 23089 3290
rect 22843 3236 22849 3238
rect 22905 3236 22929 3238
rect 22985 3236 23009 3238
rect 23065 3236 23089 3238
rect 23145 3236 23151 3238
rect 22843 3227 23151 3236
rect 23388 2848 23440 2854
rect 22664 2746 22784 2774
rect 23308 2808 23388 2836
rect 22664 1601 22692 2746
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 22836 2304 22888 2310
rect 22756 2264 22836 2292
rect 22650 1592 22706 1601
rect 22650 1527 22706 1536
rect 22282 54 22416 82
rect 22282 0 22338 54
rect 22558 0 22614 160
rect 22756 82 22784 2264
rect 22836 2246 22888 2252
rect 22843 2204 23151 2213
rect 22843 2202 22849 2204
rect 22905 2202 22929 2204
rect 22985 2202 23009 2204
rect 23065 2202 23089 2204
rect 23145 2202 23151 2204
rect 22905 2150 22907 2202
rect 23087 2150 23089 2202
rect 22843 2148 22849 2150
rect 22905 2148 22929 2150
rect 22985 2148 23009 2150
rect 23065 2148 23089 2150
rect 23145 2148 23151 2150
rect 22843 2139 23151 2148
rect 23216 1902 23244 2586
rect 23204 1896 23256 1902
rect 23204 1838 23256 1844
rect 22834 82 22890 160
rect 22756 54 22890 82
rect 22834 0 22890 54
rect 23110 82 23166 160
rect 23308 82 23336 2808
rect 23388 2790 23440 2796
rect 23492 2774 23520 3606
rect 23768 3194 23796 7142
rect 24030 4584 24086 4593
rect 24030 4519 24086 4528
rect 24044 3534 24072 4519
rect 24400 4004 24452 4010
rect 24400 3946 24452 3952
rect 24032 3528 24084 3534
rect 24032 3470 24084 3476
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24124 3460 24176 3466
rect 24124 3402 24176 3408
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24044 3097 24072 3130
rect 24030 3088 24086 3097
rect 24030 3023 24086 3032
rect 23492 2746 23612 2774
rect 23584 2446 23612 2746
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23572 2304 23624 2310
rect 23400 2264 23572 2292
rect 23400 160 23428 2264
rect 23572 2246 23624 2252
rect 23664 2304 23716 2310
rect 24032 2304 24084 2310
rect 23664 2246 23716 2252
rect 23952 2264 24032 2292
rect 23676 160 23704 2246
rect 23952 160 23980 2264
rect 24032 2246 24084 2252
rect 24136 1426 24164 3402
rect 24216 2848 24268 2854
rect 24320 2836 24348 3470
rect 24412 3058 24440 3946
rect 24872 3670 24900 7142
rect 25056 5846 25084 7346
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 25044 5840 25096 5846
rect 25044 5782 25096 5788
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 24780 3516 24808 3606
rect 25148 3602 25176 7210
rect 25608 7002 25636 7346
rect 27344 7200 27396 7206
rect 27344 7142 27396 7148
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 27160 6928 27212 6934
rect 27160 6870 27212 6876
rect 26608 6656 26660 6662
rect 26608 6598 26660 6604
rect 25872 6316 25924 6322
rect 25872 6258 25924 6264
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25136 3596 25188 3602
rect 25136 3538 25188 3544
rect 25228 3528 25280 3534
rect 24780 3488 24900 3516
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24504 3194 24532 3334
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 24268 2808 24348 2836
rect 24492 2848 24544 2854
rect 24216 2790 24268 2796
rect 24492 2790 24544 2796
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 24124 1420 24176 1426
rect 24124 1362 24176 1368
rect 23110 54 23336 82
rect 23110 0 23166 54
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 82 24270 160
rect 24412 82 24440 2586
rect 24504 160 24532 2790
rect 24780 2417 24808 3334
rect 24872 2446 24900 3488
rect 25226 3496 25228 3505
rect 25280 3496 25282 3505
rect 25226 3431 25282 3440
rect 25044 3392 25096 3398
rect 25320 3392 25372 3398
rect 25096 3352 25268 3380
rect 25044 3334 25096 3340
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24860 2440 24912 2446
rect 24766 2408 24822 2417
rect 24860 2382 24912 2388
rect 24766 2343 24822 2352
rect 24952 2304 25004 2310
rect 24780 2264 24952 2292
rect 24780 160 24808 2264
rect 24952 2246 25004 2252
rect 25056 160 25084 2790
rect 25240 2446 25268 3352
rect 25320 3334 25372 3340
rect 25332 3194 25360 3334
rect 25424 3194 25452 3878
rect 25884 3670 25912 6258
rect 26516 4820 26568 4826
rect 26516 4762 26568 4768
rect 26528 4010 26556 4762
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26620 3670 26648 6598
rect 26790 6352 26846 6361
rect 26790 6287 26846 6296
rect 26804 4146 26832 6287
rect 26976 5092 27028 5098
rect 26976 5034 27028 5040
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 25872 3664 25924 3670
rect 25872 3606 25924 3612
rect 26608 3664 26660 3670
rect 26608 3606 26660 3612
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25700 3369 25728 3470
rect 25964 3392 26016 3398
rect 25686 3360 25742 3369
rect 25964 3334 26016 3340
rect 25686 3295 25742 3304
rect 25976 3194 26004 3334
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 25412 2916 25464 2922
rect 25412 2858 25464 2864
rect 25424 2446 25452 2858
rect 25596 2848 25648 2854
rect 25596 2790 25648 2796
rect 26056 2848 26108 2854
rect 26608 2848 26660 2854
rect 26056 2790 26108 2796
rect 26436 2808 26608 2836
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 24214 54 24440 82
rect 24214 0 24270 54
rect 24490 0 24546 160
rect 24766 0 24822 160
rect 25042 0 25098 160
rect 25318 82 25374 160
rect 25516 82 25544 2586
rect 25608 160 25636 2790
rect 25318 54 25544 82
rect 25318 0 25374 54
rect 25594 0 25650 160
rect 25870 82 25926 160
rect 26068 82 26096 2790
rect 26332 2372 26384 2378
rect 26160 2332 26332 2360
rect 26160 160 26188 2332
rect 26332 2314 26384 2320
rect 26436 160 26464 2808
rect 26608 2790 26660 2796
rect 26514 2680 26570 2689
rect 26514 2615 26516 2624
rect 26568 2615 26570 2624
rect 26516 2586 26568 2592
rect 26712 2553 26740 4082
rect 26988 3670 27016 5034
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 27080 3670 27108 4966
rect 27172 4826 27200 6870
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 26976 3664 27028 3670
rect 26976 3606 27028 3612
rect 27068 3664 27120 3670
rect 27068 3606 27120 3612
rect 26792 3460 26844 3466
rect 26792 3402 26844 3408
rect 26698 2544 26754 2553
rect 26698 2479 26754 2488
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26620 1698 26648 2382
rect 26804 1737 26832 3402
rect 27172 3194 27200 3878
rect 27356 3466 27384 7142
rect 27618 3632 27674 3641
rect 27816 3602 27844 7414
rect 27618 3567 27674 3576
rect 27712 3596 27764 3602
rect 27632 3534 27660 3567
rect 27712 3538 27764 3544
rect 27804 3596 27856 3602
rect 27804 3538 27856 3544
rect 27528 3528 27580 3534
rect 27526 3496 27528 3505
rect 27620 3528 27672 3534
rect 27580 3496 27582 3505
rect 27344 3460 27396 3466
rect 27620 3470 27672 3476
rect 27724 3482 27752 3538
rect 27724 3454 27844 3482
rect 27526 3431 27582 3440
rect 27344 3402 27396 3408
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 26976 2916 27028 2922
rect 26976 2858 27028 2864
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26790 1728 26846 1737
rect 26608 1692 26660 1698
rect 26790 1663 26846 1672
rect 26608 1634 26660 1640
rect 25870 54 26096 82
rect 25870 0 25926 54
rect 26146 0 26202 160
rect 26422 0 26478 160
rect 26698 82 26754 160
rect 26896 82 26924 2586
rect 26988 160 27016 2858
rect 27068 2372 27120 2378
rect 27068 2314 27120 2320
rect 27436 2372 27488 2378
rect 27436 2314 27488 2320
rect 27080 1970 27108 2314
rect 27160 2032 27212 2038
rect 27344 2032 27396 2038
rect 27212 1980 27344 1986
rect 27160 1974 27396 1980
rect 27068 1964 27120 1970
rect 27172 1958 27384 1974
rect 27068 1906 27120 1912
rect 27160 1624 27212 1630
rect 27160 1566 27212 1572
rect 27172 1426 27200 1566
rect 27160 1420 27212 1426
rect 27160 1362 27212 1368
rect 26698 54 26924 82
rect 26698 0 26754 54
rect 26974 0 27030 160
rect 27250 82 27306 160
rect 27448 82 27476 2314
rect 27540 160 27568 3130
rect 27724 3126 27752 3334
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27816 2774 27844 3454
rect 27632 2746 27844 2774
rect 27632 2417 27660 2746
rect 27908 2446 27936 7482
rect 28092 7410 28120 9840
rect 28828 8242 28856 9840
rect 28828 8214 29132 8242
rect 28998 7984 29054 7993
rect 28998 7919 29054 7928
rect 29012 7478 29040 7919
rect 29000 7472 29052 7478
rect 29000 7414 29052 7420
rect 29104 7410 29132 8214
rect 29276 7744 29328 7750
rect 29276 7686 29328 7692
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 29092 7404 29144 7410
rect 29092 7346 29144 7352
rect 29288 7342 29316 7686
rect 29564 7410 29592 9840
rect 29552 7404 29604 7410
rect 29552 7346 29604 7352
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 30300 7290 30328 9840
rect 30748 8220 30800 8226
rect 30748 8162 30800 8168
rect 30760 7478 30788 8162
rect 31036 7546 31064 9840
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 30748 7472 30800 7478
rect 30748 7414 30800 7420
rect 30838 7440 30894 7449
rect 30380 7404 30432 7410
rect 30838 7375 30894 7384
rect 30380 7346 30432 7352
rect 30392 7290 30420 7346
rect 29000 7268 29052 7274
rect 29000 7210 29052 7216
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28724 7200 28776 7206
rect 28776 7160 28856 7188
rect 28724 7142 28776 7148
rect 27988 6180 28040 6186
rect 27988 6122 28040 6128
rect 28000 3482 28028 6122
rect 28184 3516 28212 7142
rect 28317 7100 28625 7109
rect 28317 7098 28323 7100
rect 28379 7098 28403 7100
rect 28459 7098 28483 7100
rect 28539 7098 28563 7100
rect 28619 7098 28625 7100
rect 28379 7046 28381 7098
rect 28561 7046 28563 7098
rect 28317 7044 28323 7046
rect 28379 7044 28403 7046
rect 28459 7044 28483 7046
rect 28539 7044 28563 7046
rect 28619 7044 28625 7046
rect 28317 7035 28625 7044
rect 28317 6012 28625 6021
rect 28317 6010 28323 6012
rect 28379 6010 28403 6012
rect 28459 6010 28483 6012
rect 28539 6010 28563 6012
rect 28619 6010 28625 6012
rect 28379 5958 28381 6010
rect 28561 5958 28563 6010
rect 28317 5956 28323 5958
rect 28379 5956 28403 5958
rect 28459 5956 28483 5958
rect 28539 5956 28563 5958
rect 28619 5956 28625 5958
rect 28317 5947 28625 5956
rect 28317 4924 28625 4933
rect 28317 4922 28323 4924
rect 28379 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28625 4924
rect 28379 4870 28381 4922
rect 28561 4870 28563 4922
rect 28317 4868 28323 4870
rect 28379 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28625 4870
rect 28317 4859 28625 4868
rect 28317 3836 28625 3845
rect 28317 3834 28323 3836
rect 28379 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28625 3836
rect 28379 3782 28381 3834
rect 28561 3782 28563 3834
rect 28317 3780 28323 3782
rect 28379 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28625 3782
rect 28317 3771 28625 3780
rect 28722 3768 28778 3777
rect 28722 3703 28724 3712
rect 28776 3703 28778 3712
rect 28724 3674 28776 3680
rect 28828 3618 28856 7160
rect 28736 3590 28856 3618
rect 29012 3602 29040 7210
rect 29196 3602 29224 7278
rect 30300 7262 30420 7290
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29460 3664 29512 3670
rect 29460 3606 29512 3612
rect 29000 3596 29052 3602
rect 28264 3528 28316 3534
rect 28184 3488 28264 3516
rect 28000 3454 28120 3482
rect 28264 3470 28316 3476
rect 27988 3392 28040 3398
rect 28092 3380 28120 3454
rect 28172 3392 28224 3398
rect 28092 3352 28172 3380
rect 27988 3334 28040 3340
rect 28172 3334 28224 3340
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28000 2961 28028 3334
rect 28644 3194 28672 3334
rect 28632 3188 28684 3194
rect 28632 3130 28684 3136
rect 27986 2952 28042 2961
rect 27986 2887 28042 2896
rect 28448 2848 28500 2854
rect 28184 2808 28448 2836
rect 28080 2508 28132 2514
rect 28000 2468 28080 2496
rect 27896 2440 27948 2446
rect 27618 2408 27674 2417
rect 27896 2382 27948 2388
rect 27618 2343 27674 2352
rect 27250 54 27476 82
rect 27250 0 27306 54
rect 27526 0 27582 160
rect 27802 82 27858 160
rect 28000 82 28028 2468
rect 28080 2450 28132 2456
rect 27802 54 28028 82
rect 28078 82 28134 160
rect 28184 82 28212 2808
rect 28448 2790 28500 2796
rect 28317 2748 28625 2757
rect 28317 2746 28323 2748
rect 28379 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28625 2748
rect 28379 2694 28381 2746
rect 28561 2694 28563 2746
rect 28317 2692 28323 2694
rect 28379 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28625 2694
rect 28317 2683 28625 2692
rect 28632 2644 28684 2650
rect 28632 2586 28684 2592
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28552 2106 28580 2382
rect 28540 2100 28592 2106
rect 28540 2042 28592 2048
rect 28644 490 28672 2586
rect 28736 2446 28764 3590
rect 29000 3538 29052 3544
rect 29184 3596 29236 3602
rect 29184 3538 29236 3544
rect 28908 3392 28960 3398
rect 29184 3392 29236 3398
rect 28960 3352 29132 3380
rect 28908 3334 28960 3340
rect 28908 2848 28960 2854
rect 28828 2808 28908 2836
rect 28724 2440 28776 2446
rect 28724 2382 28776 2388
rect 28552 462 28672 490
rect 28078 54 28212 82
rect 28354 82 28410 160
rect 28552 82 28580 462
rect 28354 54 28580 82
rect 28630 82 28686 160
rect 28828 82 28856 2808
rect 28908 2790 28960 2796
rect 28998 2816 29054 2825
rect 28998 2751 29054 2760
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 28920 160 28948 2518
rect 29012 2378 29040 2751
rect 29104 2446 29132 3352
rect 29184 3334 29236 3340
rect 29196 3194 29224 3334
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29184 2916 29236 2922
rect 29184 2858 29236 2864
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 29000 2372 29052 2378
rect 29000 2314 29052 2320
rect 29000 2032 29052 2038
rect 28998 2000 29000 2009
rect 29052 2000 29054 2009
rect 28998 1935 29054 1944
rect 29196 160 29224 2858
rect 29472 2446 29500 3606
rect 29656 3534 29684 7142
rect 29826 6216 29882 6225
rect 29826 6151 29882 6160
rect 29840 3738 29868 6151
rect 30380 5908 30432 5914
rect 30380 5850 30432 5856
rect 30286 4040 30342 4049
rect 30286 3975 30342 3984
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30300 3534 30328 3975
rect 29644 3528 29696 3534
rect 29644 3470 29696 3476
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 30012 3392 30064 3398
rect 30012 3334 30064 3340
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 29736 3188 29788 3194
rect 29736 3130 29788 3136
rect 29552 2508 29604 2514
rect 29552 2450 29604 2456
rect 29368 2440 29420 2446
rect 29368 2382 29420 2388
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29380 2038 29408 2382
rect 29368 2032 29420 2038
rect 29368 1974 29420 1980
rect 28630 54 28856 82
rect 27802 0 27858 54
rect 28078 0 28134 54
rect 28354 0 28410 54
rect 28630 0 28686 54
rect 28906 0 28962 160
rect 29182 0 29238 160
rect 29458 82 29514 160
rect 29564 82 29592 2450
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29656 2106 29684 2246
rect 29644 2100 29696 2106
rect 29644 2042 29696 2048
rect 29748 160 29776 3130
rect 30024 3126 30052 3334
rect 30012 3120 30064 3126
rect 30012 3062 30064 3068
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 30104 2304 30156 2310
rect 30104 2246 30156 2252
rect 29458 54 29592 82
rect 29458 0 29514 54
rect 29734 0 29790 160
rect 30010 82 30066 160
rect 30116 82 30144 2246
rect 30010 54 30144 82
rect 30208 82 30236 2790
rect 30300 1970 30328 3334
rect 30392 3126 30420 5850
rect 30748 4276 30800 4282
rect 30748 4218 30800 4224
rect 30760 3618 30788 4218
rect 30852 3738 30880 7375
rect 31496 7274 31524 7822
rect 31772 7546 31800 9840
rect 32508 7546 32536 9840
rect 33244 7546 33272 9840
rect 33980 9738 34008 9840
rect 34072 9738 34100 9846
rect 33980 9710 34100 9738
rect 33790 7644 34098 7653
rect 33790 7642 33796 7644
rect 33852 7642 33876 7644
rect 33932 7642 33956 7644
rect 34012 7642 34036 7644
rect 34092 7642 34098 7644
rect 33852 7590 33854 7642
rect 34034 7590 34036 7642
rect 33790 7588 33796 7590
rect 33852 7588 33876 7590
rect 33932 7588 33956 7590
rect 34012 7588 34036 7590
rect 34092 7588 34098 7590
rect 33790 7579 34098 7588
rect 34256 7546 34284 9846
rect 34702 9840 34758 10000
rect 35438 9840 35494 10000
rect 35544 9846 35848 9874
rect 34716 7546 34744 9840
rect 35452 9738 35480 9840
rect 35544 9738 35572 9846
rect 35452 9710 35572 9738
rect 31760 7540 31812 7546
rect 31760 7482 31812 7488
rect 32496 7540 32548 7546
rect 32496 7482 32548 7488
rect 33232 7540 33284 7546
rect 33232 7482 33284 7488
rect 34244 7540 34296 7546
rect 34244 7482 34296 7488
rect 34704 7540 34756 7546
rect 35820 7528 35848 9846
rect 36174 9840 36230 10000
rect 36910 9840 36966 10000
rect 37016 9846 37228 9874
rect 36188 7546 36216 9840
rect 36924 9738 36952 9840
rect 37016 9738 37044 9846
rect 36924 9710 37044 9738
rect 36912 7812 36964 7818
rect 36912 7754 36964 7760
rect 36924 7546 36952 7754
rect 37200 7546 37228 9846
rect 37646 9840 37702 10000
rect 38382 9840 38438 10000
rect 39118 9840 39174 10000
rect 39854 9840 39910 10000
rect 40590 9840 40646 10000
rect 41326 9840 41382 10000
rect 42062 9840 42118 10000
rect 42168 9846 42656 9874
rect 37660 7546 37688 9840
rect 35900 7540 35952 7546
rect 35820 7500 35900 7528
rect 34704 7482 34756 7488
rect 35900 7482 35952 7488
rect 36176 7540 36228 7546
rect 36176 7482 36228 7488
rect 36912 7540 36964 7546
rect 36912 7482 36964 7488
rect 37188 7540 37240 7546
rect 37188 7482 37240 7488
rect 37648 7540 37700 7546
rect 38396 7528 38424 9840
rect 39132 7546 39160 9840
rect 39868 7546 39896 9840
rect 40604 7546 40632 9840
rect 41340 7546 41368 9840
rect 42076 9738 42104 9840
rect 42168 9738 42196 9846
rect 42076 9710 42196 9738
rect 42628 7546 42656 9846
rect 42798 9840 42854 10000
rect 43534 9840 43590 10000
rect 44270 9840 44326 10000
rect 45006 9840 45062 10000
rect 42708 7880 42760 7886
rect 42708 7822 42760 7828
rect 42720 7546 42748 7822
rect 42812 7546 42840 9840
rect 43548 7546 43576 9840
rect 38660 7540 38712 7546
rect 38396 7500 38660 7528
rect 37648 7482 37700 7488
rect 38660 7482 38712 7488
rect 39120 7540 39172 7546
rect 39120 7482 39172 7488
rect 39856 7540 39908 7546
rect 39856 7482 39908 7488
rect 40592 7540 40644 7546
rect 40592 7482 40644 7488
rect 41328 7540 41380 7546
rect 41328 7482 41380 7488
rect 42616 7540 42668 7546
rect 42616 7482 42668 7488
rect 42708 7540 42760 7546
rect 42708 7482 42760 7488
rect 42800 7540 42852 7546
rect 42800 7482 42852 7488
rect 43536 7540 43588 7546
rect 43536 7482 43588 7488
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 34152 7404 34204 7410
rect 34152 7346 34204 7352
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 35624 7404 35676 7410
rect 35624 7346 35676 7352
rect 35900 7404 35952 7410
rect 35900 7346 35952 7352
rect 37004 7404 37056 7410
rect 37004 7346 37056 7352
rect 37372 7404 37424 7410
rect 37372 7346 37424 7352
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 38936 7404 38988 7410
rect 38936 7346 38988 7352
rect 39396 7404 39448 7410
rect 39396 7346 39448 7352
rect 42616 7404 42668 7410
rect 42616 7346 42668 7352
rect 32784 7313 32812 7346
rect 32770 7304 32826 7313
rect 31484 7268 31536 7274
rect 32770 7239 32826 7248
rect 31484 7210 31536 7216
rect 31944 7200 31996 7206
rect 31944 7142 31996 7148
rect 33048 7200 33100 7206
rect 33048 7142 33100 7148
rect 31206 4176 31262 4185
rect 31206 4111 31262 4120
rect 31024 4072 31076 4078
rect 31024 4014 31076 4020
rect 30840 3732 30892 3738
rect 30840 3674 30892 3680
rect 30564 3596 30616 3602
rect 30760 3590 30880 3618
rect 30564 3538 30616 3544
rect 30576 3194 30604 3538
rect 30656 3460 30708 3466
rect 30656 3402 30708 3408
rect 30668 3369 30696 3402
rect 30654 3360 30710 3369
rect 30654 3295 30710 3304
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 30656 3120 30708 3126
rect 30656 3062 30708 3068
rect 30746 3088 30802 3097
rect 30564 2916 30616 2922
rect 30564 2858 30616 2864
rect 30380 2372 30432 2378
rect 30380 2314 30432 2320
rect 30392 2281 30420 2314
rect 30378 2272 30434 2281
rect 30378 2207 30434 2216
rect 30288 1964 30340 1970
rect 30288 1906 30340 1912
rect 30576 160 30604 2858
rect 30668 2281 30696 3062
rect 30746 3023 30748 3032
rect 30800 3023 30802 3032
rect 30748 2994 30800 3000
rect 30852 2774 30880 3590
rect 31036 3058 31064 4014
rect 31220 3534 31248 4111
rect 31208 3528 31260 3534
rect 31484 3528 31536 3534
rect 31208 3470 31260 3476
rect 31404 3488 31484 3516
rect 31300 3392 31352 3398
rect 31300 3334 31352 3340
rect 31312 3194 31340 3334
rect 31300 3188 31352 3194
rect 31300 3130 31352 3136
rect 31404 3126 31432 3488
rect 31484 3470 31536 3476
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 31392 3120 31444 3126
rect 31392 3062 31444 3068
rect 31024 3052 31076 3058
rect 31024 2994 31076 3000
rect 31668 2848 31720 2854
rect 30760 2746 30880 2774
rect 31588 2808 31668 2836
rect 30760 2446 30788 2746
rect 31116 2644 31168 2650
rect 31116 2586 31168 2592
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 30654 2272 30710 2281
rect 30654 2207 30710 2216
rect 30852 2038 30880 2382
rect 30840 2032 30892 2038
rect 30840 1974 30892 1980
rect 31128 490 31156 2586
rect 31392 2440 31444 2446
rect 31312 2400 31392 2428
rect 31206 2136 31262 2145
rect 31206 2071 31262 2080
rect 31220 1766 31248 2071
rect 31208 1760 31260 1766
rect 31208 1702 31260 1708
rect 31208 1624 31260 1630
rect 31208 1566 31260 1572
rect 31220 1426 31248 1566
rect 31208 1420 31260 1426
rect 31208 1362 31260 1368
rect 31036 462 31156 490
rect 30286 82 30342 160
rect 30208 54 30342 82
rect 30010 0 30066 54
rect 30286 0 30342 54
rect 30562 0 30618 160
rect 30838 82 30894 160
rect 31036 82 31064 462
rect 30838 54 31064 82
rect 31114 82 31170 160
rect 31312 82 31340 2400
rect 31392 2382 31444 2388
rect 31392 1692 31444 1698
rect 31392 1634 31444 1640
rect 31404 1154 31432 1634
rect 31392 1148 31444 1154
rect 31392 1090 31444 1096
rect 31114 54 31340 82
rect 31390 82 31446 160
rect 31588 82 31616 2808
rect 31772 2825 31800 3470
rect 31852 3392 31904 3398
rect 31852 3334 31904 3340
rect 31864 3194 31892 3334
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 31668 2790 31720 2796
rect 31758 2816 31814 2825
rect 31758 2751 31814 2760
rect 31668 2508 31720 2514
rect 31668 2450 31720 2456
rect 31680 160 31708 2450
rect 31956 2446 31984 7142
rect 33060 6118 33088 7142
rect 33140 6724 33192 6730
rect 33140 6666 33192 6672
rect 33152 6390 33180 6666
rect 33140 6384 33192 6390
rect 33140 6326 33192 6332
rect 33048 6112 33100 6118
rect 33048 6054 33100 6060
rect 33428 5166 33456 7346
rect 34164 7002 34192 7346
rect 34900 7002 34928 7346
rect 35636 7002 35664 7346
rect 34152 6996 34204 7002
rect 34152 6938 34204 6944
rect 34428 6996 34480 7002
rect 34428 6938 34480 6944
rect 34888 6996 34940 7002
rect 34888 6938 34940 6944
rect 35624 6996 35676 7002
rect 35624 6938 35676 6944
rect 33790 6556 34098 6565
rect 33790 6554 33796 6556
rect 33852 6554 33876 6556
rect 33932 6554 33956 6556
rect 34012 6554 34036 6556
rect 34092 6554 34098 6556
rect 33852 6502 33854 6554
rect 34034 6502 34036 6554
rect 33790 6500 33796 6502
rect 33852 6500 33876 6502
rect 33932 6500 33956 6502
rect 34012 6500 34036 6502
rect 34092 6500 34098 6502
rect 33790 6491 34098 6500
rect 33790 5468 34098 5477
rect 33790 5466 33796 5468
rect 33852 5466 33876 5468
rect 33932 5466 33956 5468
rect 34012 5466 34036 5468
rect 34092 5466 34098 5468
rect 33852 5414 33854 5466
rect 34034 5414 34036 5466
rect 33790 5412 33796 5414
rect 33852 5412 33876 5414
rect 33932 5412 33956 5414
rect 34012 5412 34036 5414
rect 34092 5412 34098 5414
rect 33790 5403 34098 5412
rect 33416 5160 33468 5166
rect 33416 5102 33468 5108
rect 33790 4380 34098 4389
rect 33790 4378 33796 4380
rect 33852 4378 33876 4380
rect 33932 4378 33956 4380
rect 34012 4378 34036 4380
rect 34092 4378 34098 4380
rect 33852 4326 33854 4378
rect 34034 4326 34036 4378
rect 33790 4324 33796 4326
rect 33852 4324 33876 4326
rect 33932 4324 33956 4326
rect 34012 4324 34036 4326
rect 34092 4324 34098 4326
rect 33790 4315 34098 4324
rect 32036 4208 32088 4214
rect 32036 4150 32088 4156
rect 32048 3534 32076 4150
rect 32680 4140 32732 4146
rect 32680 4082 32732 4088
rect 32036 3528 32088 3534
rect 32036 3470 32088 3476
rect 32312 3528 32364 3534
rect 32312 3470 32364 3476
rect 32588 3528 32640 3534
rect 32692 3505 32720 4082
rect 33416 3936 33468 3942
rect 33416 3878 33468 3884
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 33140 3732 33192 3738
rect 33140 3674 33192 3680
rect 32588 3470 32640 3476
rect 32678 3496 32734 3505
rect 32128 3392 32180 3398
rect 32128 3334 32180 3340
rect 32140 3058 32168 3334
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 32036 2916 32088 2922
rect 32036 2858 32088 2864
rect 31944 2440 31996 2446
rect 31944 2382 31996 2388
rect 32048 1306 32076 2858
rect 32220 2372 32272 2378
rect 32220 2314 32272 2320
rect 32128 1964 32180 1970
rect 32128 1906 32180 1912
rect 32140 1426 32168 1906
rect 32232 1601 32260 2314
rect 32324 1873 32352 3470
rect 32496 3460 32548 3466
rect 32496 3402 32548 3408
rect 32508 3126 32536 3402
rect 32496 3120 32548 3126
rect 32496 3062 32548 3068
rect 32496 2848 32548 2854
rect 32496 2790 32548 2796
rect 32310 1864 32366 1873
rect 32310 1799 32366 1808
rect 32218 1592 32274 1601
rect 32218 1527 32274 1536
rect 32128 1420 32180 1426
rect 32128 1362 32180 1368
rect 32404 1420 32456 1426
rect 32404 1362 32456 1368
rect 31956 1278 32076 1306
rect 31956 160 31984 1278
rect 31390 54 31616 82
rect 30838 0 30894 54
rect 31114 0 31170 54
rect 31390 0 31446 54
rect 31666 0 31722 160
rect 31942 0 31998 160
rect 32218 82 32274 160
rect 32416 82 32444 1362
rect 32508 160 32536 2790
rect 32600 1329 32628 3470
rect 32678 3431 32734 3440
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 32692 2446 32720 3062
rect 32680 2440 32732 2446
rect 32680 2382 32732 2388
rect 32586 1320 32642 1329
rect 32586 1255 32642 1264
rect 32784 160 32812 3674
rect 32956 3460 33008 3466
rect 32956 3402 33008 3408
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 32876 3194 32904 3334
rect 32864 3188 32916 3194
rect 32864 3130 32916 3136
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 32876 2446 32904 2994
rect 32968 2650 32996 3402
rect 33048 2916 33100 2922
rect 33048 2858 33100 2864
rect 32956 2644 33008 2650
rect 32956 2586 33008 2592
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 33060 160 33088 2858
rect 33152 2446 33180 3674
rect 33428 3058 33456 3878
rect 34334 3768 34390 3777
rect 34334 3703 34390 3712
rect 33790 3292 34098 3301
rect 33790 3290 33796 3292
rect 33852 3290 33876 3292
rect 33932 3290 33956 3292
rect 34012 3290 34036 3292
rect 34092 3290 34098 3292
rect 33852 3238 33854 3290
rect 34034 3238 34036 3290
rect 33790 3236 33796 3238
rect 33852 3236 33876 3238
rect 33932 3236 33956 3238
rect 34012 3236 34036 3238
rect 34092 3236 34098 3238
rect 33790 3227 34098 3236
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33416 3052 33468 3058
rect 33416 2994 33468 3000
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 33140 2440 33192 2446
rect 33140 2382 33192 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33152 1426 33180 2246
rect 33428 2145 33456 2382
rect 33414 2136 33470 2145
rect 33414 2071 33470 2080
rect 33140 1420 33192 1426
rect 33140 1362 33192 1368
rect 32218 54 32444 82
rect 32218 0 32274 54
rect 32494 0 32550 160
rect 32770 0 32826 160
rect 33046 0 33102 160
rect 33322 82 33378 160
rect 33520 82 33548 2586
rect 33612 160 33640 3130
rect 34348 3058 34376 3703
rect 34336 3052 34388 3058
rect 34336 2994 34388 3000
rect 34152 2848 34204 2854
rect 34152 2790 34204 2796
rect 33790 2204 34098 2213
rect 33790 2202 33796 2204
rect 33852 2202 33876 2204
rect 33932 2202 33956 2204
rect 34012 2202 34036 2204
rect 34092 2202 34098 2204
rect 33852 2150 33854 2202
rect 34034 2150 34036 2202
rect 33790 2148 33796 2150
rect 33852 2148 33876 2150
rect 33932 2148 33956 2150
rect 34012 2148 34036 2150
rect 34092 2148 34098 2150
rect 33790 2139 34098 2148
rect 34060 1420 34112 1426
rect 34060 1362 34112 1368
rect 33322 54 33548 82
rect 33322 0 33378 54
rect 33598 0 33654 160
rect 33874 82 33930 160
rect 34072 82 34100 1362
rect 34164 160 34192 2790
rect 34440 2582 34468 6938
rect 35348 6860 35400 6866
rect 35348 6802 35400 6808
rect 34612 6792 34664 6798
rect 34612 6734 34664 6740
rect 34624 6458 34652 6734
rect 35256 6724 35308 6730
rect 35360 6712 35388 6802
rect 35308 6684 35388 6712
rect 35256 6666 35308 6672
rect 34612 6452 34664 6458
rect 34612 6394 34664 6400
rect 35912 6254 35940 7346
rect 37016 6934 37044 7346
rect 37004 6928 37056 6934
rect 37004 6870 37056 6876
rect 37384 6798 37412 7346
rect 37476 7002 37504 7346
rect 38212 7002 38240 7346
rect 38948 7002 38976 7346
rect 39408 7290 39436 7346
rect 39224 7262 39436 7290
rect 39224 7206 39252 7262
rect 39212 7200 39264 7206
rect 39212 7142 39264 7148
rect 39264 7100 39572 7109
rect 39264 7098 39270 7100
rect 39326 7098 39350 7100
rect 39406 7098 39430 7100
rect 39486 7098 39510 7100
rect 39566 7098 39572 7100
rect 39326 7046 39328 7098
rect 39508 7046 39510 7098
rect 39264 7044 39270 7046
rect 39326 7044 39350 7046
rect 39406 7044 39430 7046
rect 39486 7044 39510 7046
rect 39566 7044 39572 7046
rect 39264 7035 39572 7044
rect 37464 6996 37516 7002
rect 37464 6938 37516 6944
rect 38200 6996 38252 7002
rect 38200 6938 38252 6944
rect 38936 6996 38988 7002
rect 38936 6938 38988 6944
rect 37372 6792 37424 6798
rect 37372 6734 37424 6740
rect 38844 6792 38896 6798
rect 38844 6734 38896 6740
rect 36728 6724 36780 6730
rect 36728 6666 36780 6672
rect 36268 6656 36320 6662
rect 36268 6598 36320 6604
rect 36280 6458 36308 6598
rect 36268 6452 36320 6458
rect 36268 6394 36320 6400
rect 36740 6390 36768 6666
rect 38856 6458 38884 6734
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 36728 6384 36780 6390
rect 36728 6326 36780 6332
rect 35900 6248 35952 6254
rect 35900 6190 35952 6196
rect 39264 6012 39572 6021
rect 39264 6010 39270 6012
rect 39326 6010 39350 6012
rect 39406 6010 39430 6012
rect 39486 6010 39510 6012
rect 39566 6010 39572 6012
rect 39326 5958 39328 6010
rect 39508 5958 39510 6010
rect 39264 5956 39270 5958
rect 39326 5956 39350 5958
rect 39406 5956 39430 5958
rect 39486 5956 39510 5958
rect 39566 5956 39572 5958
rect 39264 5947 39572 5956
rect 37464 5840 37516 5846
rect 37464 5782 37516 5788
rect 37094 3632 37150 3641
rect 35440 3596 35492 3602
rect 37094 3567 37150 3576
rect 35440 3538 35492 3544
rect 35452 3194 35480 3538
rect 36634 3496 36690 3505
rect 36634 3431 36690 3440
rect 35440 3188 35492 3194
rect 35440 3130 35492 3136
rect 35072 3052 35124 3058
rect 35072 2994 35124 3000
rect 34428 2576 34480 2582
rect 34428 2518 34480 2524
rect 34336 2372 34388 2378
rect 34336 2314 34388 2320
rect 34796 2372 34848 2378
rect 34796 2314 34848 2320
rect 33874 54 34100 82
rect 33874 0 33930 54
rect 34150 0 34206 160
rect 34348 82 34376 2314
rect 34808 2106 34836 2314
rect 34796 2100 34848 2106
rect 34796 2042 34848 2048
rect 34426 82 34482 160
rect 34348 54 34482 82
rect 34426 0 34482 54
rect 34702 0 34758 160
rect 34978 82 35034 160
rect 35084 82 35112 2994
rect 35898 2952 35954 2961
rect 35898 2887 35954 2896
rect 35912 2650 35940 2887
rect 36648 2650 36676 3431
rect 37108 2650 37136 3567
rect 37476 2650 37504 5782
rect 39028 5228 39080 5234
rect 39028 5170 39080 5176
rect 37830 3088 37886 3097
rect 37830 3023 37886 3032
rect 38936 3052 38988 3058
rect 37844 2650 37872 3023
rect 38936 2994 38988 3000
rect 35900 2644 35952 2650
rect 35900 2586 35952 2592
rect 36636 2644 36688 2650
rect 36636 2586 36688 2592
rect 37096 2644 37148 2650
rect 37096 2586 37148 2592
rect 37464 2644 37516 2650
rect 37464 2586 37516 2592
rect 37832 2644 37884 2650
rect 37832 2586 37884 2592
rect 37004 2576 37056 2582
rect 36924 2524 37004 2530
rect 38108 2576 38160 2582
rect 36924 2518 37056 2524
rect 38106 2544 38108 2553
rect 38844 2576 38896 2582
rect 38160 2544 38162 2553
rect 35256 2508 35308 2514
rect 36544 2508 36596 2514
rect 35256 2450 35308 2456
rect 36372 2468 36544 2496
rect 35268 160 35296 2450
rect 35348 2372 35400 2378
rect 35900 2372 35952 2378
rect 35348 2314 35400 2320
rect 35728 2332 35900 2360
rect 35360 2106 35388 2314
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35348 2100 35400 2106
rect 35348 2042 35400 2048
rect 35452 1426 35480 2246
rect 35440 1420 35492 1426
rect 35440 1362 35492 1368
rect 34978 54 35112 82
rect 34978 0 35034 54
rect 35254 0 35310 160
rect 35530 82 35586 160
rect 35728 82 35756 2332
rect 35900 2314 35952 2320
rect 36084 2304 36136 2310
rect 36084 2246 36136 2252
rect 35820 1426 35940 1442
rect 35820 1420 35952 1426
rect 35820 1414 35900 1420
rect 35820 160 35848 1414
rect 35900 1362 35952 1368
rect 36096 160 36124 2246
rect 36372 160 36400 2468
rect 36544 2450 36596 2456
rect 36924 2502 37044 2518
rect 37924 2508 37976 2514
rect 36820 2440 36872 2446
rect 36542 2408 36598 2417
rect 36820 2382 36872 2388
rect 36542 2343 36598 2352
rect 36556 2310 36584 2343
rect 36544 2304 36596 2310
rect 36544 2246 36596 2252
rect 36636 2304 36688 2310
rect 36636 2246 36688 2252
rect 36648 160 36676 2246
rect 36832 1426 36860 2382
rect 36820 1420 36872 1426
rect 36820 1362 36872 1368
rect 36924 160 36952 2502
rect 37844 2468 37924 2496
rect 37648 2372 37700 2378
rect 37200 2332 37648 2360
rect 37200 160 37228 2332
rect 37648 2314 37700 2320
rect 37740 2304 37792 2310
rect 37740 2246 37792 2252
rect 37752 1737 37780 2246
rect 37738 1728 37794 1737
rect 37738 1663 37794 1672
rect 37844 218 37872 2468
rect 38844 2518 38896 2524
rect 38476 2508 38528 2514
rect 38106 2479 38162 2488
rect 37924 2450 37976 2456
rect 38304 2468 38476 2496
rect 38200 2372 38252 2378
rect 37660 190 37872 218
rect 37936 2332 38200 2360
rect 35530 54 35756 82
rect 35530 0 35586 54
rect 35806 0 35862 160
rect 36082 0 36138 160
rect 36358 0 36414 160
rect 36634 0 36690 160
rect 36910 0 36966 160
rect 37186 0 37242 160
rect 37462 82 37518 160
rect 37660 82 37688 190
rect 37462 54 37688 82
rect 37738 82 37794 160
rect 37936 82 37964 2332
rect 38200 2314 38252 2320
rect 38304 218 38332 2468
rect 38476 2450 38528 2456
rect 38752 2372 38804 2378
rect 38488 2332 38752 2360
rect 38384 2304 38436 2310
rect 38384 2246 38436 2252
rect 38396 1222 38424 2246
rect 38384 1216 38436 1222
rect 38384 1158 38436 1164
rect 38212 190 38332 218
rect 37738 54 37964 82
rect 38014 82 38070 160
rect 38212 82 38240 190
rect 38014 54 38240 82
rect 38290 82 38346 160
rect 38488 82 38516 2332
rect 38752 2314 38804 2320
rect 38856 1442 38884 2518
rect 38580 1414 38884 1442
rect 38580 160 38608 1414
rect 38290 54 38516 82
rect 37462 0 37518 54
rect 37738 0 37794 54
rect 38014 0 38070 54
rect 38290 0 38346 54
rect 38566 0 38622 160
rect 38842 82 38898 160
rect 38948 82 38976 2994
rect 39040 2650 39068 5170
rect 42628 5137 42656 7346
rect 44284 7002 44312 9840
rect 45020 7834 45048 9840
rect 45020 7806 45140 7834
rect 44737 7644 45045 7653
rect 44737 7642 44743 7644
rect 44799 7642 44823 7644
rect 44879 7642 44903 7644
rect 44959 7642 44983 7644
rect 45039 7642 45045 7644
rect 44799 7590 44801 7642
rect 44981 7590 44983 7642
rect 44737 7588 44743 7590
rect 44799 7588 44823 7590
rect 44879 7588 44903 7590
rect 44959 7588 44983 7590
rect 45039 7588 45045 7590
rect 44737 7579 45045 7588
rect 44272 6996 44324 7002
rect 44272 6938 44324 6944
rect 45112 6866 45140 7806
rect 45100 6860 45152 6866
rect 45100 6802 45152 6808
rect 43628 6724 43680 6730
rect 43628 6666 43680 6672
rect 43640 5914 43668 6666
rect 44737 6556 45045 6565
rect 44737 6554 44743 6556
rect 44799 6554 44823 6556
rect 44879 6554 44903 6556
rect 44959 6554 44983 6556
rect 45039 6554 45045 6556
rect 44799 6502 44801 6554
rect 44981 6502 44983 6554
rect 44737 6500 44743 6502
rect 44799 6500 44823 6502
rect 44879 6500 44903 6502
rect 44959 6500 44983 6502
rect 45039 6500 45045 6502
rect 44737 6491 45045 6500
rect 43628 5908 43680 5914
rect 43628 5850 43680 5856
rect 44737 5468 45045 5477
rect 44737 5466 44743 5468
rect 44799 5466 44823 5468
rect 44879 5466 44903 5468
rect 44959 5466 44983 5468
rect 45039 5466 45045 5468
rect 44799 5414 44801 5466
rect 44981 5414 44983 5466
rect 44737 5412 44743 5414
rect 44799 5412 44823 5414
rect 44879 5412 44903 5414
rect 44959 5412 44983 5414
rect 45039 5412 45045 5414
rect 44737 5403 45045 5412
rect 42614 5128 42670 5137
rect 42614 5063 42670 5072
rect 39264 4924 39572 4933
rect 39264 4922 39270 4924
rect 39326 4922 39350 4924
rect 39406 4922 39430 4924
rect 39486 4922 39510 4924
rect 39566 4922 39572 4924
rect 39326 4870 39328 4922
rect 39508 4870 39510 4922
rect 39264 4868 39270 4870
rect 39326 4868 39350 4870
rect 39406 4868 39430 4870
rect 39486 4868 39510 4870
rect 39566 4868 39572 4870
rect 39264 4859 39572 4868
rect 39120 4820 39172 4826
rect 39120 4762 39172 4768
rect 39132 3194 39160 4762
rect 44737 4380 45045 4389
rect 44737 4378 44743 4380
rect 44799 4378 44823 4380
rect 44879 4378 44903 4380
rect 44959 4378 44983 4380
rect 45039 4378 45045 4380
rect 44799 4326 44801 4378
rect 44981 4326 44983 4378
rect 44737 4324 44743 4326
rect 44799 4324 44823 4326
rect 44879 4324 44903 4326
rect 44959 4324 44983 4326
rect 45039 4324 45045 4326
rect 44737 4315 45045 4324
rect 39264 3836 39572 3845
rect 39264 3834 39270 3836
rect 39326 3834 39350 3836
rect 39406 3834 39430 3836
rect 39486 3834 39510 3836
rect 39566 3834 39572 3836
rect 39326 3782 39328 3834
rect 39508 3782 39510 3834
rect 39264 3780 39270 3782
rect 39326 3780 39350 3782
rect 39406 3780 39430 3782
rect 39486 3780 39510 3782
rect 39566 3780 39572 3782
rect 39264 3771 39572 3780
rect 44737 3292 45045 3301
rect 44737 3290 44743 3292
rect 44799 3290 44823 3292
rect 44879 3290 44903 3292
rect 44959 3290 44983 3292
rect 45039 3290 45045 3292
rect 44799 3238 44801 3290
rect 44981 3238 44983 3290
rect 44737 3236 44743 3238
rect 44799 3236 44823 3238
rect 44879 3236 44903 3238
rect 44959 3236 44983 3238
rect 45039 3236 45045 3238
rect 44737 3227 45045 3236
rect 39120 3188 39172 3194
rect 39120 3130 39172 3136
rect 39264 2748 39572 2757
rect 39264 2746 39270 2748
rect 39326 2746 39350 2748
rect 39406 2746 39430 2748
rect 39486 2746 39510 2748
rect 39566 2746 39572 2748
rect 39326 2694 39328 2746
rect 39508 2694 39510 2746
rect 39264 2692 39270 2694
rect 39326 2692 39350 2694
rect 39406 2692 39430 2694
rect 39486 2692 39510 2694
rect 39566 2692 39572 2694
rect 39264 2683 39572 2692
rect 39028 2644 39080 2650
rect 39028 2586 39080 2592
rect 39396 2508 39448 2514
rect 40040 2508 40092 2514
rect 39396 2450 39448 2456
rect 39960 2468 40040 2496
rect 39120 2372 39172 2378
rect 39120 2314 39172 2320
rect 39028 2304 39080 2310
rect 39028 2246 39080 2252
rect 39040 2106 39068 2246
rect 39028 2100 39080 2106
rect 39028 2042 39080 2048
rect 39132 160 39160 2314
rect 39304 2304 39356 2310
rect 39304 2246 39356 2252
rect 39316 1970 39344 2246
rect 39304 1964 39356 1970
rect 39304 1906 39356 1912
rect 39408 160 39436 2450
rect 39672 2304 39724 2310
rect 39672 2246 39724 2252
rect 39684 1562 39712 2246
rect 39672 1556 39724 1562
rect 39672 1498 39724 1504
rect 39856 1420 39908 1426
rect 39856 1362 39908 1368
rect 38842 54 38976 82
rect 38842 0 38898 54
rect 39118 0 39174 160
rect 39394 0 39450 160
rect 39670 82 39726 160
rect 39868 82 39896 1362
rect 39960 160 39988 2468
rect 40040 2450 40092 2456
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 40224 2372 40276 2378
rect 40224 2314 40276 2320
rect 40040 2304 40092 2310
rect 40040 2246 40092 2252
rect 40052 2009 40080 2246
rect 40038 2000 40094 2009
rect 40038 1935 40094 1944
rect 40236 160 40264 2314
rect 40316 2304 40368 2310
rect 40316 2246 40368 2252
rect 40328 1562 40356 2246
rect 40316 1556 40368 1562
rect 40316 1498 40368 1504
rect 40420 1426 40448 2382
rect 40684 2304 40736 2310
rect 40684 2246 40736 2252
rect 40868 2304 40920 2310
rect 40868 2246 40920 2252
rect 41144 2304 41196 2310
rect 41144 2246 41196 2252
rect 40696 1766 40724 2246
rect 40684 1760 40736 1766
rect 40684 1702 40736 1708
rect 40408 1420 40460 1426
rect 40408 1362 40460 1368
rect 40880 1358 40908 2246
rect 40868 1352 40920 1358
rect 40868 1294 40920 1300
rect 41156 1290 41184 2246
rect 44737 2204 45045 2213
rect 44737 2202 44743 2204
rect 44799 2202 44823 2204
rect 44879 2202 44903 2204
rect 44959 2202 44983 2204
rect 45039 2202 45045 2204
rect 44799 2150 44801 2202
rect 44981 2150 44983 2202
rect 44737 2148 44743 2150
rect 44799 2148 44823 2150
rect 44879 2148 44903 2150
rect 44959 2148 44983 2150
rect 45039 2148 45045 2150
rect 44737 2139 45045 2148
rect 41144 1284 41196 1290
rect 41144 1226 41196 1232
rect 39670 54 39896 82
rect 39670 0 39726 54
rect 39946 0 40002 160
rect 40222 0 40278 160
<< via2 >>
rect 1766 7404 1822 7440
rect 1766 7384 1768 7404
rect 1768 7384 1820 7404
rect 1820 7384 1822 7404
rect 6429 7098 6485 7100
rect 6509 7098 6565 7100
rect 6589 7098 6645 7100
rect 6669 7098 6725 7100
rect 6429 7046 6475 7098
rect 6475 7046 6485 7098
rect 6509 7046 6539 7098
rect 6539 7046 6551 7098
rect 6551 7046 6565 7098
rect 6589 7046 6603 7098
rect 6603 7046 6615 7098
rect 6615 7046 6645 7098
rect 6669 7046 6679 7098
rect 6679 7046 6725 7098
rect 6429 7044 6485 7046
rect 6509 7044 6565 7046
rect 6589 7044 6645 7046
rect 6669 7044 6725 7046
rect 4618 6160 4674 6216
rect 6429 6010 6485 6012
rect 6509 6010 6565 6012
rect 6589 6010 6645 6012
rect 6669 6010 6725 6012
rect 6429 5958 6475 6010
rect 6475 5958 6485 6010
rect 6509 5958 6539 6010
rect 6539 5958 6551 6010
rect 6551 5958 6565 6010
rect 6589 5958 6603 6010
rect 6603 5958 6615 6010
rect 6615 5958 6645 6010
rect 6669 5958 6679 6010
rect 6679 5958 6725 6010
rect 6429 5956 6485 5958
rect 6509 5956 6565 5958
rect 6589 5956 6645 5958
rect 6669 5956 6725 5958
rect 6429 4922 6485 4924
rect 6509 4922 6565 4924
rect 6589 4922 6645 4924
rect 6669 4922 6725 4924
rect 6429 4870 6475 4922
rect 6475 4870 6485 4922
rect 6509 4870 6539 4922
rect 6539 4870 6551 4922
rect 6551 4870 6565 4922
rect 6589 4870 6603 4922
rect 6603 4870 6615 4922
rect 6615 4870 6645 4922
rect 6669 4870 6679 4922
rect 6679 4870 6725 4922
rect 6429 4868 6485 4870
rect 6509 4868 6565 4870
rect 6589 4868 6645 4870
rect 6669 4868 6725 4870
rect 11702 7792 11758 7848
rect 11902 7642 11958 7644
rect 11982 7642 12038 7644
rect 12062 7642 12118 7644
rect 12142 7642 12198 7644
rect 11902 7590 11948 7642
rect 11948 7590 11958 7642
rect 11982 7590 12012 7642
rect 12012 7590 12024 7642
rect 12024 7590 12038 7642
rect 12062 7590 12076 7642
rect 12076 7590 12088 7642
rect 12088 7590 12118 7642
rect 12142 7590 12152 7642
rect 12152 7590 12198 7642
rect 11902 7588 11958 7590
rect 11982 7588 12038 7590
rect 12062 7588 12118 7590
rect 12142 7588 12198 7590
rect 7930 4528 7986 4584
rect 6429 3834 6485 3836
rect 6509 3834 6565 3836
rect 6589 3834 6645 3836
rect 6669 3834 6725 3836
rect 6429 3782 6475 3834
rect 6475 3782 6485 3834
rect 6509 3782 6539 3834
rect 6539 3782 6551 3834
rect 6551 3782 6565 3834
rect 6589 3782 6603 3834
rect 6603 3782 6615 3834
rect 6615 3782 6645 3834
rect 6669 3782 6679 3834
rect 6679 3782 6725 3834
rect 6429 3780 6485 3782
rect 6509 3780 6565 3782
rect 6589 3780 6645 3782
rect 6669 3780 6725 3782
rect 6826 2760 6882 2816
rect 6429 2746 6485 2748
rect 6509 2746 6565 2748
rect 6589 2746 6645 2748
rect 6669 2746 6725 2748
rect 6429 2694 6475 2746
rect 6475 2694 6485 2746
rect 6509 2694 6539 2746
rect 6539 2694 6551 2746
rect 6551 2694 6565 2746
rect 6589 2694 6603 2746
rect 6603 2694 6615 2746
rect 6615 2694 6645 2746
rect 6669 2694 6679 2746
rect 6679 2694 6725 2746
rect 6429 2692 6485 2694
rect 6509 2692 6565 2694
rect 6589 2692 6645 2694
rect 6669 2692 6725 2694
rect 7102 992 7158 1048
rect 8482 3440 8538 3496
rect 8758 3032 8814 3088
rect 9402 2896 9458 2952
rect 9954 2488 10010 2544
rect 9586 2352 9642 2408
rect 10230 1672 10286 1728
rect 11902 6554 11958 6556
rect 11982 6554 12038 6556
rect 12062 6554 12118 6556
rect 12142 6554 12198 6556
rect 11902 6502 11948 6554
rect 11948 6502 11958 6554
rect 11982 6502 12012 6554
rect 12012 6502 12024 6554
rect 12024 6502 12038 6554
rect 12062 6502 12076 6554
rect 12076 6502 12088 6554
rect 12088 6502 12118 6554
rect 12142 6502 12152 6554
rect 12152 6502 12198 6554
rect 11902 6500 11958 6502
rect 11982 6500 12038 6502
rect 12062 6500 12118 6502
rect 12142 6500 12198 6502
rect 11902 5466 11958 5468
rect 11982 5466 12038 5468
rect 12062 5466 12118 5468
rect 12142 5466 12198 5468
rect 11902 5414 11948 5466
rect 11948 5414 11958 5466
rect 11982 5414 12012 5466
rect 12012 5414 12024 5466
rect 12024 5414 12038 5466
rect 12062 5414 12076 5466
rect 12076 5414 12088 5466
rect 12088 5414 12118 5466
rect 12142 5414 12152 5466
rect 12152 5414 12198 5466
rect 11902 5412 11958 5414
rect 11982 5412 12038 5414
rect 12062 5412 12118 5414
rect 12142 5412 12198 5414
rect 11902 4378 11958 4380
rect 11982 4378 12038 4380
rect 12062 4378 12118 4380
rect 12142 4378 12198 4380
rect 11902 4326 11948 4378
rect 11948 4326 11958 4378
rect 11982 4326 12012 4378
rect 12012 4326 12024 4378
rect 12024 4326 12038 4378
rect 12062 4326 12076 4378
rect 12076 4326 12088 4378
rect 12088 4326 12118 4378
rect 12142 4326 12152 4378
rect 12152 4326 12198 4378
rect 11902 4324 11958 4326
rect 11982 4324 12038 4326
rect 12062 4324 12118 4326
rect 12142 4324 12198 4326
rect 11334 3984 11390 4040
rect 11902 3290 11958 3292
rect 11982 3290 12038 3292
rect 12062 3290 12118 3292
rect 12142 3290 12198 3292
rect 11902 3238 11948 3290
rect 11948 3238 11958 3290
rect 11982 3238 12012 3290
rect 12012 3238 12024 3290
rect 12024 3238 12038 3290
rect 12062 3238 12076 3290
rect 12076 3238 12088 3290
rect 12088 3238 12118 3290
rect 12142 3238 12152 3290
rect 12152 3238 12198 3290
rect 11902 3236 11958 3238
rect 11982 3236 12038 3238
rect 12062 3236 12118 3238
rect 12142 3236 12198 3238
rect 13358 3576 13414 3632
rect 11902 2202 11958 2204
rect 11982 2202 12038 2204
rect 12062 2202 12118 2204
rect 12142 2202 12198 2204
rect 11902 2150 11948 2202
rect 11948 2150 11958 2202
rect 11982 2150 12012 2202
rect 12012 2150 12024 2202
rect 12024 2150 12038 2202
rect 12062 2150 12076 2202
rect 12076 2150 12088 2202
rect 12088 2150 12118 2202
rect 12142 2150 12152 2202
rect 12152 2150 12198 2202
rect 11902 2148 11958 2150
rect 11982 2148 12038 2150
rect 12062 2148 12118 2150
rect 12142 2148 12198 2150
rect 12990 2216 13046 2272
rect 13082 1808 13138 1864
rect 14554 4120 14610 4176
rect 14462 3168 14518 3224
rect 14186 1944 14242 2000
rect 14462 2760 14518 2816
rect 15566 3304 15622 3360
rect 15198 1128 15254 1184
rect 17376 7098 17432 7100
rect 17456 7098 17512 7100
rect 17536 7098 17592 7100
rect 17616 7098 17672 7100
rect 17376 7046 17422 7098
rect 17422 7046 17432 7098
rect 17456 7046 17486 7098
rect 17486 7046 17498 7098
rect 17498 7046 17512 7098
rect 17536 7046 17550 7098
rect 17550 7046 17562 7098
rect 17562 7046 17592 7098
rect 17616 7046 17626 7098
rect 17626 7046 17672 7098
rect 17376 7044 17432 7046
rect 17456 7044 17512 7046
rect 17536 7044 17592 7046
rect 17616 7044 17672 7046
rect 17376 6010 17432 6012
rect 17456 6010 17512 6012
rect 17536 6010 17592 6012
rect 17616 6010 17672 6012
rect 17376 5958 17422 6010
rect 17422 5958 17432 6010
rect 17456 5958 17486 6010
rect 17486 5958 17498 6010
rect 17498 5958 17512 6010
rect 17536 5958 17550 6010
rect 17550 5958 17562 6010
rect 17562 5958 17592 6010
rect 17616 5958 17626 6010
rect 17626 5958 17672 6010
rect 17376 5956 17432 5958
rect 17456 5956 17512 5958
rect 17536 5956 17592 5958
rect 17616 5956 17672 5958
rect 17376 4922 17432 4924
rect 17456 4922 17512 4924
rect 17536 4922 17592 4924
rect 17616 4922 17672 4924
rect 17376 4870 17422 4922
rect 17422 4870 17432 4922
rect 17456 4870 17486 4922
rect 17486 4870 17498 4922
rect 17498 4870 17512 4922
rect 17536 4870 17550 4922
rect 17550 4870 17562 4922
rect 17562 4870 17592 4922
rect 17616 4870 17626 4922
rect 17626 4870 17672 4922
rect 17376 4868 17432 4870
rect 17456 4868 17512 4870
rect 17536 4868 17592 4870
rect 17616 4868 17672 4870
rect 17376 3834 17432 3836
rect 17456 3834 17512 3836
rect 17536 3834 17592 3836
rect 17616 3834 17672 3836
rect 17376 3782 17422 3834
rect 17422 3782 17432 3834
rect 17456 3782 17486 3834
rect 17486 3782 17498 3834
rect 17498 3782 17512 3834
rect 17536 3782 17550 3834
rect 17550 3782 17562 3834
rect 17562 3782 17592 3834
rect 17616 3782 17626 3834
rect 17626 3782 17672 3834
rect 17376 3780 17432 3782
rect 17456 3780 17512 3782
rect 17536 3780 17592 3782
rect 17616 3780 17672 3782
rect 17866 7248 17922 7304
rect 18050 6296 18106 6352
rect 17376 2746 17432 2748
rect 17456 2746 17512 2748
rect 17536 2746 17592 2748
rect 17616 2746 17672 2748
rect 17376 2694 17422 2746
rect 17422 2694 17432 2746
rect 17456 2694 17486 2746
rect 17486 2694 17498 2746
rect 17498 2694 17512 2746
rect 17536 2694 17550 2746
rect 17550 2694 17562 2746
rect 17562 2694 17592 2746
rect 17616 2694 17626 2746
rect 17626 2694 17672 2746
rect 17376 2692 17432 2694
rect 17456 2692 17512 2694
rect 17536 2692 17592 2694
rect 17616 2692 17672 2694
rect 17958 2760 18014 2816
rect 18234 5072 18290 5128
rect 18970 4256 19026 4312
rect 19246 3848 19302 3904
rect 18326 2644 18382 2680
rect 18326 2624 18328 2644
rect 18328 2624 18380 2644
rect 18380 2624 18382 2644
rect 18510 2388 18512 2408
rect 18512 2388 18564 2408
rect 18564 2388 18566 2408
rect 18510 2352 18566 2388
rect 19154 2760 19210 2816
rect 19062 2624 19118 2680
rect 19338 2624 19394 2680
rect 19338 2216 19394 2272
rect 19154 1264 19210 1320
rect 18786 40 18842 96
rect 19062 40 19118 96
rect 20258 7928 20314 7984
rect 22849 7642 22905 7644
rect 22929 7642 22985 7644
rect 23009 7642 23065 7644
rect 23089 7642 23145 7644
rect 22849 7590 22895 7642
rect 22895 7590 22905 7642
rect 22929 7590 22959 7642
rect 22959 7590 22971 7642
rect 22971 7590 22985 7642
rect 23009 7590 23023 7642
rect 23023 7590 23035 7642
rect 23035 7590 23065 7642
rect 23089 7590 23099 7642
rect 23099 7590 23145 7642
rect 22849 7588 22905 7590
rect 22929 7588 22985 7590
rect 23009 7588 23065 7590
rect 23089 7588 23145 7590
rect 24950 7792 25006 7848
rect 19982 3168 20038 3224
rect 21546 2896 21602 2952
rect 21638 2488 21694 2544
rect 22006 3052 22062 3088
rect 22006 3032 22008 3052
rect 22008 3032 22060 3052
rect 22060 3032 22062 3052
rect 22849 6554 22905 6556
rect 22929 6554 22985 6556
rect 23009 6554 23065 6556
rect 23089 6554 23145 6556
rect 22849 6502 22895 6554
rect 22895 6502 22905 6554
rect 22929 6502 22959 6554
rect 22959 6502 22971 6554
rect 22971 6502 22985 6554
rect 23009 6502 23023 6554
rect 23023 6502 23035 6554
rect 23035 6502 23065 6554
rect 23089 6502 23099 6554
rect 23099 6502 23145 6554
rect 22849 6500 22905 6502
rect 22929 6500 22985 6502
rect 23009 6500 23065 6502
rect 23089 6500 23145 6502
rect 22849 5466 22905 5468
rect 22929 5466 22985 5468
rect 23009 5466 23065 5468
rect 23089 5466 23145 5468
rect 22849 5414 22895 5466
rect 22895 5414 22905 5466
rect 22929 5414 22959 5466
rect 22959 5414 22971 5466
rect 22971 5414 22985 5466
rect 23009 5414 23023 5466
rect 23023 5414 23035 5466
rect 23035 5414 23065 5466
rect 23089 5414 23099 5466
rect 23099 5414 23145 5466
rect 22849 5412 22905 5414
rect 22929 5412 22985 5414
rect 23009 5412 23065 5414
rect 23089 5412 23145 5414
rect 22190 3304 22246 3360
rect 22849 4378 22905 4380
rect 22929 4378 22985 4380
rect 23009 4378 23065 4380
rect 23089 4378 23145 4380
rect 22849 4326 22895 4378
rect 22895 4326 22905 4378
rect 22929 4326 22959 4378
rect 22959 4326 22971 4378
rect 22971 4326 22985 4378
rect 23009 4326 23023 4378
rect 23023 4326 23035 4378
rect 23035 4326 23065 4378
rect 23089 4326 23099 4378
rect 23099 4326 23145 4378
rect 22849 4324 22905 4326
rect 22929 4324 22985 4326
rect 23009 4324 23065 4326
rect 23089 4324 23145 4326
rect 23202 3476 23204 3496
rect 23204 3476 23256 3496
rect 23256 3476 23258 3496
rect 23202 3440 23258 3476
rect 22466 1672 22522 1728
rect 22849 3290 22905 3292
rect 22929 3290 22985 3292
rect 23009 3290 23065 3292
rect 23089 3290 23145 3292
rect 22849 3238 22895 3290
rect 22895 3238 22905 3290
rect 22929 3238 22959 3290
rect 22959 3238 22971 3290
rect 22971 3238 22985 3290
rect 23009 3238 23023 3290
rect 23023 3238 23035 3290
rect 23035 3238 23065 3290
rect 23089 3238 23099 3290
rect 23099 3238 23145 3290
rect 22849 3236 22905 3238
rect 22929 3236 22985 3238
rect 23009 3236 23065 3238
rect 23089 3236 23145 3238
rect 22650 1536 22706 1592
rect 22849 2202 22905 2204
rect 22929 2202 22985 2204
rect 23009 2202 23065 2204
rect 23089 2202 23145 2204
rect 22849 2150 22895 2202
rect 22895 2150 22905 2202
rect 22929 2150 22959 2202
rect 22959 2150 22971 2202
rect 22971 2150 22985 2202
rect 23009 2150 23023 2202
rect 23023 2150 23035 2202
rect 23035 2150 23065 2202
rect 23089 2150 23099 2202
rect 23099 2150 23145 2202
rect 22849 2148 22905 2150
rect 22929 2148 22985 2150
rect 23009 2148 23065 2150
rect 23089 2148 23145 2150
rect 24030 4528 24086 4584
rect 24030 3032 24086 3088
rect 25226 3476 25228 3496
rect 25228 3476 25280 3496
rect 25280 3476 25282 3496
rect 25226 3440 25282 3476
rect 24766 2352 24822 2408
rect 26790 6296 26846 6352
rect 25686 3304 25742 3360
rect 26514 2644 26570 2680
rect 26514 2624 26516 2644
rect 26516 2624 26568 2644
rect 26568 2624 26570 2644
rect 26698 2488 26754 2544
rect 27618 3576 27674 3632
rect 27526 3476 27528 3496
rect 27528 3476 27580 3496
rect 27580 3476 27582 3496
rect 27526 3440 27582 3476
rect 26790 1672 26846 1728
rect 28998 7928 29054 7984
rect 30838 7384 30894 7440
rect 28323 7098 28379 7100
rect 28403 7098 28459 7100
rect 28483 7098 28539 7100
rect 28563 7098 28619 7100
rect 28323 7046 28369 7098
rect 28369 7046 28379 7098
rect 28403 7046 28433 7098
rect 28433 7046 28445 7098
rect 28445 7046 28459 7098
rect 28483 7046 28497 7098
rect 28497 7046 28509 7098
rect 28509 7046 28539 7098
rect 28563 7046 28573 7098
rect 28573 7046 28619 7098
rect 28323 7044 28379 7046
rect 28403 7044 28459 7046
rect 28483 7044 28539 7046
rect 28563 7044 28619 7046
rect 28323 6010 28379 6012
rect 28403 6010 28459 6012
rect 28483 6010 28539 6012
rect 28563 6010 28619 6012
rect 28323 5958 28369 6010
rect 28369 5958 28379 6010
rect 28403 5958 28433 6010
rect 28433 5958 28445 6010
rect 28445 5958 28459 6010
rect 28483 5958 28497 6010
rect 28497 5958 28509 6010
rect 28509 5958 28539 6010
rect 28563 5958 28573 6010
rect 28573 5958 28619 6010
rect 28323 5956 28379 5958
rect 28403 5956 28459 5958
rect 28483 5956 28539 5958
rect 28563 5956 28619 5958
rect 28323 4922 28379 4924
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28323 4870 28369 4922
rect 28369 4870 28379 4922
rect 28403 4870 28433 4922
rect 28433 4870 28445 4922
rect 28445 4870 28459 4922
rect 28483 4870 28497 4922
rect 28497 4870 28509 4922
rect 28509 4870 28539 4922
rect 28563 4870 28573 4922
rect 28573 4870 28619 4922
rect 28323 4868 28379 4870
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 28323 3834 28379 3836
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28323 3782 28369 3834
rect 28369 3782 28379 3834
rect 28403 3782 28433 3834
rect 28433 3782 28445 3834
rect 28445 3782 28459 3834
rect 28483 3782 28497 3834
rect 28497 3782 28509 3834
rect 28509 3782 28539 3834
rect 28563 3782 28573 3834
rect 28573 3782 28619 3834
rect 28323 3780 28379 3782
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28722 3732 28778 3768
rect 28722 3712 28724 3732
rect 28724 3712 28776 3732
rect 28776 3712 28778 3732
rect 27986 2896 28042 2952
rect 27618 2352 27674 2408
rect 28323 2746 28379 2748
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28323 2694 28369 2746
rect 28369 2694 28379 2746
rect 28403 2694 28433 2746
rect 28433 2694 28445 2746
rect 28445 2694 28459 2746
rect 28483 2694 28497 2746
rect 28497 2694 28509 2746
rect 28509 2694 28539 2746
rect 28563 2694 28573 2746
rect 28573 2694 28619 2746
rect 28323 2692 28379 2694
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 28998 2760 29054 2816
rect 28998 1980 29000 2000
rect 29000 1980 29052 2000
rect 29052 1980 29054 2000
rect 28998 1944 29054 1980
rect 29826 6160 29882 6216
rect 30286 3984 30342 4040
rect 33796 7642 33852 7644
rect 33876 7642 33932 7644
rect 33956 7642 34012 7644
rect 34036 7642 34092 7644
rect 33796 7590 33842 7642
rect 33842 7590 33852 7642
rect 33876 7590 33906 7642
rect 33906 7590 33918 7642
rect 33918 7590 33932 7642
rect 33956 7590 33970 7642
rect 33970 7590 33982 7642
rect 33982 7590 34012 7642
rect 34036 7590 34046 7642
rect 34046 7590 34092 7642
rect 33796 7588 33852 7590
rect 33876 7588 33932 7590
rect 33956 7588 34012 7590
rect 34036 7588 34092 7590
rect 32770 7248 32826 7304
rect 31206 4120 31262 4176
rect 30654 3304 30710 3360
rect 30378 2216 30434 2272
rect 30746 3052 30802 3088
rect 30746 3032 30748 3052
rect 30748 3032 30800 3052
rect 30800 3032 30802 3052
rect 30654 2216 30710 2272
rect 31206 2080 31262 2136
rect 31758 2760 31814 2816
rect 33796 6554 33852 6556
rect 33876 6554 33932 6556
rect 33956 6554 34012 6556
rect 34036 6554 34092 6556
rect 33796 6502 33842 6554
rect 33842 6502 33852 6554
rect 33876 6502 33906 6554
rect 33906 6502 33918 6554
rect 33918 6502 33932 6554
rect 33956 6502 33970 6554
rect 33970 6502 33982 6554
rect 33982 6502 34012 6554
rect 34036 6502 34046 6554
rect 34046 6502 34092 6554
rect 33796 6500 33852 6502
rect 33876 6500 33932 6502
rect 33956 6500 34012 6502
rect 34036 6500 34092 6502
rect 33796 5466 33852 5468
rect 33876 5466 33932 5468
rect 33956 5466 34012 5468
rect 34036 5466 34092 5468
rect 33796 5414 33842 5466
rect 33842 5414 33852 5466
rect 33876 5414 33906 5466
rect 33906 5414 33918 5466
rect 33918 5414 33932 5466
rect 33956 5414 33970 5466
rect 33970 5414 33982 5466
rect 33982 5414 34012 5466
rect 34036 5414 34046 5466
rect 34046 5414 34092 5466
rect 33796 5412 33852 5414
rect 33876 5412 33932 5414
rect 33956 5412 34012 5414
rect 34036 5412 34092 5414
rect 33796 4378 33852 4380
rect 33876 4378 33932 4380
rect 33956 4378 34012 4380
rect 34036 4378 34092 4380
rect 33796 4326 33842 4378
rect 33842 4326 33852 4378
rect 33876 4326 33906 4378
rect 33906 4326 33918 4378
rect 33918 4326 33932 4378
rect 33956 4326 33970 4378
rect 33970 4326 33982 4378
rect 33982 4326 34012 4378
rect 34036 4326 34046 4378
rect 34046 4326 34092 4378
rect 33796 4324 33852 4326
rect 33876 4324 33932 4326
rect 33956 4324 34012 4326
rect 34036 4324 34092 4326
rect 32310 1808 32366 1864
rect 32218 1536 32274 1592
rect 32678 3440 32734 3496
rect 32586 1264 32642 1320
rect 34334 3712 34390 3768
rect 33796 3290 33852 3292
rect 33876 3290 33932 3292
rect 33956 3290 34012 3292
rect 34036 3290 34092 3292
rect 33796 3238 33842 3290
rect 33842 3238 33852 3290
rect 33876 3238 33906 3290
rect 33906 3238 33918 3290
rect 33918 3238 33932 3290
rect 33956 3238 33970 3290
rect 33970 3238 33982 3290
rect 33982 3238 34012 3290
rect 34036 3238 34046 3290
rect 34046 3238 34092 3290
rect 33796 3236 33852 3238
rect 33876 3236 33932 3238
rect 33956 3236 34012 3238
rect 34036 3236 34092 3238
rect 33414 2080 33470 2136
rect 33796 2202 33852 2204
rect 33876 2202 33932 2204
rect 33956 2202 34012 2204
rect 34036 2202 34092 2204
rect 33796 2150 33842 2202
rect 33842 2150 33852 2202
rect 33876 2150 33906 2202
rect 33906 2150 33918 2202
rect 33918 2150 33932 2202
rect 33956 2150 33970 2202
rect 33970 2150 33982 2202
rect 33982 2150 34012 2202
rect 34036 2150 34046 2202
rect 34046 2150 34092 2202
rect 33796 2148 33852 2150
rect 33876 2148 33932 2150
rect 33956 2148 34012 2150
rect 34036 2148 34092 2150
rect 39270 7098 39326 7100
rect 39350 7098 39406 7100
rect 39430 7098 39486 7100
rect 39510 7098 39566 7100
rect 39270 7046 39316 7098
rect 39316 7046 39326 7098
rect 39350 7046 39380 7098
rect 39380 7046 39392 7098
rect 39392 7046 39406 7098
rect 39430 7046 39444 7098
rect 39444 7046 39456 7098
rect 39456 7046 39486 7098
rect 39510 7046 39520 7098
rect 39520 7046 39566 7098
rect 39270 7044 39326 7046
rect 39350 7044 39406 7046
rect 39430 7044 39486 7046
rect 39510 7044 39566 7046
rect 39270 6010 39326 6012
rect 39350 6010 39406 6012
rect 39430 6010 39486 6012
rect 39510 6010 39566 6012
rect 39270 5958 39316 6010
rect 39316 5958 39326 6010
rect 39350 5958 39380 6010
rect 39380 5958 39392 6010
rect 39392 5958 39406 6010
rect 39430 5958 39444 6010
rect 39444 5958 39456 6010
rect 39456 5958 39486 6010
rect 39510 5958 39520 6010
rect 39520 5958 39566 6010
rect 39270 5956 39326 5958
rect 39350 5956 39406 5958
rect 39430 5956 39486 5958
rect 39510 5956 39566 5958
rect 37094 3576 37150 3632
rect 36634 3440 36690 3496
rect 35898 2896 35954 2952
rect 37830 3032 37886 3088
rect 38106 2524 38108 2544
rect 38108 2524 38160 2544
rect 38160 2524 38162 2544
rect 36542 2352 36598 2408
rect 37738 1672 37794 1728
rect 38106 2488 38162 2524
rect 44743 7642 44799 7644
rect 44823 7642 44879 7644
rect 44903 7642 44959 7644
rect 44983 7642 45039 7644
rect 44743 7590 44789 7642
rect 44789 7590 44799 7642
rect 44823 7590 44853 7642
rect 44853 7590 44865 7642
rect 44865 7590 44879 7642
rect 44903 7590 44917 7642
rect 44917 7590 44929 7642
rect 44929 7590 44959 7642
rect 44983 7590 44993 7642
rect 44993 7590 45039 7642
rect 44743 7588 44799 7590
rect 44823 7588 44879 7590
rect 44903 7588 44959 7590
rect 44983 7588 45039 7590
rect 44743 6554 44799 6556
rect 44823 6554 44879 6556
rect 44903 6554 44959 6556
rect 44983 6554 45039 6556
rect 44743 6502 44789 6554
rect 44789 6502 44799 6554
rect 44823 6502 44853 6554
rect 44853 6502 44865 6554
rect 44865 6502 44879 6554
rect 44903 6502 44917 6554
rect 44917 6502 44929 6554
rect 44929 6502 44959 6554
rect 44983 6502 44993 6554
rect 44993 6502 45039 6554
rect 44743 6500 44799 6502
rect 44823 6500 44879 6502
rect 44903 6500 44959 6502
rect 44983 6500 45039 6502
rect 44743 5466 44799 5468
rect 44823 5466 44879 5468
rect 44903 5466 44959 5468
rect 44983 5466 45039 5468
rect 44743 5414 44789 5466
rect 44789 5414 44799 5466
rect 44823 5414 44853 5466
rect 44853 5414 44865 5466
rect 44865 5414 44879 5466
rect 44903 5414 44917 5466
rect 44917 5414 44929 5466
rect 44929 5414 44959 5466
rect 44983 5414 44993 5466
rect 44993 5414 45039 5466
rect 44743 5412 44799 5414
rect 44823 5412 44879 5414
rect 44903 5412 44959 5414
rect 44983 5412 45039 5414
rect 42614 5072 42670 5128
rect 39270 4922 39326 4924
rect 39350 4922 39406 4924
rect 39430 4922 39486 4924
rect 39510 4922 39566 4924
rect 39270 4870 39316 4922
rect 39316 4870 39326 4922
rect 39350 4870 39380 4922
rect 39380 4870 39392 4922
rect 39392 4870 39406 4922
rect 39430 4870 39444 4922
rect 39444 4870 39456 4922
rect 39456 4870 39486 4922
rect 39510 4870 39520 4922
rect 39520 4870 39566 4922
rect 39270 4868 39326 4870
rect 39350 4868 39406 4870
rect 39430 4868 39486 4870
rect 39510 4868 39566 4870
rect 44743 4378 44799 4380
rect 44823 4378 44879 4380
rect 44903 4378 44959 4380
rect 44983 4378 45039 4380
rect 44743 4326 44789 4378
rect 44789 4326 44799 4378
rect 44823 4326 44853 4378
rect 44853 4326 44865 4378
rect 44865 4326 44879 4378
rect 44903 4326 44917 4378
rect 44917 4326 44929 4378
rect 44929 4326 44959 4378
rect 44983 4326 44993 4378
rect 44993 4326 45039 4378
rect 44743 4324 44799 4326
rect 44823 4324 44879 4326
rect 44903 4324 44959 4326
rect 44983 4324 45039 4326
rect 39270 3834 39326 3836
rect 39350 3834 39406 3836
rect 39430 3834 39486 3836
rect 39510 3834 39566 3836
rect 39270 3782 39316 3834
rect 39316 3782 39326 3834
rect 39350 3782 39380 3834
rect 39380 3782 39392 3834
rect 39392 3782 39406 3834
rect 39430 3782 39444 3834
rect 39444 3782 39456 3834
rect 39456 3782 39486 3834
rect 39510 3782 39520 3834
rect 39520 3782 39566 3834
rect 39270 3780 39326 3782
rect 39350 3780 39406 3782
rect 39430 3780 39486 3782
rect 39510 3780 39566 3782
rect 44743 3290 44799 3292
rect 44823 3290 44879 3292
rect 44903 3290 44959 3292
rect 44983 3290 45039 3292
rect 44743 3238 44789 3290
rect 44789 3238 44799 3290
rect 44823 3238 44853 3290
rect 44853 3238 44865 3290
rect 44865 3238 44879 3290
rect 44903 3238 44917 3290
rect 44917 3238 44929 3290
rect 44929 3238 44959 3290
rect 44983 3238 44993 3290
rect 44993 3238 45039 3290
rect 44743 3236 44799 3238
rect 44823 3236 44879 3238
rect 44903 3236 44959 3238
rect 44983 3236 45039 3238
rect 39270 2746 39326 2748
rect 39350 2746 39406 2748
rect 39430 2746 39486 2748
rect 39510 2746 39566 2748
rect 39270 2694 39316 2746
rect 39316 2694 39326 2746
rect 39350 2694 39380 2746
rect 39380 2694 39392 2746
rect 39392 2694 39406 2746
rect 39430 2694 39444 2746
rect 39444 2694 39456 2746
rect 39456 2694 39486 2746
rect 39510 2694 39520 2746
rect 39520 2694 39566 2746
rect 39270 2692 39326 2694
rect 39350 2692 39406 2694
rect 39430 2692 39486 2694
rect 39510 2692 39566 2694
rect 40038 1944 40094 2000
rect 44743 2202 44799 2204
rect 44823 2202 44879 2204
rect 44903 2202 44959 2204
rect 44983 2202 45039 2204
rect 44743 2150 44789 2202
rect 44789 2150 44799 2202
rect 44823 2150 44853 2202
rect 44853 2150 44865 2202
rect 44865 2150 44879 2202
rect 44903 2150 44917 2202
rect 44917 2150 44929 2202
rect 44929 2150 44959 2202
rect 44983 2150 44993 2202
rect 44993 2150 45039 2202
rect 44743 2148 44799 2150
rect 44823 2148 44879 2150
rect 44903 2148 44959 2150
rect 44983 2148 45039 2150
<< metal3 >>
rect 20253 7986 20319 7989
rect 28993 7986 29059 7989
rect 20253 7984 29059 7986
rect 20253 7928 20258 7984
rect 20314 7928 28998 7984
rect 29054 7928 29059 7984
rect 20253 7926 29059 7928
rect 20253 7923 20319 7926
rect 28993 7923 29059 7926
rect 11697 7850 11763 7853
rect 24945 7850 25011 7853
rect 11697 7848 25011 7850
rect 11697 7792 11702 7848
rect 11758 7792 24950 7848
rect 25006 7792 25011 7848
rect 11697 7790 25011 7792
rect 11697 7787 11763 7790
rect 24945 7787 25011 7790
rect 11892 7648 12208 7649
rect 11892 7584 11898 7648
rect 11962 7584 11978 7648
rect 12042 7584 12058 7648
rect 12122 7584 12138 7648
rect 12202 7584 12208 7648
rect 11892 7583 12208 7584
rect 22839 7648 23155 7649
rect 22839 7584 22845 7648
rect 22909 7584 22925 7648
rect 22989 7584 23005 7648
rect 23069 7584 23085 7648
rect 23149 7584 23155 7648
rect 22839 7583 23155 7584
rect 33786 7648 34102 7649
rect 33786 7584 33792 7648
rect 33856 7584 33872 7648
rect 33936 7584 33952 7648
rect 34016 7584 34032 7648
rect 34096 7584 34102 7648
rect 33786 7583 34102 7584
rect 44733 7648 45049 7649
rect 44733 7584 44739 7648
rect 44803 7584 44819 7648
rect 44883 7584 44899 7648
rect 44963 7584 44979 7648
rect 45043 7584 45049 7648
rect 44733 7583 45049 7584
rect 1761 7442 1827 7445
rect 30833 7442 30899 7445
rect 1761 7440 30899 7442
rect 1761 7384 1766 7440
rect 1822 7384 30838 7440
rect 30894 7384 30899 7440
rect 1761 7382 30899 7384
rect 1761 7379 1827 7382
rect 30833 7379 30899 7382
rect 17861 7306 17927 7309
rect 32765 7306 32831 7309
rect 17861 7304 32831 7306
rect 17861 7248 17866 7304
rect 17922 7248 32770 7304
rect 32826 7248 32831 7304
rect 17861 7246 32831 7248
rect 17861 7243 17927 7246
rect 32765 7243 32831 7246
rect 6419 7104 6735 7105
rect 6419 7040 6425 7104
rect 6489 7040 6505 7104
rect 6569 7040 6585 7104
rect 6649 7040 6665 7104
rect 6729 7040 6735 7104
rect 6419 7039 6735 7040
rect 17366 7104 17682 7105
rect 17366 7040 17372 7104
rect 17436 7040 17452 7104
rect 17516 7040 17532 7104
rect 17596 7040 17612 7104
rect 17676 7040 17682 7104
rect 17366 7039 17682 7040
rect 28313 7104 28629 7105
rect 28313 7040 28319 7104
rect 28383 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28629 7104
rect 28313 7039 28629 7040
rect 39260 7104 39576 7105
rect 39260 7040 39266 7104
rect 39330 7040 39346 7104
rect 39410 7040 39426 7104
rect 39490 7040 39506 7104
rect 39570 7040 39576 7104
rect 39260 7039 39576 7040
rect 11892 6560 12208 6561
rect 11892 6496 11898 6560
rect 11962 6496 11978 6560
rect 12042 6496 12058 6560
rect 12122 6496 12138 6560
rect 12202 6496 12208 6560
rect 11892 6495 12208 6496
rect 22839 6560 23155 6561
rect 22839 6496 22845 6560
rect 22909 6496 22925 6560
rect 22989 6496 23005 6560
rect 23069 6496 23085 6560
rect 23149 6496 23155 6560
rect 22839 6495 23155 6496
rect 33786 6560 34102 6561
rect 33786 6496 33792 6560
rect 33856 6496 33872 6560
rect 33936 6496 33952 6560
rect 34016 6496 34032 6560
rect 34096 6496 34102 6560
rect 33786 6495 34102 6496
rect 44733 6560 45049 6561
rect 44733 6496 44739 6560
rect 44803 6496 44819 6560
rect 44883 6496 44899 6560
rect 44963 6496 44979 6560
rect 45043 6496 45049 6560
rect 44733 6495 45049 6496
rect 18045 6354 18111 6357
rect 26785 6354 26851 6357
rect 18045 6352 26851 6354
rect 18045 6296 18050 6352
rect 18106 6296 26790 6352
rect 26846 6296 26851 6352
rect 18045 6294 26851 6296
rect 18045 6291 18111 6294
rect 26785 6291 26851 6294
rect 4613 6218 4679 6221
rect 29821 6218 29887 6221
rect 4613 6216 29887 6218
rect 4613 6160 4618 6216
rect 4674 6160 29826 6216
rect 29882 6160 29887 6216
rect 4613 6158 29887 6160
rect 4613 6155 4679 6158
rect 29821 6155 29887 6158
rect 6419 6016 6735 6017
rect 6419 5952 6425 6016
rect 6489 5952 6505 6016
rect 6569 5952 6585 6016
rect 6649 5952 6665 6016
rect 6729 5952 6735 6016
rect 6419 5951 6735 5952
rect 17366 6016 17682 6017
rect 17366 5952 17372 6016
rect 17436 5952 17452 6016
rect 17516 5952 17532 6016
rect 17596 5952 17612 6016
rect 17676 5952 17682 6016
rect 17366 5951 17682 5952
rect 28313 6016 28629 6017
rect 28313 5952 28319 6016
rect 28383 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28629 6016
rect 28313 5951 28629 5952
rect 39260 6016 39576 6017
rect 39260 5952 39266 6016
rect 39330 5952 39346 6016
rect 39410 5952 39426 6016
rect 39490 5952 39506 6016
rect 39570 5952 39576 6016
rect 39260 5951 39576 5952
rect 11892 5472 12208 5473
rect 11892 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12208 5472
rect 11892 5407 12208 5408
rect 22839 5472 23155 5473
rect 22839 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23155 5472
rect 22839 5407 23155 5408
rect 33786 5472 34102 5473
rect 33786 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34102 5472
rect 33786 5407 34102 5408
rect 44733 5472 45049 5473
rect 44733 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45049 5472
rect 44733 5407 45049 5408
rect 18229 5130 18295 5133
rect 42609 5130 42675 5133
rect 18229 5128 42675 5130
rect 18229 5072 18234 5128
rect 18290 5072 42614 5128
rect 42670 5072 42675 5128
rect 18229 5070 42675 5072
rect 18229 5067 18295 5070
rect 42609 5067 42675 5070
rect 6419 4928 6735 4929
rect 6419 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6735 4928
rect 6419 4863 6735 4864
rect 17366 4928 17682 4929
rect 17366 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17682 4928
rect 17366 4863 17682 4864
rect 28313 4928 28629 4929
rect 28313 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28629 4928
rect 28313 4863 28629 4864
rect 39260 4928 39576 4929
rect 39260 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39576 4928
rect 39260 4863 39576 4864
rect 7925 4586 7991 4589
rect 24025 4586 24091 4589
rect 7925 4584 24091 4586
rect 7925 4528 7930 4584
rect 7986 4528 24030 4584
rect 24086 4528 24091 4584
rect 7925 4526 24091 4528
rect 7925 4523 7991 4526
rect 24025 4523 24091 4526
rect 11892 4384 12208 4385
rect 11892 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12208 4384
rect 11892 4319 12208 4320
rect 22839 4384 23155 4385
rect 22839 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23155 4384
rect 22839 4319 23155 4320
rect 33786 4384 34102 4385
rect 33786 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34102 4384
rect 33786 4319 34102 4320
rect 44733 4384 45049 4385
rect 44733 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45049 4384
rect 44733 4319 45049 4320
rect 18822 4252 18828 4316
rect 18892 4314 18898 4316
rect 18965 4314 19031 4317
rect 18892 4312 19031 4314
rect 18892 4256 18970 4312
rect 19026 4256 19031 4312
rect 18892 4254 19031 4256
rect 18892 4252 18898 4254
rect 18965 4251 19031 4254
rect 14549 4178 14615 4181
rect 31201 4178 31267 4181
rect 14549 4176 31267 4178
rect 14549 4120 14554 4176
rect 14610 4120 31206 4176
rect 31262 4120 31267 4176
rect 14549 4118 31267 4120
rect 14549 4115 14615 4118
rect 31201 4115 31267 4118
rect 11329 4042 11395 4045
rect 30281 4042 30347 4045
rect 11329 4040 30347 4042
rect 11329 3984 11334 4040
rect 11390 3984 30286 4040
rect 30342 3984 30347 4040
rect 11329 3982 30347 3984
rect 11329 3979 11395 3982
rect 30281 3979 30347 3982
rect 19241 3908 19307 3909
rect 19241 3906 19288 3908
rect 19196 3904 19288 3906
rect 19196 3848 19246 3904
rect 19196 3846 19288 3848
rect 19241 3844 19288 3846
rect 19352 3844 19358 3908
rect 19241 3843 19307 3844
rect 6419 3840 6735 3841
rect 6419 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6735 3840
rect 6419 3775 6735 3776
rect 17366 3840 17682 3841
rect 17366 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17682 3840
rect 17366 3775 17682 3776
rect 28313 3840 28629 3841
rect 28313 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28629 3840
rect 28313 3775 28629 3776
rect 39260 3840 39576 3841
rect 39260 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39576 3840
rect 39260 3775 39576 3776
rect 28717 3770 28783 3773
rect 34329 3770 34395 3773
rect 28717 3768 34395 3770
rect 28717 3712 28722 3768
rect 28778 3712 34334 3768
rect 34390 3712 34395 3768
rect 28717 3710 34395 3712
rect 28717 3707 28783 3710
rect 34329 3707 34395 3710
rect 13353 3634 13419 3637
rect 27613 3634 27679 3637
rect 37089 3634 37155 3637
rect 13353 3632 27679 3634
rect 13353 3576 13358 3632
rect 13414 3576 27618 3632
rect 27674 3576 27679 3632
rect 13353 3574 27679 3576
rect 13353 3571 13419 3574
rect 27613 3571 27679 3574
rect 31710 3632 37155 3634
rect 31710 3576 37094 3632
rect 37150 3576 37155 3632
rect 31710 3574 37155 3576
rect 8477 3498 8543 3501
rect 23197 3498 23263 3501
rect 8477 3496 23263 3498
rect 8477 3440 8482 3496
rect 8538 3440 23202 3496
rect 23258 3440 23263 3496
rect 8477 3438 23263 3440
rect 8477 3435 8543 3438
rect 23197 3435 23263 3438
rect 24894 3436 24900 3500
rect 24964 3498 24970 3500
rect 25221 3498 25287 3501
rect 24964 3496 25287 3498
rect 24964 3440 25226 3496
rect 25282 3440 25287 3496
rect 24964 3438 25287 3440
rect 24964 3436 24970 3438
rect 25221 3435 25287 3438
rect 27521 3498 27587 3501
rect 31710 3498 31770 3574
rect 37089 3571 37155 3574
rect 27521 3496 31770 3498
rect 27521 3440 27526 3496
rect 27582 3440 31770 3496
rect 27521 3438 31770 3440
rect 27521 3435 27587 3438
rect 31886 3436 31892 3500
rect 31956 3498 31962 3500
rect 32673 3498 32739 3501
rect 36629 3498 36695 3501
rect 31956 3496 32739 3498
rect 31956 3440 32678 3496
rect 32734 3440 32739 3496
rect 31956 3438 32739 3440
rect 31956 3436 31962 3438
rect 32673 3435 32739 3438
rect 32814 3496 36695 3498
rect 32814 3440 36634 3496
rect 36690 3440 36695 3496
rect 32814 3438 36695 3440
rect 15561 3362 15627 3365
rect 22185 3362 22251 3365
rect 15561 3360 22251 3362
rect 15561 3304 15566 3360
rect 15622 3304 22190 3360
rect 22246 3304 22251 3360
rect 15561 3302 22251 3304
rect 15561 3299 15627 3302
rect 22185 3299 22251 3302
rect 25681 3362 25747 3365
rect 30649 3362 30715 3365
rect 32814 3362 32874 3438
rect 36629 3435 36695 3438
rect 25681 3360 29378 3362
rect 25681 3304 25686 3360
rect 25742 3304 29378 3360
rect 25681 3302 29378 3304
rect 25681 3299 25747 3302
rect 11892 3296 12208 3297
rect 11892 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12208 3296
rect 11892 3231 12208 3232
rect 22839 3296 23155 3297
rect 22839 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23155 3296
rect 22839 3231 23155 3232
rect 14457 3226 14523 3229
rect 19977 3226 20043 3229
rect 14457 3224 20043 3226
rect 14457 3168 14462 3224
rect 14518 3168 19982 3224
rect 20038 3168 20043 3224
rect 14457 3166 20043 3168
rect 29318 3226 29378 3302
rect 30649 3360 32874 3362
rect 30649 3304 30654 3360
rect 30710 3304 32874 3360
rect 30649 3302 32874 3304
rect 30649 3299 30715 3302
rect 33786 3296 34102 3297
rect 33786 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34102 3296
rect 33786 3231 34102 3232
rect 44733 3296 45049 3297
rect 44733 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45049 3296
rect 44733 3231 45049 3232
rect 29318 3166 31770 3226
rect 14457 3163 14523 3166
rect 19977 3163 20043 3166
rect 8753 3090 8819 3093
rect 22001 3090 22067 3093
rect 8753 3088 22067 3090
rect 8753 3032 8758 3088
rect 8814 3032 22006 3088
rect 22062 3032 22067 3088
rect 8753 3030 22067 3032
rect 8753 3027 8819 3030
rect 22001 3027 22067 3030
rect 24025 3090 24091 3093
rect 30741 3090 30807 3093
rect 24025 3088 30807 3090
rect 24025 3032 24030 3088
rect 24086 3032 30746 3088
rect 30802 3032 30807 3088
rect 24025 3030 30807 3032
rect 31710 3090 31770 3166
rect 37825 3090 37891 3093
rect 31710 3088 37891 3090
rect 31710 3032 37830 3088
rect 37886 3032 37891 3088
rect 31710 3030 37891 3032
rect 24025 3027 24091 3030
rect 30741 3027 30807 3030
rect 37825 3027 37891 3030
rect 9397 2954 9463 2957
rect 21541 2954 21607 2957
rect 9397 2952 21607 2954
rect 9397 2896 9402 2952
rect 9458 2896 21546 2952
rect 21602 2896 21607 2952
rect 9397 2894 21607 2896
rect 9397 2891 9463 2894
rect 21541 2891 21607 2894
rect 27981 2954 28047 2957
rect 35893 2954 35959 2957
rect 27981 2952 35959 2954
rect 27981 2896 27986 2952
rect 28042 2896 35898 2952
rect 35954 2896 35959 2952
rect 27981 2894 35959 2896
rect 27981 2891 28047 2894
rect 35893 2891 35959 2894
rect 6821 2818 6887 2821
rect 14457 2818 14523 2821
rect 6821 2816 14523 2818
rect 6821 2760 6826 2816
rect 6882 2760 14462 2816
rect 14518 2760 14523 2816
rect 6821 2758 14523 2760
rect 6821 2755 6887 2758
rect 14457 2755 14523 2758
rect 17953 2818 18019 2821
rect 19149 2818 19215 2821
rect 17953 2816 19215 2818
rect 17953 2760 17958 2816
rect 18014 2760 19154 2816
rect 19210 2760 19215 2816
rect 17953 2758 19215 2760
rect 17953 2755 18019 2758
rect 19149 2755 19215 2758
rect 28993 2818 29059 2821
rect 31753 2818 31819 2821
rect 28993 2816 31819 2818
rect 28993 2760 28998 2816
rect 29054 2760 31758 2816
rect 31814 2760 31819 2816
rect 28993 2758 31819 2760
rect 28993 2755 29059 2758
rect 31753 2755 31819 2758
rect 6419 2752 6735 2753
rect 6419 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6735 2752
rect 6419 2687 6735 2688
rect 17366 2752 17682 2753
rect 17366 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17682 2752
rect 17366 2687 17682 2688
rect 28313 2752 28629 2753
rect 28313 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28629 2752
rect 28313 2687 28629 2688
rect 39260 2752 39576 2753
rect 39260 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39576 2752
rect 39260 2687 39576 2688
rect 18321 2682 18387 2685
rect 19057 2682 19123 2685
rect 18321 2680 19123 2682
rect 18321 2624 18326 2680
rect 18382 2624 19062 2680
rect 19118 2624 19123 2680
rect 18321 2622 19123 2624
rect 18321 2619 18387 2622
rect 19057 2619 19123 2622
rect 19333 2682 19399 2685
rect 26509 2682 26575 2685
rect 19333 2680 26575 2682
rect 19333 2624 19338 2680
rect 19394 2624 26514 2680
rect 26570 2624 26575 2680
rect 19333 2622 26575 2624
rect 19333 2619 19399 2622
rect 26509 2619 26575 2622
rect 9949 2546 10015 2549
rect 21633 2546 21699 2549
rect 9949 2544 21699 2546
rect 9949 2488 9954 2544
rect 10010 2488 21638 2544
rect 21694 2488 21699 2544
rect 9949 2486 21699 2488
rect 9949 2483 10015 2486
rect 21633 2483 21699 2486
rect 26693 2546 26759 2549
rect 38101 2546 38167 2549
rect 26693 2544 38167 2546
rect 26693 2488 26698 2544
rect 26754 2488 38106 2544
rect 38162 2488 38167 2544
rect 26693 2486 38167 2488
rect 26693 2483 26759 2486
rect 38101 2483 38167 2486
rect 9581 2410 9647 2413
rect 18505 2410 18571 2413
rect 9581 2408 18571 2410
rect 9581 2352 9586 2408
rect 9642 2352 18510 2408
rect 18566 2352 18571 2408
rect 9581 2350 18571 2352
rect 9581 2347 9647 2350
rect 18505 2347 18571 2350
rect 24761 2410 24827 2413
rect 27613 2410 27679 2413
rect 36537 2410 36603 2413
rect 24761 2408 27538 2410
rect 24761 2352 24766 2408
rect 24822 2352 27538 2408
rect 24761 2350 27538 2352
rect 24761 2347 24827 2350
rect 12985 2274 13051 2277
rect 19333 2274 19399 2277
rect 12985 2272 19399 2274
rect 12985 2216 12990 2272
rect 13046 2216 19338 2272
rect 19394 2216 19399 2272
rect 12985 2214 19399 2216
rect 27478 2274 27538 2350
rect 27613 2408 36603 2410
rect 27613 2352 27618 2408
rect 27674 2352 36542 2408
rect 36598 2352 36603 2408
rect 27613 2350 36603 2352
rect 27613 2347 27679 2350
rect 36537 2347 36603 2350
rect 30373 2274 30439 2277
rect 30649 2274 30715 2277
rect 27478 2272 30439 2274
rect 27478 2216 30378 2272
rect 30434 2216 30439 2272
rect 27478 2214 30439 2216
rect 12985 2211 13051 2214
rect 19333 2211 19399 2214
rect 30373 2211 30439 2214
rect 30606 2272 30715 2274
rect 30606 2216 30654 2272
rect 30710 2216 30715 2272
rect 30606 2211 30715 2216
rect 11892 2208 12208 2209
rect 11892 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12208 2208
rect 11892 2143 12208 2144
rect 22839 2208 23155 2209
rect 22839 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23155 2208
rect 22839 2143 23155 2144
rect 30606 2138 30666 2211
rect 33786 2208 34102 2209
rect 33786 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34102 2208
rect 33786 2143 34102 2144
rect 44733 2208 45049 2209
rect 44733 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45049 2208
rect 44733 2143 45049 2144
rect 26374 2078 30666 2138
rect 31201 2138 31267 2141
rect 33409 2138 33475 2141
rect 31201 2136 33475 2138
rect 31201 2080 31206 2136
rect 31262 2080 33414 2136
rect 33470 2080 33475 2136
rect 31201 2078 33475 2080
rect 14181 2002 14247 2005
rect 26374 2002 26434 2078
rect 31201 2075 31267 2078
rect 33409 2075 33475 2078
rect 14181 2000 26434 2002
rect 14181 1944 14186 2000
rect 14242 1944 26434 2000
rect 14181 1942 26434 1944
rect 28993 2002 29059 2005
rect 40033 2002 40099 2005
rect 28993 2000 40099 2002
rect 28993 1944 28998 2000
rect 29054 1944 40038 2000
rect 40094 1944 40099 2000
rect 28993 1942 40099 1944
rect 14181 1939 14247 1942
rect 28993 1939 29059 1942
rect 40033 1939 40099 1942
rect 13077 1866 13143 1869
rect 32305 1866 32371 1869
rect 13077 1864 32371 1866
rect 13077 1808 13082 1864
rect 13138 1808 32310 1864
rect 32366 1808 32371 1864
rect 13077 1806 32371 1808
rect 13077 1803 13143 1806
rect 32305 1803 32371 1806
rect 10225 1730 10291 1733
rect 22461 1730 22527 1733
rect 10225 1728 22527 1730
rect 10225 1672 10230 1728
rect 10286 1672 22466 1728
rect 22522 1672 22527 1728
rect 10225 1670 22527 1672
rect 10225 1667 10291 1670
rect 22461 1667 22527 1670
rect 26785 1730 26851 1733
rect 37733 1730 37799 1733
rect 26785 1728 37799 1730
rect 26785 1672 26790 1728
rect 26846 1672 37738 1728
rect 37794 1672 37799 1728
rect 26785 1670 37799 1672
rect 26785 1667 26851 1670
rect 37733 1667 37799 1670
rect 22645 1594 22711 1597
rect 32213 1594 32279 1597
rect 22645 1592 32279 1594
rect 22645 1536 22650 1592
rect 22706 1536 32218 1592
rect 32274 1536 32279 1592
rect 22645 1534 32279 1536
rect 22645 1531 22711 1534
rect 32213 1531 32279 1534
rect 19149 1322 19215 1325
rect 32581 1322 32647 1325
rect 19149 1320 31770 1322
rect 19149 1264 19154 1320
rect 19210 1264 31770 1320
rect 19149 1262 31770 1264
rect 19149 1259 19215 1262
rect 15193 1186 15259 1189
rect 31710 1186 31770 1262
rect 32078 1320 32647 1322
rect 32078 1264 32586 1320
rect 32642 1264 32647 1320
rect 32078 1262 32647 1264
rect 31886 1186 31892 1188
rect 15193 1184 26986 1186
rect 15193 1128 15198 1184
rect 15254 1128 26986 1184
rect 15193 1126 26986 1128
rect 31710 1126 31892 1186
rect 15193 1123 15259 1126
rect 7097 1050 7163 1053
rect 24894 1050 24900 1052
rect 7097 1048 24900 1050
rect 7097 992 7102 1048
rect 7158 992 24900 1048
rect 7097 990 24900 992
rect 7097 987 7163 990
rect 24894 988 24900 990
rect 24964 988 24970 1052
rect 26926 1050 26986 1126
rect 31886 1124 31892 1126
rect 31956 1124 31962 1188
rect 32078 1050 32138 1262
rect 32581 1259 32647 1262
rect 26926 990 32138 1050
rect 18781 100 18847 101
rect 19057 100 19123 101
rect 18781 98 18828 100
rect 18736 96 18828 98
rect 18736 40 18786 96
rect 18736 38 18828 40
rect 18781 36 18828 38
rect 18892 36 18898 100
rect 19006 36 19012 100
rect 19076 98 19123 100
rect 19076 96 19168 98
rect 19118 40 19168 96
rect 19076 38 19168 40
rect 19076 36 19123 38
rect 18781 35 18847 36
rect 19057 35 19123 36
<< via3 >>
rect 11898 7644 11962 7648
rect 11898 7588 11902 7644
rect 11902 7588 11958 7644
rect 11958 7588 11962 7644
rect 11898 7584 11962 7588
rect 11978 7644 12042 7648
rect 11978 7588 11982 7644
rect 11982 7588 12038 7644
rect 12038 7588 12042 7644
rect 11978 7584 12042 7588
rect 12058 7644 12122 7648
rect 12058 7588 12062 7644
rect 12062 7588 12118 7644
rect 12118 7588 12122 7644
rect 12058 7584 12122 7588
rect 12138 7644 12202 7648
rect 12138 7588 12142 7644
rect 12142 7588 12198 7644
rect 12198 7588 12202 7644
rect 12138 7584 12202 7588
rect 22845 7644 22909 7648
rect 22845 7588 22849 7644
rect 22849 7588 22905 7644
rect 22905 7588 22909 7644
rect 22845 7584 22909 7588
rect 22925 7644 22989 7648
rect 22925 7588 22929 7644
rect 22929 7588 22985 7644
rect 22985 7588 22989 7644
rect 22925 7584 22989 7588
rect 23005 7644 23069 7648
rect 23005 7588 23009 7644
rect 23009 7588 23065 7644
rect 23065 7588 23069 7644
rect 23005 7584 23069 7588
rect 23085 7644 23149 7648
rect 23085 7588 23089 7644
rect 23089 7588 23145 7644
rect 23145 7588 23149 7644
rect 23085 7584 23149 7588
rect 33792 7644 33856 7648
rect 33792 7588 33796 7644
rect 33796 7588 33852 7644
rect 33852 7588 33856 7644
rect 33792 7584 33856 7588
rect 33872 7644 33936 7648
rect 33872 7588 33876 7644
rect 33876 7588 33932 7644
rect 33932 7588 33936 7644
rect 33872 7584 33936 7588
rect 33952 7644 34016 7648
rect 33952 7588 33956 7644
rect 33956 7588 34012 7644
rect 34012 7588 34016 7644
rect 33952 7584 34016 7588
rect 34032 7644 34096 7648
rect 34032 7588 34036 7644
rect 34036 7588 34092 7644
rect 34092 7588 34096 7644
rect 34032 7584 34096 7588
rect 44739 7644 44803 7648
rect 44739 7588 44743 7644
rect 44743 7588 44799 7644
rect 44799 7588 44803 7644
rect 44739 7584 44803 7588
rect 44819 7644 44883 7648
rect 44819 7588 44823 7644
rect 44823 7588 44879 7644
rect 44879 7588 44883 7644
rect 44819 7584 44883 7588
rect 44899 7644 44963 7648
rect 44899 7588 44903 7644
rect 44903 7588 44959 7644
rect 44959 7588 44963 7644
rect 44899 7584 44963 7588
rect 44979 7644 45043 7648
rect 44979 7588 44983 7644
rect 44983 7588 45039 7644
rect 45039 7588 45043 7644
rect 44979 7584 45043 7588
rect 6425 7100 6489 7104
rect 6425 7044 6429 7100
rect 6429 7044 6485 7100
rect 6485 7044 6489 7100
rect 6425 7040 6489 7044
rect 6505 7100 6569 7104
rect 6505 7044 6509 7100
rect 6509 7044 6565 7100
rect 6565 7044 6569 7100
rect 6505 7040 6569 7044
rect 6585 7100 6649 7104
rect 6585 7044 6589 7100
rect 6589 7044 6645 7100
rect 6645 7044 6649 7100
rect 6585 7040 6649 7044
rect 6665 7100 6729 7104
rect 6665 7044 6669 7100
rect 6669 7044 6725 7100
rect 6725 7044 6729 7100
rect 6665 7040 6729 7044
rect 17372 7100 17436 7104
rect 17372 7044 17376 7100
rect 17376 7044 17432 7100
rect 17432 7044 17436 7100
rect 17372 7040 17436 7044
rect 17452 7100 17516 7104
rect 17452 7044 17456 7100
rect 17456 7044 17512 7100
rect 17512 7044 17516 7100
rect 17452 7040 17516 7044
rect 17532 7100 17596 7104
rect 17532 7044 17536 7100
rect 17536 7044 17592 7100
rect 17592 7044 17596 7100
rect 17532 7040 17596 7044
rect 17612 7100 17676 7104
rect 17612 7044 17616 7100
rect 17616 7044 17672 7100
rect 17672 7044 17676 7100
rect 17612 7040 17676 7044
rect 28319 7100 28383 7104
rect 28319 7044 28323 7100
rect 28323 7044 28379 7100
rect 28379 7044 28383 7100
rect 28319 7040 28383 7044
rect 28399 7100 28463 7104
rect 28399 7044 28403 7100
rect 28403 7044 28459 7100
rect 28459 7044 28463 7100
rect 28399 7040 28463 7044
rect 28479 7100 28543 7104
rect 28479 7044 28483 7100
rect 28483 7044 28539 7100
rect 28539 7044 28543 7100
rect 28479 7040 28543 7044
rect 28559 7100 28623 7104
rect 28559 7044 28563 7100
rect 28563 7044 28619 7100
rect 28619 7044 28623 7100
rect 28559 7040 28623 7044
rect 39266 7100 39330 7104
rect 39266 7044 39270 7100
rect 39270 7044 39326 7100
rect 39326 7044 39330 7100
rect 39266 7040 39330 7044
rect 39346 7100 39410 7104
rect 39346 7044 39350 7100
rect 39350 7044 39406 7100
rect 39406 7044 39410 7100
rect 39346 7040 39410 7044
rect 39426 7100 39490 7104
rect 39426 7044 39430 7100
rect 39430 7044 39486 7100
rect 39486 7044 39490 7100
rect 39426 7040 39490 7044
rect 39506 7100 39570 7104
rect 39506 7044 39510 7100
rect 39510 7044 39566 7100
rect 39566 7044 39570 7100
rect 39506 7040 39570 7044
rect 11898 6556 11962 6560
rect 11898 6500 11902 6556
rect 11902 6500 11958 6556
rect 11958 6500 11962 6556
rect 11898 6496 11962 6500
rect 11978 6556 12042 6560
rect 11978 6500 11982 6556
rect 11982 6500 12038 6556
rect 12038 6500 12042 6556
rect 11978 6496 12042 6500
rect 12058 6556 12122 6560
rect 12058 6500 12062 6556
rect 12062 6500 12118 6556
rect 12118 6500 12122 6556
rect 12058 6496 12122 6500
rect 12138 6556 12202 6560
rect 12138 6500 12142 6556
rect 12142 6500 12198 6556
rect 12198 6500 12202 6556
rect 12138 6496 12202 6500
rect 22845 6556 22909 6560
rect 22845 6500 22849 6556
rect 22849 6500 22905 6556
rect 22905 6500 22909 6556
rect 22845 6496 22909 6500
rect 22925 6556 22989 6560
rect 22925 6500 22929 6556
rect 22929 6500 22985 6556
rect 22985 6500 22989 6556
rect 22925 6496 22989 6500
rect 23005 6556 23069 6560
rect 23005 6500 23009 6556
rect 23009 6500 23065 6556
rect 23065 6500 23069 6556
rect 23005 6496 23069 6500
rect 23085 6556 23149 6560
rect 23085 6500 23089 6556
rect 23089 6500 23145 6556
rect 23145 6500 23149 6556
rect 23085 6496 23149 6500
rect 33792 6556 33856 6560
rect 33792 6500 33796 6556
rect 33796 6500 33852 6556
rect 33852 6500 33856 6556
rect 33792 6496 33856 6500
rect 33872 6556 33936 6560
rect 33872 6500 33876 6556
rect 33876 6500 33932 6556
rect 33932 6500 33936 6556
rect 33872 6496 33936 6500
rect 33952 6556 34016 6560
rect 33952 6500 33956 6556
rect 33956 6500 34012 6556
rect 34012 6500 34016 6556
rect 33952 6496 34016 6500
rect 34032 6556 34096 6560
rect 34032 6500 34036 6556
rect 34036 6500 34092 6556
rect 34092 6500 34096 6556
rect 34032 6496 34096 6500
rect 44739 6556 44803 6560
rect 44739 6500 44743 6556
rect 44743 6500 44799 6556
rect 44799 6500 44803 6556
rect 44739 6496 44803 6500
rect 44819 6556 44883 6560
rect 44819 6500 44823 6556
rect 44823 6500 44879 6556
rect 44879 6500 44883 6556
rect 44819 6496 44883 6500
rect 44899 6556 44963 6560
rect 44899 6500 44903 6556
rect 44903 6500 44959 6556
rect 44959 6500 44963 6556
rect 44899 6496 44963 6500
rect 44979 6556 45043 6560
rect 44979 6500 44983 6556
rect 44983 6500 45039 6556
rect 45039 6500 45043 6556
rect 44979 6496 45043 6500
rect 6425 6012 6489 6016
rect 6425 5956 6429 6012
rect 6429 5956 6485 6012
rect 6485 5956 6489 6012
rect 6425 5952 6489 5956
rect 6505 6012 6569 6016
rect 6505 5956 6509 6012
rect 6509 5956 6565 6012
rect 6565 5956 6569 6012
rect 6505 5952 6569 5956
rect 6585 6012 6649 6016
rect 6585 5956 6589 6012
rect 6589 5956 6645 6012
rect 6645 5956 6649 6012
rect 6585 5952 6649 5956
rect 6665 6012 6729 6016
rect 6665 5956 6669 6012
rect 6669 5956 6725 6012
rect 6725 5956 6729 6012
rect 6665 5952 6729 5956
rect 17372 6012 17436 6016
rect 17372 5956 17376 6012
rect 17376 5956 17432 6012
rect 17432 5956 17436 6012
rect 17372 5952 17436 5956
rect 17452 6012 17516 6016
rect 17452 5956 17456 6012
rect 17456 5956 17512 6012
rect 17512 5956 17516 6012
rect 17452 5952 17516 5956
rect 17532 6012 17596 6016
rect 17532 5956 17536 6012
rect 17536 5956 17592 6012
rect 17592 5956 17596 6012
rect 17532 5952 17596 5956
rect 17612 6012 17676 6016
rect 17612 5956 17616 6012
rect 17616 5956 17672 6012
rect 17672 5956 17676 6012
rect 17612 5952 17676 5956
rect 28319 6012 28383 6016
rect 28319 5956 28323 6012
rect 28323 5956 28379 6012
rect 28379 5956 28383 6012
rect 28319 5952 28383 5956
rect 28399 6012 28463 6016
rect 28399 5956 28403 6012
rect 28403 5956 28459 6012
rect 28459 5956 28463 6012
rect 28399 5952 28463 5956
rect 28479 6012 28543 6016
rect 28479 5956 28483 6012
rect 28483 5956 28539 6012
rect 28539 5956 28543 6012
rect 28479 5952 28543 5956
rect 28559 6012 28623 6016
rect 28559 5956 28563 6012
rect 28563 5956 28619 6012
rect 28619 5956 28623 6012
rect 28559 5952 28623 5956
rect 39266 6012 39330 6016
rect 39266 5956 39270 6012
rect 39270 5956 39326 6012
rect 39326 5956 39330 6012
rect 39266 5952 39330 5956
rect 39346 6012 39410 6016
rect 39346 5956 39350 6012
rect 39350 5956 39406 6012
rect 39406 5956 39410 6012
rect 39346 5952 39410 5956
rect 39426 6012 39490 6016
rect 39426 5956 39430 6012
rect 39430 5956 39486 6012
rect 39486 5956 39490 6012
rect 39426 5952 39490 5956
rect 39506 6012 39570 6016
rect 39506 5956 39510 6012
rect 39510 5956 39566 6012
rect 39566 5956 39570 6012
rect 39506 5952 39570 5956
rect 11898 5468 11962 5472
rect 11898 5412 11902 5468
rect 11902 5412 11958 5468
rect 11958 5412 11962 5468
rect 11898 5408 11962 5412
rect 11978 5468 12042 5472
rect 11978 5412 11982 5468
rect 11982 5412 12038 5468
rect 12038 5412 12042 5468
rect 11978 5408 12042 5412
rect 12058 5468 12122 5472
rect 12058 5412 12062 5468
rect 12062 5412 12118 5468
rect 12118 5412 12122 5468
rect 12058 5408 12122 5412
rect 12138 5468 12202 5472
rect 12138 5412 12142 5468
rect 12142 5412 12198 5468
rect 12198 5412 12202 5468
rect 12138 5408 12202 5412
rect 22845 5468 22909 5472
rect 22845 5412 22849 5468
rect 22849 5412 22905 5468
rect 22905 5412 22909 5468
rect 22845 5408 22909 5412
rect 22925 5468 22989 5472
rect 22925 5412 22929 5468
rect 22929 5412 22985 5468
rect 22985 5412 22989 5468
rect 22925 5408 22989 5412
rect 23005 5468 23069 5472
rect 23005 5412 23009 5468
rect 23009 5412 23065 5468
rect 23065 5412 23069 5468
rect 23005 5408 23069 5412
rect 23085 5468 23149 5472
rect 23085 5412 23089 5468
rect 23089 5412 23145 5468
rect 23145 5412 23149 5468
rect 23085 5408 23149 5412
rect 33792 5468 33856 5472
rect 33792 5412 33796 5468
rect 33796 5412 33852 5468
rect 33852 5412 33856 5468
rect 33792 5408 33856 5412
rect 33872 5468 33936 5472
rect 33872 5412 33876 5468
rect 33876 5412 33932 5468
rect 33932 5412 33936 5468
rect 33872 5408 33936 5412
rect 33952 5468 34016 5472
rect 33952 5412 33956 5468
rect 33956 5412 34012 5468
rect 34012 5412 34016 5468
rect 33952 5408 34016 5412
rect 34032 5468 34096 5472
rect 34032 5412 34036 5468
rect 34036 5412 34092 5468
rect 34092 5412 34096 5468
rect 34032 5408 34096 5412
rect 44739 5468 44803 5472
rect 44739 5412 44743 5468
rect 44743 5412 44799 5468
rect 44799 5412 44803 5468
rect 44739 5408 44803 5412
rect 44819 5468 44883 5472
rect 44819 5412 44823 5468
rect 44823 5412 44879 5468
rect 44879 5412 44883 5468
rect 44819 5408 44883 5412
rect 44899 5468 44963 5472
rect 44899 5412 44903 5468
rect 44903 5412 44959 5468
rect 44959 5412 44963 5468
rect 44899 5408 44963 5412
rect 44979 5468 45043 5472
rect 44979 5412 44983 5468
rect 44983 5412 45039 5468
rect 45039 5412 45043 5468
rect 44979 5408 45043 5412
rect 6425 4924 6489 4928
rect 6425 4868 6429 4924
rect 6429 4868 6485 4924
rect 6485 4868 6489 4924
rect 6425 4864 6489 4868
rect 6505 4924 6569 4928
rect 6505 4868 6509 4924
rect 6509 4868 6565 4924
rect 6565 4868 6569 4924
rect 6505 4864 6569 4868
rect 6585 4924 6649 4928
rect 6585 4868 6589 4924
rect 6589 4868 6645 4924
rect 6645 4868 6649 4924
rect 6585 4864 6649 4868
rect 6665 4924 6729 4928
rect 6665 4868 6669 4924
rect 6669 4868 6725 4924
rect 6725 4868 6729 4924
rect 6665 4864 6729 4868
rect 17372 4924 17436 4928
rect 17372 4868 17376 4924
rect 17376 4868 17432 4924
rect 17432 4868 17436 4924
rect 17372 4864 17436 4868
rect 17452 4924 17516 4928
rect 17452 4868 17456 4924
rect 17456 4868 17512 4924
rect 17512 4868 17516 4924
rect 17452 4864 17516 4868
rect 17532 4924 17596 4928
rect 17532 4868 17536 4924
rect 17536 4868 17592 4924
rect 17592 4868 17596 4924
rect 17532 4864 17596 4868
rect 17612 4924 17676 4928
rect 17612 4868 17616 4924
rect 17616 4868 17672 4924
rect 17672 4868 17676 4924
rect 17612 4864 17676 4868
rect 28319 4924 28383 4928
rect 28319 4868 28323 4924
rect 28323 4868 28379 4924
rect 28379 4868 28383 4924
rect 28319 4864 28383 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 39266 4924 39330 4928
rect 39266 4868 39270 4924
rect 39270 4868 39326 4924
rect 39326 4868 39330 4924
rect 39266 4864 39330 4868
rect 39346 4924 39410 4928
rect 39346 4868 39350 4924
rect 39350 4868 39406 4924
rect 39406 4868 39410 4924
rect 39346 4864 39410 4868
rect 39426 4924 39490 4928
rect 39426 4868 39430 4924
rect 39430 4868 39486 4924
rect 39486 4868 39490 4924
rect 39426 4864 39490 4868
rect 39506 4924 39570 4928
rect 39506 4868 39510 4924
rect 39510 4868 39566 4924
rect 39566 4868 39570 4924
rect 39506 4864 39570 4868
rect 11898 4380 11962 4384
rect 11898 4324 11902 4380
rect 11902 4324 11958 4380
rect 11958 4324 11962 4380
rect 11898 4320 11962 4324
rect 11978 4380 12042 4384
rect 11978 4324 11982 4380
rect 11982 4324 12038 4380
rect 12038 4324 12042 4380
rect 11978 4320 12042 4324
rect 12058 4380 12122 4384
rect 12058 4324 12062 4380
rect 12062 4324 12118 4380
rect 12118 4324 12122 4380
rect 12058 4320 12122 4324
rect 12138 4380 12202 4384
rect 12138 4324 12142 4380
rect 12142 4324 12198 4380
rect 12198 4324 12202 4380
rect 12138 4320 12202 4324
rect 22845 4380 22909 4384
rect 22845 4324 22849 4380
rect 22849 4324 22905 4380
rect 22905 4324 22909 4380
rect 22845 4320 22909 4324
rect 22925 4380 22989 4384
rect 22925 4324 22929 4380
rect 22929 4324 22985 4380
rect 22985 4324 22989 4380
rect 22925 4320 22989 4324
rect 23005 4380 23069 4384
rect 23005 4324 23009 4380
rect 23009 4324 23065 4380
rect 23065 4324 23069 4380
rect 23005 4320 23069 4324
rect 23085 4380 23149 4384
rect 23085 4324 23089 4380
rect 23089 4324 23145 4380
rect 23145 4324 23149 4380
rect 23085 4320 23149 4324
rect 33792 4380 33856 4384
rect 33792 4324 33796 4380
rect 33796 4324 33852 4380
rect 33852 4324 33856 4380
rect 33792 4320 33856 4324
rect 33872 4380 33936 4384
rect 33872 4324 33876 4380
rect 33876 4324 33932 4380
rect 33932 4324 33936 4380
rect 33872 4320 33936 4324
rect 33952 4380 34016 4384
rect 33952 4324 33956 4380
rect 33956 4324 34012 4380
rect 34012 4324 34016 4380
rect 33952 4320 34016 4324
rect 34032 4380 34096 4384
rect 34032 4324 34036 4380
rect 34036 4324 34092 4380
rect 34092 4324 34096 4380
rect 34032 4320 34096 4324
rect 44739 4380 44803 4384
rect 44739 4324 44743 4380
rect 44743 4324 44799 4380
rect 44799 4324 44803 4380
rect 44739 4320 44803 4324
rect 44819 4380 44883 4384
rect 44819 4324 44823 4380
rect 44823 4324 44879 4380
rect 44879 4324 44883 4380
rect 44819 4320 44883 4324
rect 44899 4380 44963 4384
rect 44899 4324 44903 4380
rect 44903 4324 44959 4380
rect 44959 4324 44963 4380
rect 44899 4320 44963 4324
rect 44979 4380 45043 4384
rect 44979 4324 44983 4380
rect 44983 4324 45039 4380
rect 45039 4324 45043 4380
rect 44979 4320 45043 4324
rect 18828 4252 18892 4316
rect 19288 3904 19352 3908
rect 19288 3848 19302 3904
rect 19302 3848 19352 3904
rect 19288 3844 19352 3848
rect 6425 3836 6489 3840
rect 6425 3780 6429 3836
rect 6429 3780 6485 3836
rect 6485 3780 6489 3836
rect 6425 3776 6489 3780
rect 6505 3836 6569 3840
rect 6505 3780 6509 3836
rect 6509 3780 6565 3836
rect 6565 3780 6569 3836
rect 6505 3776 6569 3780
rect 6585 3836 6649 3840
rect 6585 3780 6589 3836
rect 6589 3780 6645 3836
rect 6645 3780 6649 3836
rect 6585 3776 6649 3780
rect 6665 3836 6729 3840
rect 6665 3780 6669 3836
rect 6669 3780 6725 3836
rect 6725 3780 6729 3836
rect 6665 3776 6729 3780
rect 17372 3836 17436 3840
rect 17372 3780 17376 3836
rect 17376 3780 17432 3836
rect 17432 3780 17436 3836
rect 17372 3776 17436 3780
rect 17452 3836 17516 3840
rect 17452 3780 17456 3836
rect 17456 3780 17512 3836
rect 17512 3780 17516 3836
rect 17452 3776 17516 3780
rect 17532 3836 17596 3840
rect 17532 3780 17536 3836
rect 17536 3780 17592 3836
rect 17592 3780 17596 3836
rect 17532 3776 17596 3780
rect 17612 3836 17676 3840
rect 17612 3780 17616 3836
rect 17616 3780 17672 3836
rect 17672 3780 17676 3836
rect 17612 3776 17676 3780
rect 28319 3836 28383 3840
rect 28319 3780 28323 3836
rect 28323 3780 28379 3836
rect 28379 3780 28383 3836
rect 28319 3776 28383 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 39266 3836 39330 3840
rect 39266 3780 39270 3836
rect 39270 3780 39326 3836
rect 39326 3780 39330 3836
rect 39266 3776 39330 3780
rect 39346 3836 39410 3840
rect 39346 3780 39350 3836
rect 39350 3780 39406 3836
rect 39406 3780 39410 3836
rect 39346 3776 39410 3780
rect 39426 3836 39490 3840
rect 39426 3780 39430 3836
rect 39430 3780 39486 3836
rect 39486 3780 39490 3836
rect 39426 3776 39490 3780
rect 39506 3836 39570 3840
rect 39506 3780 39510 3836
rect 39510 3780 39566 3836
rect 39566 3780 39570 3836
rect 39506 3776 39570 3780
rect 24900 3436 24964 3500
rect 31892 3436 31956 3500
rect 11898 3292 11962 3296
rect 11898 3236 11902 3292
rect 11902 3236 11958 3292
rect 11958 3236 11962 3292
rect 11898 3232 11962 3236
rect 11978 3292 12042 3296
rect 11978 3236 11982 3292
rect 11982 3236 12038 3292
rect 12038 3236 12042 3292
rect 11978 3232 12042 3236
rect 12058 3292 12122 3296
rect 12058 3236 12062 3292
rect 12062 3236 12118 3292
rect 12118 3236 12122 3292
rect 12058 3232 12122 3236
rect 12138 3292 12202 3296
rect 12138 3236 12142 3292
rect 12142 3236 12198 3292
rect 12198 3236 12202 3292
rect 12138 3232 12202 3236
rect 22845 3292 22909 3296
rect 22845 3236 22849 3292
rect 22849 3236 22905 3292
rect 22905 3236 22909 3292
rect 22845 3232 22909 3236
rect 22925 3292 22989 3296
rect 22925 3236 22929 3292
rect 22929 3236 22985 3292
rect 22985 3236 22989 3292
rect 22925 3232 22989 3236
rect 23005 3292 23069 3296
rect 23005 3236 23009 3292
rect 23009 3236 23065 3292
rect 23065 3236 23069 3292
rect 23005 3232 23069 3236
rect 23085 3292 23149 3296
rect 23085 3236 23089 3292
rect 23089 3236 23145 3292
rect 23145 3236 23149 3292
rect 23085 3232 23149 3236
rect 33792 3292 33856 3296
rect 33792 3236 33796 3292
rect 33796 3236 33852 3292
rect 33852 3236 33856 3292
rect 33792 3232 33856 3236
rect 33872 3292 33936 3296
rect 33872 3236 33876 3292
rect 33876 3236 33932 3292
rect 33932 3236 33936 3292
rect 33872 3232 33936 3236
rect 33952 3292 34016 3296
rect 33952 3236 33956 3292
rect 33956 3236 34012 3292
rect 34012 3236 34016 3292
rect 33952 3232 34016 3236
rect 34032 3292 34096 3296
rect 34032 3236 34036 3292
rect 34036 3236 34092 3292
rect 34092 3236 34096 3292
rect 34032 3232 34096 3236
rect 44739 3292 44803 3296
rect 44739 3236 44743 3292
rect 44743 3236 44799 3292
rect 44799 3236 44803 3292
rect 44739 3232 44803 3236
rect 44819 3292 44883 3296
rect 44819 3236 44823 3292
rect 44823 3236 44879 3292
rect 44879 3236 44883 3292
rect 44819 3232 44883 3236
rect 44899 3292 44963 3296
rect 44899 3236 44903 3292
rect 44903 3236 44959 3292
rect 44959 3236 44963 3292
rect 44899 3232 44963 3236
rect 44979 3292 45043 3296
rect 44979 3236 44983 3292
rect 44983 3236 45039 3292
rect 45039 3236 45043 3292
rect 44979 3232 45043 3236
rect 6425 2748 6489 2752
rect 6425 2692 6429 2748
rect 6429 2692 6485 2748
rect 6485 2692 6489 2748
rect 6425 2688 6489 2692
rect 6505 2748 6569 2752
rect 6505 2692 6509 2748
rect 6509 2692 6565 2748
rect 6565 2692 6569 2748
rect 6505 2688 6569 2692
rect 6585 2748 6649 2752
rect 6585 2692 6589 2748
rect 6589 2692 6645 2748
rect 6645 2692 6649 2748
rect 6585 2688 6649 2692
rect 6665 2748 6729 2752
rect 6665 2692 6669 2748
rect 6669 2692 6725 2748
rect 6725 2692 6729 2748
rect 6665 2688 6729 2692
rect 17372 2748 17436 2752
rect 17372 2692 17376 2748
rect 17376 2692 17432 2748
rect 17432 2692 17436 2748
rect 17372 2688 17436 2692
rect 17452 2748 17516 2752
rect 17452 2692 17456 2748
rect 17456 2692 17512 2748
rect 17512 2692 17516 2748
rect 17452 2688 17516 2692
rect 17532 2748 17596 2752
rect 17532 2692 17536 2748
rect 17536 2692 17592 2748
rect 17592 2692 17596 2748
rect 17532 2688 17596 2692
rect 17612 2748 17676 2752
rect 17612 2692 17616 2748
rect 17616 2692 17672 2748
rect 17672 2692 17676 2748
rect 17612 2688 17676 2692
rect 28319 2748 28383 2752
rect 28319 2692 28323 2748
rect 28323 2692 28379 2748
rect 28379 2692 28383 2748
rect 28319 2688 28383 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 39266 2748 39330 2752
rect 39266 2692 39270 2748
rect 39270 2692 39326 2748
rect 39326 2692 39330 2748
rect 39266 2688 39330 2692
rect 39346 2748 39410 2752
rect 39346 2692 39350 2748
rect 39350 2692 39406 2748
rect 39406 2692 39410 2748
rect 39346 2688 39410 2692
rect 39426 2748 39490 2752
rect 39426 2692 39430 2748
rect 39430 2692 39486 2748
rect 39486 2692 39490 2748
rect 39426 2688 39490 2692
rect 39506 2748 39570 2752
rect 39506 2692 39510 2748
rect 39510 2692 39566 2748
rect 39566 2692 39570 2748
rect 39506 2688 39570 2692
rect 11898 2204 11962 2208
rect 11898 2148 11902 2204
rect 11902 2148 11958 2204
rect 11958 2148 11962 2204
rect 11898 2144 11962 2148
rect 11978 2204 12042 2208
rect 11978 2148 11982 2204
rect 11982 2148 12038 2204
rect 12038 2148 12042 2204
rect 11978 2144 12042 2148
rect 12058 2204 12122 2208
rect 12058 2148 12062 2204
rect 12062 2148 12118 2204
rect 12118 2148 12122 2204
rect 12058 2144 12122 2148
rect 12138 2204 12202 2208
rect 12138 2148 12142 2204
rect 12142 2148 12198 2204
rect 12198 2148 12202 2204
rect 12138 2144 12202 2148
rect 22845 2204 22909 2208
rect 22845 2148 22849 2204
rect 22849 2148 22905 2204
rect 22905 2148 22909 2204
rect 22845 2144 22909 2148
rect 22925 2204 22989 2208
rect 22925 2148 22929 2204
rect 22929 2148 22985 2204
rect 22985 2148 22989 2204
rect 22925 2144 22989 2148
rect 23005 2204 23069 2208
rect 23005 2148 23009 2204
rect 23009 2148 23065 2204
rect 23065 2148 23069 2204
rect 23005 2144 23069 2148
rect 23085 2204 23149 2208
rect 23085 2148 23089 2204
rect 23089 2148 23145 2204
rect 23145 2148 23149 2204
rect 23085 2144 23149 2148
rect 33792 2204 33856 2208
rect 33792 2148 33796 2204
rect 33796 2148 33852 2204
rect 33852 2148 33856 2204
rect 33792 2144 33856 2148
rect 33872 2204 33936 2208
rect 33872 2148 33876 2204
rect 33876 2148 33932 2204
rect 33932 2148 33936 2204
rect 33872 2144 33936 2148
rect 33952 2204 34016 2208
rect 33952 2148 33956 2204
rect 33956 2148 34012 2204
rect 34012 2148 34016 2204
rect 33952 2144 34016 2148
rect 34032 2204 34096 2208
rect 34032 2148 34036 2204
rect 34036 2148 34092 2204
rect 34092 2148 34096 2204
rect 34032 2144 34096 2148
rect 44739 2204 44803 2208
rect 44739 2148 44743 2204
rect 44743 2148 44799 2204
rect 44799 2148 44803 2204
rect 44739 2144 44803 2148
rect 44819 2204 44883 2208
rect 44819 2148 44823 2204
rect 44823 2148 44879 2204
rect 44879 2148 44883 2204
rect 44819 2144 44883 2148
rect 44899 2204 44963 2208
rect 44899 2148 44903 2204
rect 44903 2148 44959 2204
rect 44959 2148 44963 2204
rect 44899 2144 44963 2148
rect 44979 2204 45043 2208
rect 44979 2148 44983 2204
rect 44983 2148 45039 2204
rect 45039 2148 45043 2204
rect 44979 2144 45043 2148
rect 24900 988 24964 1052
rect 31892 1124 31956 1188
rect 18828 96 18892 100
rect 18828 40 18842 96
rect 18842 40 18892 96
rect 18828 36 18892 40
rect 19012 96 19076 100
rect 19012 40 19062 96
rect 19062 40 19076 96
rect 19012 36 19076 40
<< metal4 >>
rect 6417 7104 6737 7664
rect 6417 7040 6425 7104
rect 6489 7040 6505 7104
rect 6569 7040 6585 7104
rect 6649 7040 6665 7104
rect 6729 7040 6737 7104
rect 6417 6016 6737 7040
rect 6417 5952 6425 6016
rect 6489 5952 6505 6016
rect 6569 5952 6585 6016
rect 6649 5952 6665 6016
rect 6729 5952 6737 6016
rect 6417 4928 6737 5952
rect 6417 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6737 4928
rect 6417 3840 6737 4864
rect 6417 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6737 3840
rect 6417 2752 6737 3776
rect 6417 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6737 2752
rect 6417 2128 6737 2688
rect 11890 7648 12210 7664
rect 11890 7584 11898 7648
rect 11962 7584 11978 7648
rect 12042 7584 12058 7648
rect 12122 7584 12138 7648
rect 12202 7584 12210 7648
rect 11890 6560 12210 7584
rect 11890 6496 11898 6560
rect 11962 6496 11978 6560
rect 12042 6496 12058 6560
rect 12122 6496 12138 6560
rect 12202 6496 12210 6560
rect 11890 5472 12210 6496
rect 11890 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12210 5472
rect 11890 4384 12210 5408
rect 11890 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12210 4384
rect 11890 3296 12210 4320
rect 11890 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12210 3296
rect 11890 2208 12210 3232
rect 11890 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12210 2208
rect 11890 2128 12210 2144
rect 17364 7104 17684 7664
rect 17364 7040 17372 7104
rect 17436 7040 17452 7104
rect 17516 7040 17532 7104
rect 17596 7040 17612 7104
rect 17676 7040 17684 7104
rect 17364 6016 17684 7040
rect 17364 5952 17372 6016
rect 17436 5952 17452 6016
rect 17516 5952 17532 6016
rect 17596 5952 17612 6016
rect 17676 5952 17684 6016
rect 17364 4928 17684 5952
rect 17364 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17684 4928
rect 17364 3840 17684 4864
rect 22837 7648 23157 7664
rect 22837 7584 22845 7648
rect 22909 7584 22925 7648
rect 22989 7584 23005 7648
rect 23069 7584 23085 7648
rect 23149 7584 23157 7648
rect 22837 6560 23157 7584
rect 22837 6496 22845 6560
rect 22909 6496 22925 6560
rect 22989 6496 23005 6560
rect 23069 6496 23085 6560
rect 23149 6496 23157 6560
rect 22837 5472 23157 6496
rect 22837 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23157 5472
rect 22837 4384 23157 5408
rect 22837 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23157 4384
rect 18827 4316 18893 4317
rect 18827 4252 18828 4316
rect 18892 4252 18893 4316
rect 18827 4251 18893 4252
rect 17364 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17684 3840
rect 17364 2752 17684 3776
rect 17364 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17684 2752
rect 17364 2128 17684 2688
rect 18830 101 18890 4251
rect 19287 3908 19353 3909
rect 19287 3844 19288 3908
rect 19352 3844 19353 3908
rect 19287 3843 19353 3844
rect 19290 3770 19350 3843
rect 19014 3710 19350 3770
rect 19014 101 19074 3710
rect 22837 3296 23157 4320
rect 28311 7104 28631 7664
rect 28311 7040 28319 7104
rect 28383 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28631 7104
rect 28311 6016 28631 7040
rect 28311 5952 28319 6016
rect 28383 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28631 6016
rect 28311 4928 28631 5952
rect 28311 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28631 4928
rect 28311 3840 28631 4864
rect 28311 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28631 3840
rect 24899 3500 24965 3501
rect 24899 3436 24900 3500
rect 24964 3436 24965 3500
rect 24899 3435 24965 3436
rect 22837 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23157 3296
rect 22837 2208 23157 3232
rect 22837 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23157 2208
rect 22837 2128 23157 2144
rect 24902 1053 24962 3435
rect 28311 2752 28631 3776
rect 33784 7648 34104 7664
rect 33784 7584 33792 7648
rect 33856 7584 33872 7648
rect 33936 7584 33952 7648
rect 34016 7584 34032 7648
rect 34096 7584 34104 7648
rect 33784 6560 34104 7584
rect 33784 6496 33792 6560
rect 33856 6496 33872 6560
rect 33936 6496 33952 6560
rect 34016 6496 34032 6560
rect 34096 6496 34104 6560
rect 33784 5472 34104 6496
rect 33784 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34104 5472
rect 33784 4384 34104 5408
rect 33784 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34104 4384
rect 31891 3500 31957 3501
rect 31891 3436 31892 3500
rect 31956 3436 31957 3500
rect 31891 3435 31957 3436
rect 28311 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28631 2752
rect 28311 2128 28631 2688
rect 31894 1189 31954 3435
rect 33784 3296 34104 4320
rect 33784 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34104 3296
rect 33784 2208 34104 3232
rect 33784 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34104 2208
rect 33784 2128 34104 2144
rect 39258 7104 39578 7664
rect 39258 7040 39266 7104
rect 39330 7040 39346 7104
rect 39410 7040 39426 7104
rect 39490 7040 39506 7104
rect 39570 7040 39578 7104
rect 39258 6016 39578 7040
rect 39258 5952 39266 6016
rect 39330 5952 39346 6016
rect 39410 5952 39426 6016
rect 39490 5952 39506 6016
rect 39570 5952 39578 6016
rect 39258 4928 39578 5952
rect 39258 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39578 4928
rect 39258 3840 39578 4864
rect 39258 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39578 3840
rect 39258 2752 39578 3776
rect 39258 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39578 2752
rect 39258 2128 39578 2688
rect 44731 7648 45051 7664
rect 44731 7584 44739 7648
rect 44803 7584 44819 7648
rect 44883 7584 44899 7648
rect 44963 7584 44979 7648
rect 45043 7584 45051 7648
rect 44731 6560 45051 7584
rect 44731 6496 44739 6560
rect 44803 6496 44819 6560
rect 44883 6496 44899 6560
rect 44963 6496 44979 6560
rect 45043 6496 45051 6560
rect 44731 5472 45051 6496
rect 44731 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45051 5472
rect 44731 4384 45051 5408
rect 44731 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45051 4384
rect 44731 3296 45051 4320
rect 44731 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45051 3296
rect 44731 2208 45051 3232
rect 44731 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45051 2208
rect 44731 2128 45051 2144
rect 31891 1188 31957 1189
rect 31891 1124 31892 1188
rect 31956 1124 31957 1188
rect 31891 1123 31957 1124
rect 24899 1052 24965 1053
rect 24899 988 24900 1052
rect 24964 988 24965 1052
rect 24899 987 24965 988
rect 18827 100 18893 101
rect 18827 36 18828 100
rect 18892 36 18893 100
rect 18827 35 18893 36
rect 19011 100 19077 101
rect 19011 36 19012 100
rect 19076 36 19077 100
rect 19011 35 19077 36
use sky130_fd_sc_hd__buf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _01_
timestamp 1688980957
transform 1 0 26312 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _02_
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _03_
timestamp 1688980957
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _05_
timestamp 1688980957
transform 1 0 20792 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _06_
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _07_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 14260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 23736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 24472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 25024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 21160 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1688980957
transform 1 0 25944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 28428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 28336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 28612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _47_
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _48_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform 1 0 24748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _52_
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 31556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1688980957
transform 1 0 31832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1688980957
transform 1 0 32108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1688980957
transform 1 0 27416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1688980957
transform 1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1688980957
transform 1 0 32384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1688980957
transform 1 0 30268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _64_
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _65_
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _66_
timestamp 1688980957
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _67_
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _68_
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1688980957
transform 1 0 33764 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform 1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform 1 0 36800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1688980957
transform 1 0 36340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1688980957
transform 1 0 37076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1688980957
transform 1 0 37812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1688980957
transform 1 0 38548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _77_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _78_
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _79_
timestamp 1688980957
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _80_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _81_
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _82_
timestamp 1688980957
transform 1 0 17940 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _83_
timestamp 1688980957
transform 1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _84_
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _85_
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _86_
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _87_
timestamp 1688980957
transform 1 0 27968 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _88_
timestamp 1688980957
transform 1 0 26312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _89_
timestamp 1688980957
transform 1 0 29624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _90_
timestamp 1688980957
transform 1 0 27048 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _91_
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _92_
timestamp 1688980957
transform 1 0 26680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_179
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_436
timestamp 1688980957
transform 1 0 41216 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_90
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_102 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_133
timestamp 1688980957
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_138
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_147
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_155 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_199
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_376
timestamp 1688980957
transform 1 0 35696 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_388
timestamp 1688980957
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_414
timestamp 1688980957
transform 1 0 39192 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_426
timestamp 1688980957
transform 1 0 40296 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_438
timestamp 1688980957
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_446
timestamp 1688980957
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_192
timestamp 1688980957
transform 1 0 18768 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_212
timestamp 1688980957
transform 1 0 20608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_220
timestamp 1688980957
transform 1 0 21344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_236
timestamp 1688980957
transform 1 0 22816 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_266
timestamp 1688980957
transform 1 0 25576 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_273
timestamp 1688980957
transform 1 0 26220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_320
timestamp 1688980957
transform 1 0 30544 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_343
timestamp 1688980957
transform 1 0 32660 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_351
timestamp 1688980957
transform 1 0 33396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_189
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_198
timestamp 1688980957
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_210
timestamp 1688980957
transform 1 0 20424 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_228
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_240
timestamp 1688980957
transform 1 0 23184 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_252
timestamp 1688980957
transform 1 0 24288 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_264
timestamp 1688980957
transform 1 0 25392 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_272
timestamp 1688980957
transform 1 0 26128 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_344
timestamp 1688980957
transform 1 0 32752 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_356
timestamp 1688980957
transform 1 0 33856 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_368
timestamp 1688980957
transform 1 0 34960 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_380
timestamp 1688980957
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_21
timestamp 1688980957
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_353
timestamp 1688980957
transform 1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_358
timestamp 1688980957
transform 1 0 34040 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_368
timestamp 1688980957
transform 1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_374
timestamp 1688980957
transform 1 0 35512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_382
timestamp 1688980957
transform 1 0 36248 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_386
timestamp 1688980957
transform 1 0 36616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_390
timestamp 1688980957
transform 1 0 36984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_394
timestamp 1688980957
transform 1 0 37352 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_398
timestamp 1688980957
transform 1 0 37720 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_402
timestamp 1688980957
transform 1 0 38088 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_406
timestamp 1688980957
transform 1 0 38456 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_410
timestamp 1688980957
transform 1 0 38824 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_418
timestamp 1688980957
transform 1 0 39560 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_12
timestamp 1688980957
transform 1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_20
timestamp 1688980957
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_29
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_72
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_76
timestamp 1688980957
transform 1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_92
timestamp 1688980957
transform 1 0 9568 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_124
timestamp 1688980957
transform 1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_132
timestamp 1688980957
transform 1 0 13248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_141
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_148
timestamp 1688980957
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_156
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_164
timestamp 1688980957
transform 1 0 16192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_172
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_177
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_185
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_197
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_204
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_212
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_228
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_236
timestamp 1688980957
transform 1 0 22816 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_244
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_260
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_269
timestamp 1688980957
transform 1 0 25852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_276
timestamp 1688980957
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_284
timestamp 1688980957
transform 1 0 27232 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_289
timestamp 1688980957
transform 1 0 27692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_300
timestamp 1688980957
transform 1 0 28704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_309
timestamp 1688980957
transform 1 0 29532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_313
timestamp 1688980957
transform 1 0 29900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_321
timestamp 1688980957
transform 1 0 30636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_325
timestamp 1688980957
transform 1 0 31004 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_332
timestamp 1688980957
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_356
timestamp 1688980957
transform 1 0 33856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_365
timestamp 1688980957
transform 1 0 34684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_372
timestamp 1688980957
transform 1 0 35328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_380
timestamp 1688980957
transform 1 0 36064 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_412
timestamp 1688980957
transform 1 0 39008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_421
timestamp 1688980957
transform 1 0 39836 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_428
timestamp 1688980957
transform 1 0 40480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_436
timestamp 1688980957
transform 1 0 41216 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_444
timestamp 1688980957
transform 1 0 41952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_468
timestamp 1688980957
transform 1 0 44160 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_472
timestamp 1688980957
transform 1 0 44528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 38640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 39468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 38916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 40388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 40664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 36064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 36616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 10304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 19044 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1688980957
transform 1 0 15640 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 17112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform 1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1688980957
transform 1 0 19320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1688980957
transform 1 0 22264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1688980957
transform 1 0 24472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1688980957
transform 1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1688980957
transform 1 0 25944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1688980957
transform 1 0 27416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1688980957
transform 1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1688980957
transform 1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1688980957
transform 1 0 29624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output90 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 9016 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 9752 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 11960 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 12696 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 13432 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 14168 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 14904 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 15640 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 2392 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 3864 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 4600 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform -1 0 8832 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 24932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 24564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 22080 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 22080 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform 1 0 30084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 27508 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 28612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 31188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output147
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output148
timestamp 1688980957
transform 1 0 33764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output149
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output150
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output151
timestamp 1688980957
transform 1 0 35236 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output152
timestamp 1688980957
transform 1 0 34868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output153
timestamp 1688980957
transform 1 0 30820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output154
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output155
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output156
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output157
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output158
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output159
timestamp 1688980957
transform 1 0 32660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output160
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output161
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output162
timestamp 1688980957
transform 1 0 31096 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output163
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output164
timestamp 1688980957
transform 1 0 32660 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output165
timestamp 1688980957
transform 1 0 33304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output166
timestamp 1688980957
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output167
timestamp 1688980957
transform 1 0 34776 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output168
timestamp 1688980957
transform 1 0 35512 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output169
timestamp 1688980957
transform 1 0 36248 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output170
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output171
timestamp 1688980957
transform 1 0 37812 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output172
timestamp 1688980957
transform 1 0 38456 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output173
timestamp 1688980957
transform 1 0 39192 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output174
timestamp 1688980957
transform 1 0 39928 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output175
timestamp 1688980957
transform 1 0 40664 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output176
timestamp 1688980957
transform 1 0 41400 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output177
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output178
timestamp 1688980957
transform 1 0 42964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output179
timestamp 1688980957
transform 1 0 43608 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output180
timestamp 1688980957
transform 1 0 44068 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output181
timestamp 1688980957
transform 1 0 43516 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output182
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 44896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 44896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 44896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 44896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 34702 0 34758 160 0 FreeSans 224 90 0 0 Ci
port 0 nsew signal input
flabel metal2 s 34978 0 35034 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 1 nsew signal input
flabel metal2 s 37738 0 37794 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 2 nsew signal input
flabel metal2 s 38014 0 38070 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 3 nsew signal input
flabel metal2 s 38290 0 38346 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 4 nsew signal input
flabel metal2 s 38566 0 38622 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 5 nsew signal input
flabel metal2 s 38842 0 38898 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 6 nsew signal input
flabel metal2 s 39118 0 39174 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 7 nsew signal input
flabel metal2 s 39394 0 39450 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 8 nsew signal input
flabel metal2 s 39670 0 39726 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 9 nsew signal input
flabel metal2 s 39946 0 40002 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 10 nsew signal input
flabel metal2 s 40222 0 40278 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 11 nsew signal input
flabel metal2 s 35254 0 35310 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 12 nsew signal input
flabel metal2 s 35530 0 35586 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 13 nsew signal input
flabel metal2 s 35806 0 35862 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 14 nsew signal input
flabel metal2 s 36082 0 36138 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 15 nsew signal input
flabel metal2 s 36358 0 36414 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 16 nsew signal input
flabel metal2 s 36634 0 36690 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 17 nsew signal input
flabel metal2 s 36910 0 36966 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 18 nsew signal input
flabel metal2 s 37186 0 37242 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 19 nsew signal input
flabel metal2 s 37462 0 37518 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 20 nsew signal input
flabel metal2 s 1582 9840 1638 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 21 nsew signal tristate
flabel metal2 s 8942 9840 8998 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 22 nsew signal tristate
flabel metal2 s 9678 9840 9734 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 23 nsew signal tristate
flabel metal2 s 10414 9840 10470 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 24 nsew signal tristate
flabel metal2 s 11150 9840 11206 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 25 nsew signal tristate
flabel metal2 s 11886 9840 11942 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 26 nsew signal tristate
flabel metal2 s 12622 9840 12678 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 27 nsew signal tristate
flabel metal2 s 13358 9840 13414 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 28 nsew signal tristate
flabel metal2 s 14094 9840 14150 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 29 nsew signal tristate
flabel metal2 s 14830 9840 14886 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 30 nsew signal tristate
flabel metal2 s 15566 9840 15622 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 31 nsew signal tristate
flabel metal2 s 2318 9840 2374 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 32 nsew signal tristate
flabel metal2 s 3054 9840 3110 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 33 nsew signal tristate
flabel metal2 s 3790 9840 3846 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 34 nsew signal tristate
flabel metal2 s 4526 9840 4582 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 35 nsew signal tristate
flabel metal2 s 5262 9840 5318 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 36 nsew signal tristate
flabel metal2 s 5998 9840 6054 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 37 nsew signal tristate
flabel metal2 s 6734 9840 6790 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 38 nsew signal tristate
flabel metal2 s 7470 9840 7526 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 39 nsew signal tristate
flabel metal2 s 8206 9840 8262 10000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 40 nsew signal tristate
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N1END[0]
port 41 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N1END[1]
port 42 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N1END[2]
port 43 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N1END[3]
port 44 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N2END[0]
port 45 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N2END[1]
port 46 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N2END[2]
port 47 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N2END[3]
port 48 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 N2END[4]
port 49 nsew signal input
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 N2END[5]
port 50 nsew signal input
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 N2END[6]
port 51 nsew signal input
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 N2END[7]
port 52 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N2MID[0]
port 53 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N2MID[1]
port 54 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N2MID[2]
port 55 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N2MID[3]
port 56 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N2MID[4]
port 57 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N2MID[5]
port 58 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N2MID[6]
port 59 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N2MID[7]
port 60 nsew signal input
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 N4END[0]
port 61 nsew signal input
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 N4END[10]
port 62 nsew signal input
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 N4END[11]
port 63 nsew signal input
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 N4END[12]
port 64 nsew signal input
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 N4END[13]
port 65 nsew signal input
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 N4END[14]
port 66 nsew signal input
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 N4END[15]
port 67 nsew signal input
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 N4END[1]
port 68 nsew signal input
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 N4END[2]
port 69 nsew signal input
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 N4END[3]
port 70 nsew signal input
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 N4END[4]
port 71 nsew signal input
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 N4END[5]
port 72 nsew signal input
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 N4END[6]
port 73 nsew signal input
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 N4END[7]
port 74 nsew signal input
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 N4END[8]
port 75 nsew signal input
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 N4END[9]
port 76 nsew signal input
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 NN4END[0]
port 77 nsew signal input
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 NN4END[10]
port 78 nsew signal input
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 NN4END[11]
port 79 nsew signal input
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 NN4END[12]
port 80 nsew signal input
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 NN4END[13]
port 81 nsew signal input
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 NN4END[14]
port 82 nsew signal input
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 NN4END[15]
port 83 nsew signal input
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 NN4END[1]
port 84 nsew signal input
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 NN4END[2]
port 85 nsew signal input
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 NN4END[3]
port 86 nsew signal input
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 NN4END[4]
port 87 nsew signal input
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 NN4END[5]
port 88 nsew signal input
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 NN4END[6]
port 89 nsew signal input
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 NN4END[7]
port 90 nsew signal input
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 NN4END[8]
port 91 nsew signal input
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 NN4END[9]
port 92 nsew signal input
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 93 nsew signal tristate
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 94 nsew signal tristate
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 95 nsew signal tristate
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 96 nsew signal tristate
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 97 nsew signal tristate
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 98 nsew signal tristate
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 99 nsew signal tristate
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 100 nsew signal tristate
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 101 nsew signal tristate
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 102 nsew signal tristate
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 103 nsew signal tristate
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 104 nsew signal tristate
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 105 nsew signal tristate
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 106 nsew signal tristate
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 107 nsew signal tristate
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 108 nsew signal tristate
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 109 nsew signal tristate
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 110 nsew signal tristate
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 111 nsew signal tristate
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 112 nsew signal tristate
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 113 nsew signal tristate
flabel metal2 s 28354 0 28410 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 114 nsew signal tristate
flabel metal2 s 28630 0 28686 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 115 nsew signal tristate
flabel metal2 s 28906 0 28962 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 116 nsew signal tristate
flabel metal2 s 29182 0 29238 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 117 nsew signal tristate
flabel metal2 s 29458 0 29514 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 118 nsew signal tristate
flabel metal2 s 29734 0 29790 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 119 nsew signal tristate
flabel metal2 s 25870 0 25926 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 120 nsew signal tristate
flabel metal2 s 26146 0 26202 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 121 nsew signal tristate
flabel metal2 s 26422 0 26478 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 122 nsew signal tristate
flabel metal2 s 26698 0 26754 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 123 nsew signal tristate
flabel metal2 s 26974 0 27030 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 124 nsew signal tristate
flabel metal2 s 27250 0 27306 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 125 nsew signal tristate
flabel metal2 s 27526 0 27582 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 126 nsew signal tristate
flabel metal2 s 27802 0 27858 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 127 nsew signal tristate
flabel metal2 s 28078 0 28134 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 128 nsew signal tristate
flabel metal2 s 30010 0 30066 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 129 nsew signal tristate
flabel metal2 s 32770 0 32826 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 130 nsew signal tristate
flabel metal2 s 33046 0 33102 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 131 nsew signal tristate
flabel metal2 s 33322 0 33378 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 132 nsew signal tristate
flabel metal2 s 33598 0 33654 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 133 nsew signal tristate
flabel metal2 s 33874 0 33930 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 134 nsew signal tristate
flabel metal2 s 34150 0 34206 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 135 nsew signal tristate
flabel metal2 s 30286 0 30342 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 136 nsew signal tristate
flabel metal2 s 30562 0 30618 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 137 nsew signal tristate
flabel metal2 s 30838 0 30894 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 138 nsew signal tristate
flabel metal2 s 31114 0 31170 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 139 nsew signal tristate
flabel metal2 s 31390 0 31446 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 140 nsew signal tristate
flabel metal2 s 31666 0 31722 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 141 nsew signal tristate
flabel metal2 s 31942 0 31998 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 142 nsew signal tristate
flabel metal2 s 32218 0 32274 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 143 nsew signal tristate
flabel metal2 s 32494 0 32550 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 144 nsew signal tristate
flabel metal2 s 16302 9840 16358 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN0
port 145 nsew signal input
flabel metal2 s 17038 9840 17094 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN1
port 146 nsew signal input
flabel metal2 s 17774 9840 17830 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN10
port 147 nsew signal input
flabel metal2 s 18510 9840 18566 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN11
port 148 nsew signal input
flabel metal2 s 19246 9840 19302 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN12
port 149 nsew signal input
flabel metal2 s 19982 9840 20038 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN13
port 150 nsew signal input
flabel metal2 s 20718 9840 20774 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN14
port 151 nsew signal input
flabel metal2 s 21454 9840 21510 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN15
port 152 nsew signal input
flabel metal2 s 22190 9840 22246 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN16
port 153 nsew signal input
flabel metal2 s 22926 9840 22982 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN17
port 154 nsew signal input
flabel metal2 s 23662 9840 23718 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN18
port 155 nsew signal input
flabel metal2 s 24398 9840 24454 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN19
port 156 nsew signal input
flabel metal2 s 25134 9840 25190 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN2
port 157 nsew signal input
flabel metal2 s 25870 9840 25926 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN3
port 158 nsew signal input
flabel metal2 s 26606 9840 26662 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN4
port 159 nsew signal input
flabel metal2 s 27342 9840 27398 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN5
port 160 nsew signal input
flabel metal2 s 28078 9840 28134 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN6
port 161 nsew signal input
flabel metal2 s 28814 9840 28870 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN7
port 162 nsew signal input
flabel metal2 s 29550 9840 29606 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN8
port 163 nsew signal input
flabel metal2 s 30286 9840 30342 10000 0 FreeSans 224 90 0 0 UIO_TOP_UIN9
port 164 nsew signal input
flabel metal2 s 31022 9840 31078 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT0
port 165 nsew signal tristate
flabel metal2 s 31758 9840 31814 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT1
port 166 nsew signal tristate
flabel metal2 s 32494 9840 32550 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT10
port 167 nsew signal tristate
flabel metal2 s 33230 9840 33286 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT11
port 168 nsew signal tristate
flabel metal2 s 33966 9840 34022 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT12
port 169 nsew signal tristate
flabel metal2 s 34702 9840 34758 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT13
port 170 nsew signal tristate
flabel metal2 s 35438 9840 35494 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT14
port 171 nsew signal tristate
flabel metal2 s 36174 9840 36230 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT15
port 172 nsew signal tristate
flabel metal2 s 36910 9840 36966 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT16
port 173 nsew signal tristate
flabel metal2 s 37646 9840 37702 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT17
port 174 nsew signal tristate
flabel metal2 s 38382 9840 38438 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT18
port 175 nsew signal tristate
flabel metal2 s 39118 9840 39174 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT19
port 176 nsew signal tristate
flabel metal2 s 39854 9840 39910 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT2
port 177 nsew signal tristate
flabel metal2 s 40590 9840 40646 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT3
port 178 nsew signal tristate
flabel metal2 s 41326 9840 41382 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT4
port 179 nsew signal tristate
flabel metal2 s 42062 9840 42118 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT5
port 180 nsew signal tristate
flabel metal2 s 42798 9840 42854 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT6
port 181 nsew signal tristate
flabel metal2 s 43534 9840 43590 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT7
port 182 nsew signal tristate
flabel metal2 s 44270 9840 44326 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT8
port 183 nsew signal tristate
flabel metal2 s 45006 9840 45062 10000 0 FreeSans 224 90 0 0 UIO_TOP_UOUT9
port 184 nsew signal tristate
flabel metal2 s 34426 0 34482 160 0 FreeSans 224 90 0 0 UserCLK
port 185 nsew signal input
flabel metal2 s 846 9840 902 10000 0 FreeSans 224 90 0 0 UserCLKo
port 186 nsew signal tristate
flabel metal4 s 6417 2128 6737 7664 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 17364 2128 17684 7664 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 28311 2128 28631 7664 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 39258 2128 39578 7664 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 11890 2128 12210 7664 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
flabel metal4 s 22837 2128 23157 7664 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
flabel metal4 s 33784 2128 34104 7664 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
flabel metal4 s 44731 2128 45051 7664 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
rlabel metal1 23000 7072 23000 7072 0 vccd1
rlabel via1 23077 7616 23077 7616 0 vssd1
rlabel metal2 35059 68 35059 68 0 FrameStrobe[0]
rlabel metal2 37865 68 37865 68 0 FrameStrobe[10]
rlabel metal2 38141 68 38141 68 0 FrameStrobe[11]
rlabel metal2 38417 68 38417 68 0 FrameStrobe[12]
rlabel metal2 38594 755 38594 755 0 FrameStrobe[13]
rlabel metal2 38923 68 38923 68 0 FrameStrobe[14]
rlabel metal2 39146 1214 39146 1214 0 FrameStrobe[15]
rlabel metal2 39422 1282 39422 1282 0 FrameStrobe[16]
rlabel metal2 39797 68 39797 68 0 FrameStrobe[17]
rlabel metal2 39974 1282 39974 1282 0 FrameStrobe[18]
rlabel metal2 40250 1214 40250 1214 0 FrameStrobe[19]
rlabel metal2 35282 1282 35282 1282 0 FrameStrobe[1]
rlabel metal2 35657 68 35657 68 0 FrameStrobe[2]
rlabel metal2 35834 755 35834 755 0 FrameStrobe[3]
rlabel metal2 36110 1180 36110 1180 0 FrameStrobe[4]
rlabel metal2 36386 1282 36386 1282 0 FrameStrobe[5]
rlabel metal2 36662 1180 36662 1180 0 FrameStrobe[6]
rlabel metal2 36938 1299 36938 1299 0 FrameStrobe[7]
rlabel metal2 37214 1214 37214 1214 0 FrameStrobe[8]
rlabel metal2 37589 68 37589 68 0 FrameStrobe[9]
rlabel metal2 1610 8680 1610 8680 0 FrameStrobe_O[0]
rlabel metal2 8970 8680 8970 8680 0 FrameStrobe_O[10]
rlabel metal2 9706 8680 9706 8680 0 FrameStrobe_O[11]
rlabel metal2 10442 8680 10442 8680 0 FrameStrobe_O[12]
rlabel metal2 11178 8680 11178 8680 0 FrameStrobe_O[13]
rlabel metal2 11914 9173 11914 9173 0 FrameStrobe_O[14]
rlabel metal2 12650 8680 12650 8680 0 FrameStrobe_O[15]
rlabel metal2 13386 9785 13386 9785 0 FrameStrobe_O[16]
rlabel metal2 14122 8680 14122 8680 0 FrameStrobe_O[17]
rlabel metal2 14858 9173 14858 9173 0 FrameStrobe_O[18]
rlabel metal2 15594 8680 15594 8680 0 FrameStrobe_O[19]
rlabel metal2 2346 9785 2346 9785 0 FrameStrobe_O[1]
rlabel metal2 3082 8680 3082 8680 0 FrameStrobe_O[2]
rlabel metal2 3818 9173 3818 9173 0 FrameStrobe_O[3]
rlabel metal2 4554 8680 4554 8680 0 FrameStrobe_O[4]
rlabel metal2 5290 9037 5290 9037 0 FrameStrobe_O[5]
rlabel metal2 6026 9173 6026 9173 0 FrameStrobe_O[6]
rlabel metal2 6762 9241 6762 9241 0 FrameStrobe_O[7]
rlabel metal2 7498 8680 7498 8680 0 FrameStrobe_O[8]
rlabel metal2 8234 9037 8234 9037 0 FrameStrobe_O[9]
rlabel metal2 5750 1248 5750 1248 0 N1END[0]
rlabel metal2 6026 1248 6026 1248 0 N1END[1]
rlabel metal2 6302 1248 6302 1248 0 N1END[2]
rlabel metal2 6479 68 6479 68 0 N1END[3]
rlabel metal2 9115 68 9115 68 0 N2END[0]
rlabel metal2 9338 1214 9338 1214 0 N2END[1]
rlabel metal2 9515 68 9515 68 0 N2END[2]
rlabel metal2 9791 68 9791 68 0 N2END[3]
rlabel metal2 10166 1214 10166 1214 0 N2END[4]
rlabel metal2 10442 1248 10442 1248 0 N2END[5]
rlabel metal2 10619 68 10619 68 0 N2END[6]
rlabel metal2 10895 68 10895 68 0 N2END[7]
rlabel metal2 6755 68 6755 68 0 N2MID[0]
rlabel metal2 7031 68 7031 68 0 N2MID[1]
rlabel metal2 7307 68 7307 68 0 N2MID[2]
rlabel metal2 7583 68 7583 68 0 N2MID[3]
rlabel metal2 7859 68 7859 68 0 N2MID[4]
rlabel metal2 8135 68 8135 68 0 N2MID[5]
rlabel metal2 8411 68 8411 68 0 N2MID[6]
rlabel metal2 8687 68 8687 68 0 N2MID[7]
rlabel metal2 11171 68 11171 68 0 N4END[0]
rlabel metal2 13931 68 13931 68 0 N4END[10]
rlabel metal2 14359 68 14359 68 0 N4END[11]
rlabel metal2 11546 687 11546 687 0 N4END[1]
rlabel metal2 11822 1248 11822 1248 0 N4END[2]
rlabel metal2 12098 687 12098 687 0 N4END[3]
rlabel metal2 12374 1299 12374 1299 0 N4END[4]
rlabel metal2 12650 1248 12650 1248 0 N4END[5]
rlabel metal2 12926 1248 12926 1248 0 N4END[6]
rlabel metal2 13202 1248 13202 1248 0 N4END[7]
rlabel metal2 13478 1421 13478 1421 0 N4END[8]
rlabel metal2 13754 687 13754 687 0 N4END[9]
rlabel metal2 15686 1520 15686 1520 0 NN4END[0]
rlabel metal2 18446 1299 18446 1299 0 NN4END[10]
rlabel metal2 18775 68 18775 68 0 NN4END[11]
rlabel metal2 18998 143 18998 143 0 NN4END[12]
rlabel metal2 19274 1095 19274 1095 0 NN4END[13]
rlabel metal2 19497 68 19497 68 0 NN4END[14]
rlabel metal2 19826 687 19826 687 0 NN4END[15]
rlabel metal2 15909 68 15909 68 0 NN4END[1]
rlabel metal2 16337 68 16337 68 0 NN4END[2]
rlabel metal1 16560 3502 16560 3502 0 NN4END[3]
rlabel metal2 16790 1421 16790 1421 0 NN4END[4]
rlabel metal2 17066 1214 17066 1214 0 NN4END[5]
rlabel metal2 17342 823 17342 823 0 NN4END[6]
rlabel metal2 17717 68 17717 68 0 NN4END[7]
rlabel metal1 17894 3400 17894 3400 0 NN4END[8]
rlabel metal1 17848 3026 17848 3026 0 NN4END[9]
rlabel metal2 20194 2788 20194 2788 0 S1BEG[0]
rlabel metal2 20378 1282 20378 1282 0 S1BEG[1]
rlabel metal1 20746 2822 20746 2822 0 S1BEG[2]
rlabel metal2 20831 68 20831 68 0 S1BEG[3]
rlabel metal2 23414 1180 23414 1180 0 S2BEG[0]
rlabel metal2 23690 1180 23690 1180 0 S2BEG[1]
rlabel metal2 23966 1180 23966 1180 0 S2BEG[2]
rlabel metal2 24341 68 24341 68 0 S2BEG[3]
rlabel metal1 24656 2822 24656 2822 0 S2BEG[4]
rlabel metal2 24794 1180 24794 1180 0 S2BEG[5]
rlabel metal1 25208 2822 25208 2822 0 S2BEG[6]
rlabel metal2 25445 68 25445 68 0 S2BEG[7]
rlabel metal2 21305 68 21305 68 0 S2BEGb[0]
rlabel metal2 21482 1214 21482 1214 0 S2BEGb[1]
rlabel metal2 21705 68 21705 68 0 S2BEGb[2]
rlabel metal2 22034 1452 22034 1452 0 S2BEGb[3]
rlabel metal2 22363 68 22363 68 0 S2BEGb[4]
rlabel metal1 22724 2822 22724 2822 0 S2BEGb[5]
rlabel metal2 22809 68 22809 68 0 S2BEGb[6]
rlabel metal2 23237 68 23237 68 0 S2BEGb[7]
rlabel metal1 25760 2822 25760 2822 0 S4BEG[0]
rlabel metal2 28481 68 28481 68 0 S4BEG[10]
rlabel metal2 28757 68 28757 68 0 S4BEG[11]
rlabel metal2 28934 1316 28934 1316 0 S4BEG[12]
rlabel metal1 29578 2890 29578 2890 0 S4BEG[13]
rlabel metal2 29539 68 29539 68 0 S4BEG[14]
rlabel metal1 30130 3162 30130 3162 0 S4BEG[15]
rlabel metal2 25997 68 25997 68 0 S4BEG[1]
rlabel metal2 26174 1214 26174 1214 0 S4BEG[2]
rlabel metal2 26542 2822 26542 2822 0 S4BEG[3]
rlabel metal2 26825 68 26825 68 0 S4BEG[4]
rlabel metal1 27370 2890 27370 2890 0 S4BEG[5]
rlabel metal2 27377 68 27377 68 0 S4BEG[6]
rlabel metal1 27922 3162 27922 3162 0 S4BEG[7]
rlabel metal2 27929 68 27929 68 0 S4BEG[8]
rlabel metal2 28159 68 28159 68 0 S4BEG[9]
rlabel metal2 30091 68 30091 68 0 SS4BEG[0]
rlabel metal1 32936 3706 32936 3706 0 SS4BEG[10]
rlabel metal1 33534 2890 33534 2890 0 SS4BEG[11]
rlabel metal2 33449 68 33449 68 0 SS4BEG[12]
rlabel metal1 34086 3162 34086 3162 0 SS4BEG[13]
rlabel metal2 34001 68 34001 68 0 SS4BEG[14]
rlabel metal1 34638 2822 34638 2822 0 SS4BEG[15]
rlabel metal2 30261 68 30261 68 0 SS4BEG[1]
rlabel metal1 31096 2890 31096 2890 0 SS4BEG[2]
rlabel metal2 30965 68 30965 68 0 SS4BEG[3]
rlabel metal1 32154 2380 32154 2380 0 SS4BEG[4]
rlabel metal2 31517 68 31517 68 0 SS4BEG[5]
rlabel metal2 31694 1282 31694 1282 0 SS4BEG[6]
rlabel metal2 31970 687 31970 687 0 SS4BEG[7]
rlabel metal2 32345 68 32345 68 0 SS4BEG[8]
rlabel metal1 32982 2822 32982 2822 0 SS4BEG[9]
rlabel metal2 16330 8612 16330 8612 0 UIO_TOP_UIN0
rlabel metal2 17066 8612 17066 8612 0 UIO_TOP_UIN1
rlabel metal2 17802 8612 17802 8612 0 UIO_TOP_UIN10
rlabel metal2 18538 8612 18538 8612 0 UIO_TOP_UIN11
rlabel metal1 19274 7446 19274 7446 0 UIO_TOP_UIN12
rlabel metal2 20010 8612 20010 8612 0 UIO_TOP_UIN13
rlabel metal2 20746 8612 20746 8612 0 UIO_TOP_UIN14
rlabel metal2 21482 8612 21482 8612 0 UIO_TOP_UIN15
rlabel metal2 22218 8612 22218 8612 0 UIO_TOP_UIN16
rlabel metal2 22954 9785 22954 9785 0 UIO_TOP_UIN17
rlabel metal2 23690 8612 23690 8612 0 UIO_TOP_UIN18
rlabel metal2 24426 8612 24426 8612 0 UIO_TOP_UIN19
rlabel metal2 25162 8612 25162 8612 0 UIO_TOP_UIN2
rlabel metal2 25898 8612 25898 8612 0 UIO_TOP_UIN3
rlabel metal2 26634 8612 26634 8612 0 UIO_TOP_UIN4
rlabel metal2 27370 8612 27370 8612 0 UIO_TOP_UIN5
rlabel metal2 28106 8612 28106 8612 0 UIO_TOP_UIN6
rlabel metal2 28842 9037 28842 9037 0 UIO_TOP_UIN7
rlabel metal2 29578 8612 29578 8612 0 UIO_TOP_UIN8
rlabel metal2 30314 8561 30314 8561 0 UIO_TOP_UIN9
rlabel metal2 31050 8680 31050 8680 0 UIO_TOP_UOUT0
rlabel metal2 31786 8680 31786 8680 0 UIO_TOP_UOUT1
rlabel metal2 32522 8680 32522 8680 0 UIO_TOP_UOUT10
rlabel metal2 33258 8680 33258 8680 0 UIO_TOP_UOUT11
rlabel metal2 33994 9785 33994 9785 0 UIO_TOP_UOUT12
rlabel metal2 34730 8680 34730 8680 0 UIO_TOP_UOUT13
rlabel metal2 35466 9785 35466 9785 0 UIO_TOP_UOUT14
rlabel metal2 36202 8680 36202 8680 0 UIO_TOP_UOUT15
rlabel metal2 36938 9785 36938 9785 0 UIO_TOP_UOUT16
rlabel metal2 37674 8680 37674 8680 0 UIO_TOP_UOUT17
rlabel metal2 38410 8680 38410 8680 0 UIO_TOP_UOUT18
rlabel metal2 39146 8680 39146 8680 0 UIO_TOP_UOUT19
rlabel metal2 39882 8680 39882 8680 0 UIO_TOP_UOUT2
rlabel metal2 40618 8680 40618 8680 0 UIO_TOP_UOUT3
rlabel metal2 41354 8680 41354 8680 0 UIO_TOP_UOUT4
rlabel metal2 42090 9785 42090 9785 0 UIO_TOP_UOUT5
rlabel metal2 42826 8680 42826 8680 0 UIO_TOP_UOUT6
rlabel metal2 43562 8680 43562 8680 0 UIO_TOP_UOUT7
rlabel metal2 44298 8408 44298 8408 0 UIO_TOP_UOUT8
rlabel metal1 44528 6834 44528 6834 0 UIO_TOP_UOUT9
rlabel metal2 34401 68 34401 68 0 UserCLK
rlabel metal1 1334 6834 1334 6834 0 UserCLKo
rlabel metal2 35466 3366 35466 3366 0 net1
rlabel metal2 14766 1870 14766 1870 0 net10
rlabel metal1 14858 2312 14858 2312 0 net100
rlabel metal1 2852 7378 2852 7378 0 net101
rlabel metal1 5014 7344 5014 7344 0 net102
rlabel metal1 4324 7378 4324 7378 0 net103
rlabel metal1 4738 7276 4738 7276 0 net104
rlabel metal1 8234 7412 8234 7412 0 net105
rlabel metal1 5842 7344 5842 7344 0 net106
rlabel metal2 6808 7378 6808 7378 0 net107
rlabel metal2 7314 6086 7314 6086 0 net108
rlabel metal1 8372 7514 8372 7514 0 net109
rlabel metal2 15134 1751 15134 1751 0 net11
rlabel metal1 20194 3128 20194 3128 0 net110
rlabel metal1 19734 2414 19734 2414 0 net111
rlabel via2 18354 2635 18354 2635 0 net112
rlabel metal1 19412 2346 19412 2346 0 net113
rlabel metal2 21850 2652 21850 2652 0 net114
rlabel metal1 23736 2414 23736 2414 0 net115
rlabel metal1 21850 2312 21850 2312 0 net116
rlabel metal1 24978 2414 24978 2414 0 net117
rlabel metal1 24702 2992 24702 2992 0 net118
rlabel metal1 25530 2414 25530 2414 0 net119
rlabel metal1 36018 2618 36018 2618 0 net12
rlabel metal1 24886 3094 24886 3094 0 net120
rlabel metal1 25714 2346 25714 2346 0 net121
rlabel metal1 19458 2618 19458 2618 0 net122
rlabel metal1 20746 2312 20746 2312 0 net123
rlabel metal1 21252 2414 21252 2414 0 net124
rlabel metal1 21482 3060 21482 3060 0 net125
rlabel metal1 22172 2414 22172 2414 0 net126
rlabel metal2 21758 3264 21758 3264 0 net127
rlabel metal2 21988 3366 21988 3366 0 net128
rlabel metal1 23322 3128 23322 3128 0 net129
rlabel metal2 36570 2329 36570 2329 0 net13
rlabel metal1 25576 3094 25576 3094 0 net130
rlabel metal1 29578 2414 29578 2414 0 net131
rlabel metal1 29164 3026 29164 3026 0 net132
rlabel metal1 29670 2346 29670 2346 0 net133
rlabel metal1 29532 3094 29532 3094 0 net134
rlabel metal2 17250 3706 17250 3706 0 net135
rlabel metal2 19366 6647 19366 6647 0 net136
rlabel metal1 21114 3400 21114 3400 0 net137
rlabel metal2 21022 2349 21022 2349 0 net138
rlabel metal1 27094 3128 27094 3128 0 net139
rlabel metal3 32844 3400 32844 3400 0 net14
rlabel metal1 27784 2414 27784 2414 0 net140
rlabel metal1 27416 3094 27416 3094 0 net141
rlabel metal1 30958 2482 30958 2482 0 net142
rlabel metal1 28198 2992 28198 2992 0 net143
rlabel metal2 28796 3604 28796 3604 0 net144
rlabel metal1 28520 3026 28520 3026 0 net145
rlabel metal1 30866 2346 30866 2346 0 net146
rlabel metal1 33672 2550 33672 2550 0 net147
rlabel metal1 33672 3026 33672 3026 0 net148
rlabel metal2 34822 2210 34822 2210 0 net149
rlabel metal2 37122 3111 37122 3111 0 net15
rlabel metal1 33672 3094 33672 3094 0 net150
rlabel metal1 35374 2040 35374 2040 0 net151
rlabel metal1 34684 3026 34684 3026 0 net152
rlabel metal1 30866 3026 30866 3026 0 net153
rlabel metal1 31280 3026 31280 3026 0 net154
rlabel metal2 32246 1955 32246 1955 0 net155
rlabel metal1 32752 2414 32752 2414 0 net156
rlabel metal1 31993 3094 31993 3094 0 net157
rlabel metal1 33258 2414 33258 2414 0 net158
rlabel metal1 32798 3128 32798 3128 0 net159
rlabel metal2 25070 6596 25070 6596 0 net16
rlabel metal1 33488 2346 33488 2346 0 net160
rlabel metal1 33350 2992 33350 2992 0 net161
rlabel metal2 20286 5831 20286 5831 0 net162
rlabel metal1 20562 7310 20562 7310 0 net163
rlabel metal1 17618 3434 17618 3434 0 net164
rlabel metal1 17618 3638 17618 3638 0 net165
rlabel metal1 33994 6970 33994 6970 0 net166
rlabel metal1 34822 6970 34822 6970 0 net167
rlabel metal1 35466 6970 35466 6970 0 net168
rlabel metal1 36616 7446 36616 7446 0 net169
rlabel metal2 37766 1989 37766 1989 0 net17
rlabel metal1 36892 6630 36892 6630 0 net170
rlabel metal1 37306 6970 37306 6970 0 net171
rlabel metal1 38042 6970 38042 6970 0 net172
rlabel metal1 38778 6970 38778 6970 0 net173
rlabel metal1 19826 2958 19826 2958 0 net174
rlabel metal2 19826 7650 19826 7650 0 net175
rlabel metal1 19504 2958 19504 2958 0 net176
rlabel metal2 29302 7514 29302 7514 0 net177
rlabel metal1 31740 7990 31740 7990 0 net178
rlabel metal2 18170 4131 18170 4131 0 net179
rlabel metal1 37950 2618 37950 2618 0 net18
rlabel metal1 17572 2822 17572 2822 0 net180
rlabel metal1 18032 2482 18032 2482 0 net181
rlabel metal2 17250 7276 17250 7276 0 net182
rlabel via2 38134 2533 38134 2533 0 net19
rlabel metal1 39054 1972 39054 1972 0 net2
rlabel metal2 26634 2040 26634 2040 0 net20
rlabel metal2 5658 1972 5658 1972 0 net21
rlabel metal1 6394 2550 6394 2550 0 net22
rlabel metal1 6854 2414 6854 2414 0 net23
rlabel metal1 6670 2618 6670 2618 0 net24
rlabel metal1 22494 2958 22494 2958 0 net25
rlabel metal1 9200 2278 9200 2278 0 net26
rlabel metal1 9476 2278 9476 2278 0 net27
rlabel metal2 9706 3366 9706 3366 0 net28
rlabel metal2 9982 2567 9982 2567 0 net29
rlabel metal1 39100 2618 39100 2618 0 net3
rlabel metal1 10258 2312 10258 2312 0 net30
rlabel metal2 19366 2329 19366 2329 0 net31
rlabel metal1 18722 1496 18722 1496 0 net32
rlabel metal2 7130 1649 7130 1649 0 net33
rlabel metal2 10258 2125 10258 2125 0 net34
rlabel metal2 7406 1972 7406 1972 0 net35
rlabel metal1 7682 2312 7682 2312 0 net36
rlabel metal2 7958 3417 7958 3417 0 net37
rlabel metal2 21574 1802 21574 1802 0 net38
rlabel metal1 8510 2346 8510 2346 0 net39
rlabel metal1 39330 1870 39330 1870 0 net4
rlabel metal1 8786 2346 8786 2346 0 net40
rlabel metal1 21390 3570 21390 3570 0 net41
rlabel metal2 14214 2125 14214 2125 0 net42
rlabel metal2 14582 3655 14582 3655 0 net43
rlabel metal2 11362 3281 11362 3281 0 net44
rlabel metal2 15226 1377 15226 1377 0 net45
rlabel metal1 27278 2006 27278 2006 0 net46
rlabel metal2 19182 1615 19182 1615 0 net47
rlabel metal2 12558 2006 12558 2006 0 net48
rlabel metal1 12834 2312 12834 2312 0 net49
rlabel metal2 39698 1904 39698 1904 0 net5
rlabel metal2 13110 2057 13110 2057 0 net50
rlabel metal2 13754 3876 13754 3876 0 net51
rlabel metal2 31786 3145 31786 3145 0 net52
rlabel metal2 16882 4624 16882 4624 0 net53
rlabel metal1 18814 3128 18814 3128 0 net54
rlabel metal1 19090 3026 19090 3026 0 net55
rlabel metal2 19090 5644 19090 5644 0 net56
rlabel metal1 19320 3094 19320 3094 0 net57
rlabel metal1 19550 3706 19550 3706 0 net58
rlabel metal2 18078 2074 18078 2074 0 net59
rlabel metal2 39146 3978 39146 3978 0 net6
rlabel metal2 15962 4658 15962 4658 0 net60
rlabel metal1 16928 2482 16928 2482 0 net61
rlabel metal2 16790 3808 16790 3808 0 net62
rlabel metal1 17158 3536 17158 3536 0 net63
rlabel metal1 16192 2618 16192 2618 0 net64
rlabel metal1 17480 2414 17480 2414 0 net65
rlabel via1 17711 3094 17711 3094 0 net66
rlabel metal1 18032 3094 18032 3094 0 net67
rlabel metal1 18446 2992 18446 2992 0 net68
rlabel metal1 16698 7412 16698 7412 0 net69
rlabel metal1 15318 2040 15318 2040 0 net7
rlabel metal1 17112 3026 17112 3026 0 net70
rlabel metal2 18078 6749 18078 6749 0 net71
rlabel metal1 26450 7412 26450 7412 0 net72
rlabel metal1 21574 3638 21574 3638 0 net73
rlabel metal1 20470 3502 20470 3502 0 net74
rlabel metal1 21206 3502 21206 3502 0 net75
rlabel metal1 21965 7242 21965 7242 0 net76
rlabel metal1 22586 3570 22586 3570 0 net77
rlabel metal1 23506 3536 23506 3536 0 net78
rlabel metal1 24242 3060 24242 3060 0 net79
rlabel metal1 16560 1632 16560 1632 0 net8
rlabel metal1 24932 3502 24932 3502 0 net80
rlabel metal1 29302 3502 29302 3502 0 net81
rlabel metal1 29072 3502 29072 3502 0 net82
rlabel metal1 28842 3468 28842 3468 0 net83
rlabel metal1 28428 3502 28428 3502 0 net84
rlabel metal1 27876 3502 27876 3502 0 net85
rlabel metal1 28796 7378 28796 7378 0 net86
rlabel metal1 29946 3502 29946 3502 0 net87
rlabel metal2 31970 4794 31970 4794 0 net88
rlabel metal1 35236 2550 35236 2550 0 net89
rlabel metal1 16560 1836 16560 1836 0 net9
rlabel via2 1794 7395 1794 7395 0 net90
rlabel metal2 9154 7174 9154 7174 0 net91
rlabel metal1 9890 7854 9890 7854 0 net92
rlabel metal2 10810 7718 10810 7718 0 net93
rlabel metal2 10994 5542 10994 5542 0 net94
rlabel metal1 12098 7310 12098 7310 0 net95
rlabel metal1 14214 2618 14214 2618 0 net96
rlabel metal1 13386 7310 13386 7310 0 net97
rlabel metal2 14306 4828 14306 4828 0 net98
rlabel metal1 14628 2550 14628 2550 0 net99
<< properties >>
string FIXED_BBOX 0 0 46000 10000
<< end >>
