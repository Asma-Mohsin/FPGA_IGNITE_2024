VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_IO
  CLASS BLOCK ;
  FOREIGN RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 181.000 BY 250.000 ;
  PIN Config_accessC_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 235.430 181.000 235.810 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 238.150 181.000 238.530 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 241.550 181.000 241.930 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 244.270 181.000 244.650 ;
    END
  END Config_accessC_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.550 0.700 3.930 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.590 0.700 5.970 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.950 0.700 7.330 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.990 0.700 9.370 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.990 0.700 26.370 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.030 0.700 28.410 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.070 0.700 30.450 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.110 0.700 32.490 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.470 0.700 33.850 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.510 0.700 35.890 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.550 0.700 37.930 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.590 0.700 39.970 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.030 0.700 11.410 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.070 0.700 13.450 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.430 0.700 14.810 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.470 0.700 16.850 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.510 0.700 18.890 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.550 0.700 20.930 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.590 0.700 22.970 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.950 0.700 24.330 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.550 0.700 71.930 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.590 0.700 90.970 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.630 0.700 93.010 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.590 0.700 73.970 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.630 0.700 76.010 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.670 0.700 78.050 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.030 0.700 79.410 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.070 0.700 81.450 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.110 0.700 83.490 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.150 0.700 85.530 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.190 0.700 87.570 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.550 0.700 88.930 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.630 0.700 42.010 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.670 0.700 61.050 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.030 0.700 62.410 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.070 0.700 64.450 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.110 0.700 66.490 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.150 0.700 68.530 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.510 0.700 69.890 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.990 0.700 43.370 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.030 0.700 45.410 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.070 0.700 47.450 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.110 0.700 49.490 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.150 0.700 51.530 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.510 0.700 52.890 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.550 0.700 54.930 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.590 0.700 56.970 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.630 0.700 59.010 ;
    END
  END EE4END[9]
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 198.710 181.000 199.090 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 202.110 181.000 202.490 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 204.830 181.000 205.210 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 208.230 181.000 208.610 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 210.950 181.000 211.330 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 214.350 181.000 214.730 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 217.070 181.000 217.450 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 220.470 181.000 220.850 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 223.190 181.000 223.570 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 225.910 181.000 226.290 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 229.310 181.000 229.690 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 232.030 181.000 232.410 ;
    END
  END FAB2RAM_C_O3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 150.430 181.000 150.810 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 153.150 181.000 153.530 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 156.550 181.000 156.930 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 159.270 181.000 159.650 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 162.670 181.000 163.050 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 165.390 181.000 165.770 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 168.790 181.000 169.170 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 171.510 181.000 171.890 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 174.910 181.000 175.290 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 177.630 181.000 178.010 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 180.350 181.000 180.730 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 183.750 181.000 184.130 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 186.470 181.000 186.850 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 189.870 181.000 190.250 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 192.590 181.000 192.970 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 195.990 181.000 196.370 ;
    END
  END FAB2RAM_D3_O3
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.790 0.700 186.170 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.830 0.700 205.210 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.870 0.700 207.250 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.230 0.700 208.610 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.270 0.700 210.650 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.310 0.700 212.690 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.350 0.700 214.730 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.390 0.700 216.770 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.750 0.700 218.130 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.790 0.700 220.170 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.830 0.700 222.210 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.830 0.700 188.210 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.870 0.700 224.250 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.230 0.700 225.610 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.270 0.700 227.650 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.310 0.700 229.690 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.350 0.700 231.730 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.390 0.700 233.770 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.750 0.700 235.130 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.790 0.700 237.170 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.830 0.700 239.210 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.870 0.700 241.250 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.190 0.700 189.570 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.910 0.700 243.290 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.270 0.700 244.650 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.230 0.700 191.610 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.270 0.700 193.650 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.310 0.700 195.690 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.350 0.700 197.730 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.710 0.700 199.090 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.750 0.700 201.130 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.790 0.700 203.170 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 4.230 181.000 4.610 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 34.830 181.000 35.210 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 38.230 181.000 38.610 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 40.950 181.000 41.330 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 43.670 181.000 44.050 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 47.070 181.000 47.450 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 49.790 181.000 50.170 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 53.190 181.000 53.570 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 55.910 181.000 56.290 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 59.310 181.000 59.690 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 62.030 181.000 62.410 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 7.630 181.000 8.010 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 65.430 181.000 65.810 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 68.150 181.000 68.530 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 71.550 181.000 71.930 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 74.270 181.000 74.650 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 77.670 181.000 78.050 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 80.390 181.000 80.770 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 83.790 181.000 84.170 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 86.510 181.000 86.890 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 89.230 181.000 89.610 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 92.630 181.000 93.010 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 10.350 181.000 10.730 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 95.350 181.000 95.730 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 98.750 181.000 99.130 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 13.750 181.000 14.130 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 16.470 181.000 16.850 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 19.870 181.000 20.250 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 22.590 181.000 22.970 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 25.990 181.000 26.370 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 28.710 181.000 29.090 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 32.110 181.000 32.490 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 138.960 0.000 139.340 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 157.820 0.000 158.200 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 159.660 0.000 160.040 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.500 0.000 161.880 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.340 0.000 163.720 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 165.180 0.000 165.560 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.480 0.000 167.860 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 169.320 0.000 169.700 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 171.160 0.000 171.540 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 173.000 0.000 173.380 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 174.840 0.000 175.220 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 140.800 0.000 141.180 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 142.640 0.000 143.020 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 144.480 0.000 144.860 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 146.780 0.000 147.160 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 148.620 0.000 149.000 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 150.460 0.000 150.840 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 152.300 0.000 152.680 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 154.140 0.000 154.520 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 155.980 0.000 156.360 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.960 249.300 139.340 250.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.820 249.300 158.200 250.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 159.660 249.300 160.040 250.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.500 249.300 161.880 250.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 163.340 249.300 163.720 250.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 165.180 249.300 165.560 250.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.480 249.300 167.860 250.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 169.320 249.300 169.700 250.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 171.160 249.300 171.540 250.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 173.000 249.300 173.380 250.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 174.840 249.300 175.220 250.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.800 249.300 141.180 250.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.640 249.300 143.020 250.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.480 249.300 144.860 250.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.780 249.300 147.160 250.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.620 249.300 149.000 250.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.460 249.300 150.840 250.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.300 249.300 152.680 250.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.140 249.300 154.520 250.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.980 249.300 156.360 250.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.260 249.300 3.640 250.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 5.560 249.300 5.940 250.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 7.400 249.300 7.780 250.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.240 249.300 9.620 250.000 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 3.260 0.000 3.640 0.700 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 5.560 0.000 5.940 0.700 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 7.400 0.000 7.780 0.700 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 9.240 0.000 9.620 0.700 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 11.080 249.300 11.460 250.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 12.920 249.300 13.300 250.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 14.760 249.300 15.140 250.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.600 249.300 16.980 250.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 18.440 249.300 18.820 250.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 20.280 249.300 20.660 250.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.120 249.300 22.500 250.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 23.960 249.300 24.340 250.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 26.260 249.300 26.640 250.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.100 249.300 28.480 250.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.940 249.300 30.320 250.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 31.780 249.300 32.160 250.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.620 249.300 34.000 250.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.460 249.300 35.840 250.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.300 249.300 37.680 250.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.140 249.300 39.520 250.000 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 26.260 0.000 26.640 0.700 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 28.100 0.000 28.480 0.700 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 29.940 0.000 30.320 0.700 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 31.780 0.000 32.160 0.700 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 33.620 0.000 34.000 0.700 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.460 0.000 35.840 0.700 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 37.300 0.000 37.680 0.700 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.140 0.000 39.520 0.700 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 11.080 0.000 11.460 0.700 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.920 0.000 13.300 0.700 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 14.760 0.000 15.140 0.700 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.600 0.000 16.980 0.700 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 18.440 0.000 18.820 0.700 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 20.280 0.000 20.660 0.700 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 22.120 0.000 22.500 0.700 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.960 0.000 24.340 0.700 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 40.980 249.300 41.360 250.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.840 249.300 60.220 250.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.680 249.300 62.060 250.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 63.520 249.300 63.900 250.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.820 249.300 66.200 250.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.660 249.300 68.040 250.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.500 249.300 69.880 250.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 42.820 249.300 43.200 250.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 44.660 249.300 45.040 250.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.960 249.300 47.340 250.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.800 249.300 49.180 250.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.640 249.300 51.020 250.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.480 249.300 52.860 250.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.320 249.300 54.700 250.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 56.160 249.300 56.540 250.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 249.300 58.380 250.000 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 40.980 0.000 41.360 0.700 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 59.840 0.000 60.220 0.700 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 61.680 0.000 62.060 0.700 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 63.520 0.000 63.900 0.700 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 65.820 0.000 66.200 0.700 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 67.660 0.000 68.040 0.700 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 69.500 0.000 69.880 0.700 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 42.820 0.000 43.200 0.700 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 44.660 0.000 45.040 0.700 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 46.960 0.000 47.340 0.700 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 48.800 0.000 49.180 0.700 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 50.640 0.000 51.020 0.700 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 52.480 0.000 52.860 0.700 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.320 0.000 54.700 0.700 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 56.160 0.000 56.540 0.700 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 58.000 0.000 58.380 0.700 ;
    END
  END N4END[9]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 101.470 181.000 101.850 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 104.870 181.000 105.250 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 107.590 181.000 107.970 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 110.990 181.000 111.370 ;
    END
  END RAM2FAB_D0_I3
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 113.710 181.000 114.090 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 117.110 181.000 117.490 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 119.830 181.000 120.210 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 123.230 181.000 123.610 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 125.950 181.000 126.330 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 129.350 181.000 129.730 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 132.070 181.000 132.450 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 134.790 181.000 135.170 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 138.190 181.000 138.570 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 140.910 181.000 141.290 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 144.310 181.000 144.690 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 147.030 181.000 147.410 ;
    END
  END RAM2FAB_D3_I3
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.340 0.000 71.720 0.700 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.180 0.000 73.560 0.700 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.020 0.000 75.400 0.700 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.860 0.000 77.240 0.700 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 71.340 249.300 71.720 250.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 73.180 249.300 73.560 250.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 75.020 249.300 75.400 250.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 76.860 249.300 77.240 250.000 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.700 0.000 79.080 0.700 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.540 0.000 80.920 0.700 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.380 0.000 82.760 0.700 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 84.220 0.000 84.600 0.700 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 0.000 86.900 0.700 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 88.360 0.000 88.740 0.700 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.200 0.000 90.580 0.700 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.040 0.000 92.420 0.700 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.880 0.000 94.260 0.700 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 95.720 0.000 96.100 0.700 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 97.560 0.000 97.940 0.700 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.400 0.000 99.780 0.700 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 101.240 0.000 101.620 0.700 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 103.080 0.000 103.460 0.700 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.920 0.000 105.300 0.700 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 107.220 0.000 107.600 0.700 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 93.880 249.300 94.260 250.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 95.720 249.300 96.100 250.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 97.560 249.300 97.940 250.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.400 249.300 99.780 250.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 101.240 249.300 101.620 250.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 103.080 249.300 103.460 250.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 104.920 249.300 105.300 250.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 107.220 249.300 107.600 250.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 78.700 249.300 79.080 250.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 80.540 249.300 80.920 250.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.380 249.300 82.760 250.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 84.220 249.300 84.600 250.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 249.300 86.900 250.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 88.360 249.300 88.740 250.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.200 249.300 90.580 250.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 92.040 249.300 92.420 250.000 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.060 0.000 109.440 0.700 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 127.920 0.000 128.300 0.700 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 129.760 0.000 130.140 0.700 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 131.600 0.000 131.980 0.700 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 133.440 0.000 133.820 0.700 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 135.280 0.000 135.660 0.700 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 137.120 0.000 137.500 0.700 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.900 0.000 111.280 0.700 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.740 0.000 113.120 0.700 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 114.580 0.000 114.960 0.700 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 116.420 0.000 116.800 0.700 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.260 0.000 118.640 0.700 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 120.100 0.000 120.480 0.700 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.940 0.000 122.320 0.700 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.780 0.000 124.160 0.700 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 126.080 0.000 126.460 0.700 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 109.060 249.300 109.440 250.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 127.920 249.300 128.300 250.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 129.760 249.300 130.140 250.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 131.600 249.300 131.980 250.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 133.440 249.300 133.820 250.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.280 249.300 135.660 250.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 137.120 249.300 137.500 250.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 110.900 249.300 111.280 250.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 112.740 249.300 113.120 250.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 114.580 249.300 114.960 250.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.420 249.300 116.800 250.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 118.260 249.300 118.640 250.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 120.100 249.300 120.480 250.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 121.940 249.300 122.320 250.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 123.780 249.300 124.160 250.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 126.080 249.300 126.460 250.000 ;
    END
  END S4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 176.680 0.000 177.060 0.700 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 176.680 249.300 177.060 250.000 ;
    END
  END UserCLKo
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.670 0.700 95.050 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.710 0.700 97.090 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.070 0.700 98.450 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.110 0.700 100.490 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.150 0.700 102.530 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.190 0.700 104.570 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.230 0.700 106.610 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.590 0.700 107.970 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.630 0.700 110.010 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.670 0.700 112.050 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.710 0.700 114.090 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.750 0.700 116.130 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.110 0.700 117.490 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.150 0.700 119.530 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.190 0.700 121.570 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.230 0.700 123.610 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.590 0.700 124.970 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.630 0.700 127.010 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.670 0.700 129.050 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.710 0.700 131.090 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.670 0.700 163.050 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.710 0.700 182.090 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.750 0.700 184.130 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.710 0.700 165.090 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.750 0.700 167.130 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.790 0.700 169.170 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.150 0.700 170.530 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.190 0.700 172.570 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.230 0.700 174.610 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.270 0.700 176.650 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.310 0.700 178.690 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.670 0.700 180.050 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.750 0.700 133.130 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.790 0.700 152.170 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.150 0.700 153.530 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.190 0.700 155.570 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.230 0.700 157.610 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.270 0.700 159.650 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.310 0.700 161.690 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.110 0.700 134.490 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.150 0.700 136.530 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.190 0.700 138.570 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.230 0.700 140.610 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.270 0.700 142.650 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.630 0.700 144.010 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.670 0.700 146.050 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.710 0.700 148.090 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.750 0.700 150.130 ;
    END
  END WW4BEG[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.580 5.200 22.180 245.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 5.200 175.780 245.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 21.290 175.960 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 174.470 175.960 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.880 5.200 25.480 245.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 175.720 244.885 ;
      LAYER met1 ;
        RECT 3.290 2.080 180.710 248.840 ;
      LAYER met2 ;
        RECT 3.920 249.020 5.280 249.300 ;
        RECT 6.220 249.020 7.120 249.300 ;
        RECT 8.060 249.020 8.960 249.300 ;
        RECT 9.900 249.020 10.800 249.300 ;
        RECT 11.740 249.020 12.640 249.300 ;
        RECT 13.580 249.020 14.480 249.300 ;
        RECT 15.420 249.020 16.320 249.300 ;
        RECT 17.260 249.020 18.160 249.300 ;
        RECT 19.100 249.020 20.000 249.300 ;
        RECT 20.940 249.020 21.840 249.300 ;
        RECT 22.780 249.020 23.680 249.300 ;
        RECT 24.620 249.020 25.980 249.300 ;
        RECT 26.920 249.020 27.820 249.300 ;
        RECT 28.760 249.020 29.660 249.300 ;
        RECT 30.600 249.020 31.500 249.300 ;
        RECT 32.440 249.020 33.340 249.300 ;
        RECT 34.280 249.020 35.180 249.300 ;
        RECT 36.120 249.020 37.020 249.300 ;
        RECT 37.960 249.020 38.860 249.300 ;
        RECT 39.800 249.020 40.700 249.300 ;
        RECT 41.640 249.020 42.540 249.300 ;
        RECT 43.480 249.020 44.380 249.300 ;
        RECT 45.320 249.020 46.680 249.300 ;
        RECT 47.620 249.020 48.520 249.300 ;
        RECT 49.460 249.020 50.360 249.300 ;
        RECT 51.300 249.020 52.200 249.300 ;
        RECT 53.140 249.020 54.040 249.300 ;
        RECT 54.980 249.020 55.880 249.300 ;
        RECT 56.820 249.020 57.720 249.300 ;
        RECT 58.660 249.020 59.560 249.300 ;
        RECT 60.500 249.020 61.400 249.300 ;
        RECT 62.340 249.020 63.240 249.300 ;
        RECT 64.180 249.020 65.540 249.300 ;
        RECT 66.480 249.020 67.380 249.300 ;
        RECT 68.320 249.020 69.220 249.300 ;
        RECT 70.160 249.020 71.060 249.300 ;
        RECT 72.000 249.020 72.900 249.300 ;
        RECT 73.840 249.020 74.740 249.300 ;
        RECT 75.680 249.020 76.580 249.300 ;
        RECT 77.520 249.020 78.420 249.300 ;
        RECT 79.360 249.020 80.260 249.300 ;
        RECT 81.200 249.020 82.100 249.300 ;
        RECT 83.040 249.020 83.940 249.300 ;
        RECT 84.880 249.020 86.240 249.300 ;
        RECT 87.180 249.020 88.080 249.300 ;
        RECT 89.020 249.020 89.920 249.300 ;
        RECT 90.860 249.020 91.760 249.300 ;
        RECT 92.700 249.020 93.600 249.300 ;
        RECT 94.540 249.020 95.440 249.300 ;
        RECT 96.380 249.020 97.280 249.300 ;
        RECT 98.220 249.020 99.120 249.300 ;
        RECT 100.060 249.020 100.960 249.300 ;
        RECT 101.900 249.020 102.800 249.300 ;
        RECT 103.740 249.020 104.640 249.300 ;
        RECT 105.580 249.020 106.940 249.300 ;
        RECT 107.880 249.020 108.780 249.300 ;
        RECT 109.720 249.020 110.620 249.300 ;
        RECT 111.560 249.020 112.460 249.300 ;
        RECT 113.400 249.020 114.300 249.300 ;
        RECT 115.240 249.020 116.140 249.300 ;
        RECT 117.080 249.020 117.980 249.300 ;
        RECT 118.920 249.020 119.820 249.300 ;
        RECT 120.760 249.020 121.660 249.300 ;
        RECT 122.600 249.020 123.500 249.300 ;
        RECT 124.440 249.020 125.800 249.300 ;
        RECT 126.740 249.020 127.640 249.300 ;
        RECT 128.580 249.020 129.480 249.300 ;
        RECT 130.420 249.020 131.320 249.300 ;
        RECT 132.260 249.020 133.160 249.300 ;
        RECT 134.100 249.020 135.000 249.300 ;
        RECT 135.940 249.020 136.840 249.300 ;
        RECT 137.780 249.020 138.680 249.300 ;
        RECT 139.620 249.020 140.520 249.300 ;
        RECT 141.460 249.020 142.360 249.300 ;
        RECT 143.300 249.020 144.200 249.300 ;
        RECT 145.140 249.020 146.500 249.300 ;
        RECT 147.440 249.020 148.340 249.300 ;
        RECT 149.280 249.020 150.180 249.300 ;
        RECT 151.120 249.020 152.020 249.300 ;
        RECT 152.960 249.020 153.860 249.300 ;
        RECT 154.800 249.020 155.700 249.300 ;
        RECT 156.640 249.020 157.540 249.300 ;
        RECT 158.480 249.020 159.380 249.300 ;
        RECT 160.320 249.020 161.220 249.300 ;
        RECT 162.160 249.020 163.060 249.300 ;
        RECT 164.000 249.020 164.900 249.300 ;
        RECT 165.840 249.020 167.200 249.300 ;
        RECT 168.140 249.020 169.040 249.300 ;
        RECT 169.980 249.020 170.880 249.300 ;
        RECT 171.820 249.020 172.720 249.300 ;
        RECT 173.660 249.020 174.560 249.300 ;
        RECT 175.500 249.020 176.400 249.300 ;
        RECT 177.340 249.020 180.680 249.300 ;
        RECT 3.320 0.980 180.680 249.020 ;
        RECT 3.920 0.270 5.280 0.980 ;
        RECT 6.220 0.270 7.120 0.980 ;
        RECT 8.060 0.270 8.960 0.980 ;
        RECT 9.900 0.270 10.800 0.980 ;
        RECT 11.740 0.270 12.640 0.980 ;
        RECT 13.580 0.270 14.480 0.980 ;
        RECT 15.420 0.270 16.320 0.980 ;
        RECT 17.260 0.270 18.160 0.980 ;
        RECT 19.100 0.270 20.000 0.980 ;
        RECT 20.940 0.270 21.840 0.980 ;
        RECT 22.780 0.270 23.680 0.980 ;
        RECT 24.620 0.270 25.980 0.980 ;
        RECT 26.920 0.270 27.820 0.980 ;
        RECT 28.760 0.270 29.660 0.980 ;
        RECT 30.600 0.270 31.500 0.980 ;
        RECT 32.440 0.270 33.340 0.980 ;
        RECT 34.280 0.270 35.180 0.980 ;
        RECT 36.120 0.270 37.020 0.980 ;
        RECT 37.960 0.270 38.860 0.980 ;
        RECT 39.800 0.270 40.700 0.980 ;
        RECT 41.640 0.270 42.540 0.980 ;
        RECT 43.480 0.270 44.380 0.980 ;
        RECT 45.320 0.270 46.680 0.980 ;
        RECT 47.620 0.270 48.520 0.980 ;
        RECT 49.460 0.270 50.360 0.980 ;
        RECT 51.300 0.270 52.200 0.980 ;
        RECT 53.140 0.270 54.040 0.980 ;
        RECT 54.980 0.270 55.880 0.980 ;
        RECT 56.820 0.270 57.720 0.980 ;
        RECT 58.660 0.270 59.560 0.980 ;
        RECT 60.500 0.270 61.400 0.980 ;
        RECT 62.340 0.270 63.240 0.980 ;
        RECT 64.180 0.270 65.540 0.980 ;
        RECT 66.480 0.270 67.380 0.980 ;
        RECT 68.320 0.270 69.220 0.980 ;
        RECT 70.160 0.270 71.060 0.980 ;
        RECT 72.000 0.270 72.900 0.980 ;
        RECT 73.840 0.270 74.740 0.980 ;
        RECT 75.680 0.270 76.580 0.980 ;
        RECT 77.520 0.270 78.420 0.980 ;
        RECT 79.360 0.270 80.260 0.980 ;
        RECT 81.200 0.270 82.100 0.980 ;
        RECT 83.040 0.270 83.940 0.980 ;
        RECT 84.880 0.270 86.240 0.980 ;
        RECT 87.180 0.270 88.080 0.980 ;
        RECT 89.020 0.270 89.920 0.980 ;
        RECT 90.860 0.270 91.760 0.980 ;
        RECT 92.700 0.270 93.600 0.980 ;
        RECT 94.540 0.270 95.440 0.980 ;
        RECT 96.380 0.270 97.280 0.980 ;
        RECT 98.220 0.270 99.120 0.980 ;
        RECT 100.060 0.270 100.960 0.980 ;
        RECT 101.900 0.270 102.800 0.980 ;
        RECT 103.740 0.270 104.640 0.980 ;
        RECT 105.580 0.270 106.940 0.980 ;
        RECT 107.880 0.270 108.780 0.980 ;
        RECT 109.720 0.270 110.620 0.980 ;
        RECT 111.560 0.270 112.460 0.980 ;
        RECT 113.400 0.270 114.300 0.980 ;
        RECT 115.240 0.270 116.140 0.980 ;
        RECT 117.080 0.270 117.980 0.980 ;
        RECT 118.920 0.270 119.820 0.980 ;
        RECT 120.760 0.270 121.660 0.980 ;
        RECT 122.600 0.270 123.500 0.980 ;
        RECT 124.440 0.270 125.800 0.980 ;
        RECT 126.740 0.270 127.640 0.980 ;
        RECT 128.580 0.270 129.480 0.980 ;
        RECT 130.420 0.270 131.320 0.980 ;
        RECT 132.260 0.270 133.160 0.980 ;
        RECT 134.100 0.270 135.000 0.980 ;
        RECT 135.940 0.270 136.840 0.980 ;
        RECT 137.780 0.270 138.680 0.980 ;
        RECT 139.620 0.270 140.520 0.980 ;
        RECT 141.460 0.270 142.360 0.980 ;
        RECT 143.300 0.270 144.200 0.980 ;
        RECT 145.140 0.270 146.500 0.980 ;
        RECT 147.440 0.270 148.340 0.980 ;
        RECT 149.280 0.270 150.180 0.980 ;
        RECT 151.120 0.270 152.020 0.980 ;
        RECT 152.960 0.270 153.860 0.980 ;
        RECT 154.800 0.270 155.700 0.980 ;
        RECT 156.640 0.270 157.540 0.980 ;
        RECT 158.480 0.270 159.380 0.980 ;
        RECT 160.320 0.270 161.220 0.980 ;
        RECT 162.160 0.270 163.060 0.980 ;
        RECT 164.000 0.270 164.900 0.980 ;
        RECT 165.840 0.270 167.200 0.980 ;
        RECT 168.140 0.270 169.040 0.980 ;
        RECT 169.980 0.270 170.880 0.980 ;
        RECT 171.820 0.270 172.720 0.980 ;
        RECT 173.660 0.270 174.560 0.980 ;
        RECT 175.500 0.270 176.400 0.980 ;
        RECT 177.340 0.270 180.680 0.980 ;
      LAYER met3 ;
        RECT 1.100 243.870 179.900 244.965 ;
        RECT 0.700 243.690 180.300 243.870 ;
        RECT 1.100 242.510 180.300 243.690 ;
        RECT 0.700 242.330 180.300 242.510 ;
        RECT 0.700 241.650 179.900 242.330 ;
        RECT 1.100 241.150 179.900 241.650 ;
        RECT 1.100 240.470 180.300 241.150 ;
        RECT 0.700 239.610 180.300 240.470 ;
        RECT 1.100 238.930 180.300 239.610 ;
        RECT 1.100 238.430 179.900 238.930 ;
        RECT 0.700 237.750 179.900 238.430 ;
        RECT 0.700 237.570 180.300 237.750 ;
        RECT 1.100 236.390 180.300 237.570 ;
        RECT 0.700 236.210 180.300 236.390 ;
        RECT 0.700 235.530 179.900 236.210 ;
        RECT 1.100 235.030 179.900 235.530 ;
        RECT 1.100 234.350 180.300 235.030 ;
        RECT 0.700 234.170 180.300 234.350 ;
        RECT 1.100 232.990 180.300 234.170 ;
        RECT 0.700 232.810 180.300 232.990 ;
        RECT 0.700 232.130 179.900 232.810 ;
        RECT 1.100 231.630 179.900 232.130 ;
        RECT 1.100 230.950 180.300 231.630 ;
        RECT 0.700 230.090 180.300 230.950 ;
        RECT 1.100 228.910 179.900 230.090 ;
        RECT 0.700 228.050 180.300 228.910 ;
        RECT 1.100 226.870 180.300 228.050 ;
        RECT 0.700 226.690 180.300 226.870 ;
        RECT 0.700 226.010 179.900 226.690 ;
        RECT 1.100 225.510 179.900 226.010 ;
        RECT 1.100 224.830 180.300 225.510 ;
        RECT 0.700 224.650 180.300 224.830 ;
        RECT 1.100 223.970 180.300 224.650 ;
        RECT 1.100 223.470 179.900 223.970 ;
        RECT 0.700 222.790 179.900 223.470 ;
        RECT 0.700 222.610 180.300 222.790 ;
        RECT 1.100 221.430 180.300 222.610 ;
        RECT 0.700 221.250 180.300 221.430 ;
        RECT 0.700 220.570 179.900 221.250 ;
        RECT 1.100 220.070 179.900 220.570 ;
        RECT 1.100 219.390 180.300 220.070 ;
        RECT 0.700 218.530 180.300 219.390 ;
        RECT 1.100 217.850 180.300 218.530 ;
        RECT 1.100 217.350 179.900 217.850 ;
        RECT 0.700 217.170 179.900 217.350 ;
        RECT 1.100 216.670 179.900 217.170 ;
        RECT 1.100 215.990 180.300 216.670 ;
        RECT 0.700 215.130 180.300 215.990 ;
        RECT 1.100 213.950 179.900 215.130 ;
        RECT 0.700 213.090 180.300 213.950 ;
        RECT 1.100 211.910 180.300 213.090 ;
        RECT 0.700 211.730 180.300 211.910 ;
        RECT 0.700 211.050 179.900 211.730 ;
        RECT 1.100 210.550 179.900 211.050 ;
        RECT 1.100 209.870 180.300 210.550 ;
        RECT 0.700 209.010 180.300 209.870 ;
        RECT 1.100 207.830 179.900 209.010 ;
        RECT 0.700 207.650 180.300 207.830 ;
        RECT 1.100 206.470 180.300 207.650 ;
        RECT 0.700 205.610 180.300 206.470 ;
        RECT 1.100 204.430 179.900 205.610 ;
        RECT 0.700 203.570 180.300 204.430 ;
        RECT 1.100 202.890 180.300 203.570 ;
        RECT 1.100 202.390 179.900 202.890 ;
        RECT 0.700 201.710 179.900 202.390 ;
        RECT 0.700 201.530 180.300 201.710 ;
        RECT 1.100 200.350 180.300 201.530 ;
        RECT 0.700 199.490 180.300 200.350 ;
        RECT 1.100 198.310 179.900 199.490 ;
        RECT 0.700 198.130 180.300 198.310 ;
        RECT 1.100 196.950 180.300 198.130 ;
        RECT 0.700 196.770 180.300 196.950 ;
        RECT 0.700 196.090 179.900 196.770 ;
        RECT 1.100 195.590 179.900 196.090 ;
        RECT 1.100 194.910 180.300 195.590 ;
        RECT 0.700 194.050 180.300 194.910 ;
        RECT 1.100 193.370 180.300 194.050 ;
        RECT 1.100 192.870 179.900 193.370 ;
        RECT 0.700 192.190 179.900 192.870 ;
        RECT 0.700 192.010 180.300 192.190 ;
        RECT 1.100 190.830 180.300 192.010 ;
        RECT 0.700 190.650 180.300 190.830 ;
        RECT 0.700 189.970 179.900 190.650 ;
        RECT 1.100 189.470 179.900 189.970 ;
        RECT 1.100 188.790 180.300 189.470 ;
        RECT 0.700 188.610 180.300 188.790 ;
        RECT 1.100 187.430 180.300 188.610 ;
        RECT 0.700 187.250 180.300 187.430 ;
        RECT 0.700 186.570 179.900 187.250 ;
        RECT 1.100 186.070 179.900 186.570 ;
        RECT 1.100 185.390 180.300 186.070 ;
        RECT 0.700 184.530 180.300 185.390 ;
        RECT 1.100 183.350 179.900 184.530 ;
        RECT 0.700 182.490 180.300 183.350 ;
        RECT 1.100 181.310 180.300 182.490 ;
        RECT 0.700 181.130 180.300 181.310 ;
        RECT 0.700 180.450 179.900 181.130 ;
        RECT 1.100 179.950 179.900 180.450 ;
        RECT 1.100 179.270 180.300 179.950 ;
        RECT 0.700 179.090 180.300 179.270 ;
        RECT 1.100 178.410 180.300 179.090 ;
        RECT 1.100 177.910 179.900 178.410 ;
        RECT 0.700 177.230 179.900 177.910 ;
        RECT 0.700 177.050 180.300 177.230 ;
        RECT 1.100 175.870 180.300 177.050 ;
        RECT 0.700 175.690 180.300 175.870 ;
        RECT 0.700 175.010 179.900 175.690 ;
        RECT 1.100 174.510 179.900 175.010 ;
        RECT 1.100 173.830 180.300 174.510 ;
        RECT 0.700 172.970 180.300 173.830 ;
        RECT 1.100 172.290 180.300 172.970 ;
        RECT 1.100 171.790 179.900 172.290 ;
        RECT 0.700 171.110 179.900 171.790 ;
        RECT 0.700 170.930 180.300 171.110 ;
        RECT 1.100 169.750 180.300 170.930 ;
        RECT 0.700 169.570 180.300 169.750 ;
        RECT 1.100 168.390 179.900 169.570 ;
        RECT 0.700 167.530 180.300 168.390 ;
        RECT 1.100 166.350 180.300 167.530 ;
        RECT 0.700 166.170 180.300 166.350 ;
        RECT 0.700 165.490 179.900 166.170 ;
        RECT 1.100 164.990 179.900 165.490 ;
        RECT 1.100 164.310 180.300 164.990 ;
        RECT 0.700 163.450 180.300 164.310 ;
        RECT 1.100 162.270 179.900 163.450 ;
        RECT 0.700 162.090 180.300 162.270 ;
        RECT 1.100 160.910 180.300 162.090 ;
        RECT 0.700 160.050 180.300 160.910 ;
        RECT 1.100 158.870 179.900 160.050 ;
        RECT 0.700 158.010 180.300 158.870 ;
        RECT 1.100 157.330 180.300 158.010 ;
        RECT 1.100 156.830 179.900 157.330 ;
        RECT 0.700 156.150 179.900 156.830 ;
        RECT 0.700 155.970 180.300 156.150 ;
        RECT 1.100 154.790 180.300 155.970 ;
        RECT 0.700 153.930 180.300 154.790 ;
        RECT 1.100 152.750 179.900 153.930 ;
        RECT 0.700 152.570 180.300 152.750 ;
        RECT 1.100 151.390 180.300 152.570 ;
        RECT 0.700 151.210 180.300 151.390 ;
        RECT 0.700 150.530 179.900 151.210 ;
        RECT 1.100 150.030 179.900 150.530 ;
        RECT 1.100 149.350 180.300 150.030 ;
        RECT 0.700 148.490 180.300 149.350 ;
        RECT 1.100 147.810 180.300 148.490 ;
        RECT 1.100 147.310 179.900 147.810 ;
        RECT 0.700 146.630 179.900 147.310 ;
        RECT 0.700 146.450 180.300 146.630 ;
        RECT 1.100 145.270 180.300 146.450 ;
        RECT 0.700 145.090 180.300 145.270 ;
        RECT 0.700 144.410 179.900 145.090 ;
        RECT 1.100 143.910 179.900 144.410 ;
        RECT 1.100 143.230 180.300 143.910 ;
        RECT 0.700 143.050 180.300 143.230 ;
        RECT 1.100 141.870 180.300 143.050 ;
        RECT 0.700 141.690 180.300 141.870 ;
        RECT 0.700 141.010 179.900 141.690 ;
        RECT 1.100 140.510 179.900 141.010 ;
        RECT 1.100 139.830 180.300 140.510 ;
        RECT 0.700 138.970 180.300 139.830 ;
        RECT 1.100 137.790 179.900 138.970 ;
        RECT 0.700 136.930 180.300 137.790 ;
        RECT 1.100 135.750 180.300 136.930 ;
        RECT 0.700 135.570 180.300 135.750 ;
        RECT 0.700 134.890 179.900 135.570 ;
        RECT 1.100 134.390 179.900 134.890 ;
        RECT 1.100 133.710 180.300 134.390 ;
        RECT 0.700 133.530 180.300 133.710 ;
        RECT 1.100 132.850 180.300 133.530 ;
        RECT 1.100 132.350 179.900 132.850 ;
        RECT 0.700 131.670 179.900 132.350 ;
        RECT 0.700 131.490 180.300 131.670 ;
        RECT 1.100 130.310 180.300 131.490 ;
        RECT 0.700 130.130 180.300 130.310 ;
        RECT 0.700 129.450 179.900 130.130 ;
        RECT 1.100 128.950 179.900 129.450 ;
        RECT 1.100 128.270 180.300 128.950 ;
        RECT 0.700 127.410 180.300 128.270 ;
        RECT 1.100 126.730 180.300 127.410 ;
        RECT 1.100 126.230 179.900 126.730 ;
        RECT 0.700 125.550 179.900 126.230 ;
        RECT 0.700 125.370 180.300 125.550 ;
        RECT 1.100 124.190 180.300 125.370 ;
        RECT 0.700 124.010 180.300 124.190 ;
        RECT 1.100 122.830 179.900 124.010 ;
        RECT 0.700 121.970 180.300 122.830 ;
        RECT 1.100 120.790 180.300 121.970 ;
        RECT 0.700 120.610 180.300 120.790 ;
        RECT 0.700 119.930 179.900 120.610 ;
        RECT 1.100 119.430 179.900 119.930 ;
        RECT 1.100 118.750 180.300 119.430 ;
        RECT 0.700 117.890 180.300 118.750 ;
        RECT 1.100 116.710 179.900 117.890 ;
        RECT 0.700 116.530 180.300 116.710 ;
        RECT 1.100 115.350 180.300 116.530 ;
        RECT 0.700 114.490 180.300 115.350 ;
        RECT 1.100 113.310 179.900 114.490 ;
        RECT 0.700 112.450 180.300 113.310 ;
        RECT 1.100 111.770 180.300 112.450 ;
        RECT 1.100 111.270 179.900 111.770 ;
        RECT 0.700 110.590 179.900 111.270 ;
        RECT 0.700 110.410 180.300 110.590 ;
        RECT 1.100 109.230 180.300 110.410 ;
        RECT 0.700 108.370 180.300 109.230 ;
        RECT 1.100 107.190 179.900 108.370 ;
        RECT 0.700 107.010 180.300 107.190 ;
        RECT 1.100 105.830 180.300 107.010 ;
        RECT 0.700 105.650 180.300 105.830 ;
        RECT 0.700 104.970 179.900 105.650 ;
        RECT 1.100 104.470 179.900 104.970 ;
        RECT 1.100 103.790 180.300 104.470 ;
        RECT 0.700 102.930 180.300 103.790 ;
        RECT 1.100 102.250 180.300 102.930 ;
        RECT 1.100 101.750 179.900 102.250 ;
        RECT 0.700 101.070 179.900 101.750 ;
        RECT 0.700 100.890 180.300 101.070 ;
        RECT 1.100 99.710 180.300 100.890 ;
        RECT 0.700 99.530 180.300 99.710 ;
        RECT 0.700 98.850 179.900 99.530 ;
        RECT 1.100 98.350 179.900 98.850 ;
        RECT 1.100 97.670 180.300 98.350 ;
        RECT 0.700 97.490 180.300 97.670 ;
        RECT 1.100 96.310 180.300 97.490 ;
        RECT 0.700 96.130 180.300 96.310 ;
        RECT 0.700 95.450 179.900 96.130 ;
        RECT 1.100 94.950 179.900 95.450 ;
        RECT 1.100 94.270 180.300 94.950 ;
        RECT 0.700 93.410 180.300 94.270 ;
        RECT 1.100 92.230 179.900 93.410 ;
        RECT 0.700 91.370 180.300 92.230 ;
        RECT 1.100 90.190 180.300 91.370 ;
        RECT 0.700 90.010 180.300 90.190 ;
        RECT 0.700 89.330 179.900 90.010 ;
        RECT 1.100 88.830 179.900 89.330 ;
        RECT 1.100 88.150 180.300 88.830 ;
        RECT 0.700 87.970 180.300 88.150 ;
        RECT 1.100 87.290 180.300 87.970 ;
        RECT 1.100 86.790 179.900 87.290 ;
        RECT 0.700 86.110 179.900 86.790 ;
        RECT 0.700 85.930 180.300 86.110 ;
        RECT 1.100 84.750 180.300 85.930 ;
        RECT 0.700 84.570 180.300 84.750 ;
        RECT 0.700 83.890 179.900 84.570 ;
        RECT 1.100 83.390 179.900 83.890 ;
        RECT 1.100 82.710 180.300 83.390 ;
        RECT 0.700 81.850 180.300 82.710 ;
        RECT 1.100 81.170 180.300 81.850 ;
        RECT 1.100 80.670 179.900 81.170 ;
        RECT 0.700 79.990 179.900 80.670 ;
        RECT 0.700 79.810 180.300 79.990 ;
        RECT 1.100 78.630 180.300 79.810 ;
        RECT 0.700 78.450 180.300 78.630 ;
        RECT 1.100 77.270 179.900 78.450 ;
        RECT 0.700 76.410 180.300 77.270 ;
        RECT 1.100 75.230 180.300 76.410 ;
        RECT 0.700 75.050 180.300 75.230 ;
        RECT 0.700 74.370 179.900 75.050 ;
        RECT 1.100 73.870 179.900 74.370 ;
        RECT 1.100 73.190 180.300 73.870 ;
        RECT 0.700 72.330 180.300 73.190 ;
        RECT 1.100 71.150 179.900 72.330 ;
        RECT 0.700 70.290 180.300 71.150 ;
        RECT 1.100 69.110 180.300 70.290 ;
        RECT 0.700 68.930 180.300 69.110 ;
        RECT 1.100 67.750 179.900 68.930 ;
        RECT 0.700 66.890 180.300 67.750 ;
        RECT 1.100 66.210 180.300 66.890 ;
        RECT 1.100 65.710 179.900 66.210 ;
        RECT 0.700 65.030 179.900 65.710 ;
        RECT 0.700 64.850 180.300 65.030 ;
        RECT 1.100 63.670 180.300 64.850 ;
        RECT 0.700 62.810 180.300 63.670 ;
        RECT 1.100 61.630 179.900 62.810 ;
        RECT 0.700 61.450 180.300 61.630 ;
        RECT 1.100 60.270 180.300 61.450 ;
        RECT 0.700 60.090 180.300 60.270 ;
        RECT 0.700 59.410 179.900 60.090 ;
        RECT 1.100 58.910 179.900 59.410 ;
        RECT 1.100 58.230 180.300 58.910 ;
        RECT 0.700 57.370 180.300 58.230 ;
        RECT 1.100 56.690 180.300 57.370 ;
        RECT 1.100 56.190 179.900 56.690 ;
        RECT 0.700 55.510 179.900 56.190 ;
        RECT 0.700 55.330 180.300 55.510 ;
        RECT 1.100 54.150 180.300 55.330 ;
        RECT 0.700 53.970 180.300 54.150 ;
        RECT 0.700 53.290 179.900 53.970 ;
        RECT 1.100 52.790 179.900 53.290 ;
        RECT 1.100 52.110 180.300 52.790 ;
        RECT 0.700 51.930 180.300 52.110 ;
        RECT 1.100 50.750 180.300 51.930 ;
        RECT 0.700 50.570 180.300 50.750 ;
        RECT 0.700 49.890 179.900 50.570 ;
        RECT 1.100 49.390 179.900 49.890 ;
        RECT 1.100 48.710 180.300 49.390 ;
        RECT 0.700 47.850 180.300 48.710 ;
        RECT 1.100 46.670 179.900 47.850 ;
        RECT 0.700 45.810 180.300 46.670 ;
        RECT 1.100 44.630 180.300 45.810 ;
        RECT 0.700 44.450 180.300 44.630 ;
        RECT 0.700 43.770 179.900 44.450 ;
        RECT 1.100 43.270 179.900 43.770 ;
        RECT 1.100 42.590 180.300 43.270 ;
        RECT 0.700 42.410 180.300 42.590 ;
        RECT 1.100 41.730 180.300 42.410 ;
        RECT 1.100 41.230 179.900 41.730 ;
        RECT 0.700 40.550 179.900 41.230 ;
        RECT 0.700 40.370 180.300 40.550 ;
        RECT 1.100 39.190 180.300 40.370 ;
        RECT 0.700 39.010 180.300 39.190 ;
        RECT 0.700 38.330 179.900 39.010 ;
        RECT 1.100 37.830 179.900 38.330 ;
        RECT 1.100 37.150 180.300 37.830 ;
        RECT 0.700 36.290 180.300 37.150 ;
        RECT 1.100 35.610 180.300 36.290 ;
        RECT 1.100 35.110 179.900 35.610 ;
        RECT 0.700 34.430 179.900 35.110 ;
        RECT 0.700 34.250 180.300 34.430 ;
        RECT 1.100 33.070 180.300 34.250 ;
        RECT 0.700 32.890 180.300 33.070 ;
        RECT 1.100 31.710 179.900 32.890 ;
        RECT 0.700 30.850 180.300 31.710 ;
        RECT 1.100 29.670 180.300 30.850 ;
        RECT 0.700 29.490 180.300 29.670 ;
        RECT 0.700 28.810 179.900 29.490 ;
        RECT 1.100 28.310 179.900 28.810 ;
        RECT 1.100 27.630 180.300 28.310 ;
        RECT 0.700 26.770 180.300 27.630 ;
        RECT 1.100 25.590 179.900 26.770 ;
        RECT 0.700 24.730 180.300 25.590 ;
        RECT 1.100 23.550 180.300 24.730 ;
        RECT 0.700 23.370 180.300 23.550 ;
        RECT 1.100 22.190 179.900 23.370 ;
        RECT 0.700 21.330 180.300 22.190 ;
        RECT 1.100 20.650 180.300 21.330 ;
        RECT 1.100 20.150 179.900 20.650 ;
        RECT 0.700 19.470 179.900 20.150 ;
        RECT 0.700 19.290 180.300 19.470 ;
        RECT 1.100 18.110 180.300 19.290 ;
        RECT 0.700 17.250 180.300 18.110 ;
        RECT 1.100 16.070 179.900 17.250 ;
        RECT 0.700 15.210 180.300 16.070 ;
        RECT 1.100 14.530 180.300 15.210 ;
        RECT 1.100 14.030 179.900 14.530 ;
        RECT 0.700 13.850 179.900 14.030 ;
        RECT 1.100 13.350 179.900 13.850 ;
        RECT 1.100 12.670 180.300 13.350 ;
        RECT 0.700 11.810 180.300 12.670 ;
        RECT 1.100 11.130 180.300 11.810 ;
        RECT 1.100 10.630 179.900 11.130 ;
        RECT 0.700 9.950 179.900 10.630 ;
        RECT 0.700 9.770 180.300 9.950 ;
        RECT 1.100 8.590 180.300 9.770 ;
        RECT 0.700 8.410 180.300 8.590 ;
        RECT 0.700 7.730 179.900 8.410 ;
        RECT 1.100 7.230 179.900 7.730 ;
        RECT 1.100 6.550 180.300 7.230 ;
        RECT 0.700 6.370 180.300 6.550 ;
        RECT 1.100 5.190 180.300 6.370 ;
        RECT 0.700 5.010 180.300 5.190 ;
        RECT 0.700 4.330 179.900 5.010 ;
        RECT 1.100 3.830 179.900 4.330 ;
        RECT 1.100 3.575 180.300 3.830 ;
      LAYER met4 ;
        RECT 8.575 4.800 20.180 243.945 ;
        RECT 22.580 4.800 23.480 243.945 ;
        RECT 25.880 4.800 170.825 243.945 ;
        RECT 8.575 4.255 170.825 4.800 ;
  END
END RAM_IO
END LIBRARY

