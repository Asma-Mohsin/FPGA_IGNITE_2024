VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_RAM_IO
  CLASS BLOCK ;
  FOREIGN N_term_RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 40.000 ;
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 10.670 39.200 10.950 40.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.470 39.200 70.750 40.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 76.450 39.200 76.730 40.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.430 39.200 82.710 40.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 88.410 39.200 88.690 40.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 94.390 39.200 94.670 40.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 100.370 39.200 100.650 40.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 39.200 106.630 40.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 112.330 39.200 112.610 40.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 118.310 39.200 118.590 40.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 124.290 39.200 124.570 40.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 16.650 39.200 16.930 40.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.630 39.200 22.910 40.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.610 39.200 28.890 40.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 34.590 39.200 34.870 40.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 40.570 39.200 40.850 40.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 46.550 39.200 46.830 40.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 52.530 39.200 52.810 40.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.510 39.200 58.790 40.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 39.200 64.770 40.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 0.800 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 0.800 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 0.800 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 0.800 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 0.800 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 0.800 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 20.330 0.000 20.610 0.800 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 0.800 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 0.800 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 0.800 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 0.800 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 0.800 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 0.800 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 0.800 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 0.800 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 0.800 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 0.800 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 0.800 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 0.800 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 0.800 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 0.800 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 0.800 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.800 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 0.800 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 0.800 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 0.800 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 0.800 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 0.800 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 0.800 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 0.800 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 0.800 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.800 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 0.800 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.800 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.800 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 0.800 ;
    END
  END N4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 0.800 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 0.800 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 0.800 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 0.800 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 0.800 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 0.800 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 0.800 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 0.800 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 0.800 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 0.800 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 0.800 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 0.800 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 0.800 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 0.800 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.800 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 0.800 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 0.800 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 0.800 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 0.800 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 0.800 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 0.800 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 0.800 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 0.800 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 0.800 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 0.800 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 0.800 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 0.800 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 0.800 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 0.800 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 0.800 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 0.800 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 0.800 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 0.800 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 0.800 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 0.800 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 0.800 ;
    END
  END S4BEG[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 4.690 39.200 4.970 40.000 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.390 5.200 35.990 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.060 5.200 65.660 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.730 5.200 95.330 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.400 5.200 125.000 32.880 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.555 5.200 21.155 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.225 5.200 50.825 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.895 5.200 80.495 32.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.565 5.200 110.165 32.880 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 124.200 32.725 ;
      LAYER met1 ;
        RECT 0.990 1.060 128.270 32.880 ;
      LAYER met2 ;
        RECT 1.020 38.920 4.410 39.850 ;
        RECT 5.250 38.920 10.390 39.850 ;
        RECT 11.230 38.920 16.370 39.850 ;
        RECT 17.210 38.920 22.350 39.850 ;
        RECT 23.190 38.920 28.330 39.850 ;
        RECT 29.170 38.920 34.310 39.850 ;
        RECT 35.150 38.920 40.290 39.850 ;
        RECT 41.130 38.920 46.270 39.850 ;
        RECT 47.110 38.920 52.250 39.850 ;
        RECT 53.090 38.920 58.230 39.850 ;
        RECT 59.070 38.920 64.210 39.850 ;
        RECT 65.050 38.920 70.190 39.850 ;
        RECT 71.030 38.920 76.170 39.850 ;
        RECT 77.010 38.920 82.150 39.850 ;
        RECT 82.990 38.920 88.130 39.850 ;
        RECT 88.970 38.920 94.110 39.850 ;
        RECT 94.950 38.920 100.090 39.850 ;
        RECT 100.930 38.920 106.070 39.850 ;
        RECT 106.910 38.920 112.050 39.850 ;
        RECT 112.890 38.920 118.030 39.850 ;
        RECT 118.870 38.920 124.010 39.850 ;
        RECT 124.850 38.920 128.240 39.850 ;
        RECT 1.020 1.080 128.240 38.920 ;
        RECT 1.570 0.270 2.110 1.080 ;
        RECT 2.950 0.270 3.490 1.080 ;
        RECT 4.330 0.270 4.870 1.080 ;
        RECT 5.710 0.270 6.250 1.080 ;
        RECT 7.090 0.270 7.630 1.080 ;
        RECT 8.470 0.270 9.010 1.080 ;
        RECT 9.850 0.270 10.390 1.080 ;
        RECT 11.230 0.270 11.770 1.080 ;
        RECT 12.610 0.270 13.150 1.080 ;
        RECT 13.990 0.270 14.530 1.080 ;
        RECT 15.370 0.270 15.910 1.080 ;
        RECT 16.750 0.270 17.290 1.080 ;
        RECT 18.130 0.270 18.670 1.080 ;
        RECT 19.510 0.270 20.050 1.080 ;
        RECT 20.890 0.270 21.430 1.080 ;
        RECT 22.270 0.270 22.810 1.080 ;
        RECT 23.650 0.270 24.190 1.080 ;
        RECT 25.030 0.270 25.570 1.080 ;
        RECT 26.410 0.270 26.950 1.080 ;
        RECT 27.790 0.270 28.330 1.080 ;
        RECT 29.170 0.270 29.710 1.080 ;
        RECT 30.550 0.270 31.090 1.080 ;
        RECT 31.930 0.270 32.470 1.080 ;
        RECT 33.310 0.270 33.850 1.080 ;
        RECT 34.690 0.270 35.230 1.080 ;
        RECT 36.070 0.270 36.610 1.080 ;
        RECT 37.450 0.270 37.990 1.080 ;
        RECT 38.830 0.270 39.370 1.080 ;
        RECT 40.210 0.270 40.750 1.080 ;
        RECT 41.590 0.270 42.130 1.080 ;
        RECT 42.970 0.270 43.510 1.080 ;
        RECT 44.350 0.270 44.890 1.080 ;
        RECT 45.730 0.270 46.270 1.080 ;
        RECT 47.110 0.270 47.650 1.080 ;
        RECT 48.490 0.270 49.030 1.080 ;
        RECT 49.870 0.270 50.410 1.080 ;
        RECT 51.250 0.270 51.790 1.080 ;
        RECT 52.630 0.270 53.170 1.080 ;
        RECT 54.010 0.270 54.550 1.080 ;
        RECT 55.390 0.270 55.930 1.080 ;
        RECT 56.770 0.270 57.310 1.080 ;
        RECT 58.150 0.270 58.690 1.080 ;
        RECT 59.530 0.270 60.070 1.080 ;
        RECT 60.910 0.270 61.450 1.080 ;
        RECT 62.290 0.270 62.830 1.080 ;
        RECT 63.670 0.270 64.210 1.080 ;
        RECT 65.050 0.270 65.590 1.080 ;
        RECT 66.430 0.270 66.970 1.080 ;
        RECT 67.810 0.270 68.350 1.080 ;
        RECT 69.190 0.270 69.730 1.080 ;
        RECT 70.570 0.270 71.110 1.080 ;
        RECT 71.950 0.270 72.490 1.080 ;
        RECT 73.330 0.270 73.870 1.080 ;
        RECT 74.710 0.270 75.250 1.080 ;
        RECT 76.090 0.270 76.630 1.080 ;
        RECT 77.470 0.270 78.010 1.080 ;
        RECT 78.850 0.270 79.390 1.080 ;
        RECT 80.230 0.270 80.770 1.080 ;
        RECT 81.610 0.270 82.150 1.080 ;
        RECT 82.990 0.270 83.530 1.080 ;
        RECT 84.370 0.270 84.910 1.080 ;
        RECT 85.750 0.270 86.290 1.080 ;
        RECT 87.130 0.270 87.670 1.080 ;
        RECT 88.510 0.270 89.050 1.080 ;
        RECT 89.890 0.270 90.430 1.080 ;
        RECT 91.270 0.270 91.810 1.080 ;
        RECT 92.650 0.270 93.190 1.080 ;
        RECT 94.030 0.270 94.570 1.080 ;
        RECT 95.410 0.270 95.950 1.080 ;
        RECT 96.790 0.270 97.330 1.080 ;
        RECT 98.170 0.270 98.710 1.080 ;
        RECT 99.550 0.270 100.090 1.080 ;
        RECT 100.930 0.270 101.470 1.080 ;
        RECT 102.310 0.270 102.850 1.080 ;
        RECT 103.690 0.270 104.230 1.080 ;
        RECT 105.070 0.270 105.610 1.080 ;
        RECT 106.450 0.270 106.990 1.080 ;
        RECT 107.830 0.270 108.370 1.080 ;
        RECT 109.210 0.270 109.750 1.080 ;
        RECT 110.590 0.270 111.130 1.080 ;
        RECT 111.970 0.270 112.510 1.080 ;
        RECT 113.350 0.270 113.890 1.080 ;
        RECT 114.730 0.270 115.270 1.080 ;
        RECT 116.110 0.270 116.650 1.080 ;
        RECT 117.490 0.270 118.030 1.080 ;
        RECT 118.870 0.270 119.410 1.080 ;
        RECT 120.250 0.270 120.790 1.080 ;
        RECT 121.630 0.270 122.170 1.080 ;
        RECT 123.010 0.270 123.550 1.080 ;
        RECT 124.390 0.270 124.930 1.080 ;
        RECT 125.770 0.270 126.310 1.080 ;
        RECT 127.150 0.270 127.690 1.080 ;
      LAYER met3 ;
        RECT 7.425 2.895 124.990 32.805 ;
      LAYER met4 ;
        RECT 12.750 4.800 19.155 20.905 ;
        RECT 21.555 4.800 33.990 20.905 ;
        RECT 36.390 4.800 48.825 20.905 ;
        RECT 51.225 4.800 63.660 20.905 ;
        RECT 66.060 4.800 78.495 20.905 ;
        RECT 80.895 4.800 93.330 20.905 ;
        RECT 95.730 4.800 108.165 20.905 ;
        RECT 110.565 4.800 111.025 20.905 ;
        RECT 12.750 4.510 111.025 4.800 ;
      LAYER met5 ;
        RECT 12.540 4.300 56.460 5.900 ;
  END
END N_term_RAM_IO
END LIBRARY

