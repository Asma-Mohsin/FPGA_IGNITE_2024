module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    VGND,
    VPWR,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 input VGND;
 input VPWR;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire \E6BEG_outbuf_0.A ;
 wire \E6BEG_outbuf_0.X ;
 wire \E6BEG_outbuf_1.A ;
 wire \E6BEG_outbuf_1.X ;
 wire \E6BEG_outbuf_2.A ;
 wire \E6BEG_outbuf_2.X ;
 wire \E6BEG_outbuf_3.A ;
 wire \E6BEG_outbuf_3.X ;
 wire \E6BEG_outbuf_4.A ;
 wire \E6BEG_outbuf_4.X ;
 wire \E6BEG_outbuf_5.A ;
 wire \E6BEG_outbuf_5.X ;
 wire \E6BEG_outbuf_6.A ;
 wire \E6BEG_outbuf_6.X ;
 wire \E6BEG_outbuf_7.A ;
 wire \E6BEG_outbuf_7.X ;
 wire \E6BEG_outbuf_8.A ;
 wire \E6BEG_outbuf_8.X ;
 wire \E6BEG_outbuf_9.A ;
 wire \E6BEG_outbuf_9.X ;
 wire \EE4BEG_outbuf_0.A ;
 wire \EE4BEG_outbuf_0.X ;
 wire \EE4BEG_outbuf_1.A ;
 wire \EE4BEG_outbuf_1.X ;
 wire \EE4BEG_outbuf_10.A ;
 wire \EE4BEG_outbuf_10.X ;
 wire \EE4BEG_outbuf_11.A ;
 wire \EE4BEG_outbuf_11.X ;
 wire \EE4BEG_outbuf_2.A ;
 wire \EE4BEG_outbuf_2.X ;
 wire \EE4BEG_outbuf_3.A ;
 wire \EE4BEG_outbuf_3.X ;
 wire \EE4BEG_outbuf_4.A ;
 wire \EE4BEG_outbuf_4.X ;
 wire \EE4BEG_outbuf_5.A ;
 wire \EE4BEG_outbuf_5.X ;
 wire \EE4BEG_outbuf_6.A ;
 wire \EE4BEG_outbuf_6.X ;
 wire \EE4BEG_outbuf_7.A ;
 wire \EE4BEG_outbuf_7.X ;
 wire \EE4BEG_outbuf_8.A ;
 wire \EE4BEG_outbuf_8.X ;
 wire \EE4BEG_outbuf_9.A ;
 wire \EE4BEG_outbuf_9.X ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.Ci ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.Co ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[0] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[10] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[11] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[12] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[13] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[14] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[15] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[16] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[17] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[18] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[1] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[2] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[3] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[4] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[5] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[6] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[7] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[8] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[9] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.EN ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.I[0] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.I[1] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.I[2] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.I[3] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.LUT_out ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.O ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.SR ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._01_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._02_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._04_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._05_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._06_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._07_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._08_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr._09_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[152] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[153] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[154] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[155] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[156] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[157] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[158] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[159] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[160] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[161] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[162] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[163] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[164] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[165] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[166] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[167] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[168] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[169] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[170] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[171] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[172] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[173] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[174] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[175] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[176] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[177] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[178] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[179] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[180] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[181] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[182] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[183] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[184] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[185] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[186] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[187] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[188] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[189] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[190] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[191] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[192] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[193] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[194] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[195] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[196] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[197] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[198] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[199] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[200] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[201] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[202] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[203] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[204] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[205] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[206] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[207] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[208] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[209] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[210] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[211] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[212] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[213] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[214] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[215] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[216] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[217] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[218] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[219] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[220] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[221] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[222] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[223] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[224] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[225] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[226] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[227] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[228] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[229] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[230] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[231] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[232] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[233] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[234] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[235] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[236] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[237] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[238] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[239] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[240] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[241] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[242] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[243] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[244] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[245] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[246] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[247] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[248] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[249] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[250] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[251] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[252] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[253] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[254] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[255] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[256] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[257] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[258] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[259] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[260] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[261] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[262] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[263] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[264] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[265] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[266] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[267] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[268] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[269] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[270] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[271] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[272] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[273] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[274] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[275] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[276] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[277] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[278] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[279] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[280] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[281] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[282] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[283] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[284] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[285] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[286] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[287] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[288] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[289] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[290] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[291] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[292] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[293] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[294] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[295] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[296] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[297] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[298] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[299] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[300] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[301] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[302] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[303] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[304] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[305] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[306] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[307] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[308] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[309] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[310] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[311] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[312] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[313] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[314] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[315] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[316] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[317] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[318] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[319] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[320] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[321] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[322] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[323] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[324] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[325] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[326] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[327] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[328] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[329] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[330] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[331] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[332] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[333] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[334] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[335] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[336] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[337] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[338] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[339] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[340] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[341] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[342] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[343] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[344] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[345] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[346] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[347] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[348] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[349] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[350] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[351] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[352] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[353] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[354] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[355] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[356] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[357] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[358] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[359] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[360] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[361] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[362] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[363] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[364] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[365] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[366] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[367] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[368] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[369] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[370] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[371] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[372] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[373] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[374] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[375] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[376] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[377] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[378] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[379] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[380] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[381] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[382] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[383] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[384] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[385] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[386] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[387] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[388] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[389] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[390] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[391] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[392] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[393] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[394] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[395] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[396] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[397] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[398] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[399] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[400] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[401] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[402] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[403] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[404] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[405] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[406] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[407] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[408] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[409] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[410] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[411] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[412] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[413] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[414] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[415] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[416] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[417] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[418] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[419] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[420] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[421] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[422] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[423] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[424] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[425] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[426] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[427] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[428] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[429] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[430] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[431] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[432] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[433] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[434] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[435] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[436] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[437] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[438] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[439] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[440] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[441] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[442] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[443] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[444] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[445] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[446] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[447] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[448] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[449] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[450] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[451] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[452] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[453] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[454] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[455] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[456] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[457] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[458] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[459] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[460] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[461] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[462] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[463] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[464] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[465] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[466] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[467] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[468] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[469] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[470] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[471] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[472] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[473] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[474] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[475] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[476] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[477] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[478] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[479] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[480] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[481] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[482] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[483] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[484] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[485] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[486] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[487] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[488] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[489] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[490] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[491] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[492] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[493] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[494] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[495] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[496] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[497] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[498] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[499] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[500] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[501] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[502] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[503] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[504] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[505] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[506] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[507] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[508] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[509] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[510] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[511] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[512] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[513] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[514] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[515] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[516] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[517] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[518] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[519] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[520] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[521] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[522] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[523] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[524] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[525] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[526] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[527] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[528] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[529] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[530] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[531] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[532] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[533] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[534] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[535] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[536] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[537] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[538] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[539] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[540] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[541] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[542] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[543] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[544] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[545] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[546] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[547] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[548] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[549] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[550] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[551] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[552] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[553] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[554] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[555] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[556] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[557] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[558] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[559] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[560] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[561] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[562] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[563] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[564] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[565] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[566] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[567] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[568] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[569] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[570] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[571] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[572] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[573] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[574] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[575] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[576] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[577] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[578] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[579] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[580] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[581] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[582] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[583] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[584] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[585] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[586] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[587] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[588] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[589] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[590] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[591] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[592] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[593] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[594] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[595] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[596] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[597] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[598] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[599] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[600] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[601] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[602] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[603] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[604] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[605] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[606] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[607] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[608] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[609] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[610] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[611] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[612] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[613] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[614] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits[615] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[0] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[100] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[101] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[102] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[103] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[104] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[105] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[106] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[107] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[108] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[109] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[10] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[110] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[111] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[112] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[113] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[114] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[115] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[116] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[117] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[118] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[119] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[11] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[120] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[121] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[122] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[123] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[124] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[125] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[126] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[127] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[128] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[129] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[12] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[130] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[131] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[132] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[133] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[134] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[135] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[136] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[137] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[138] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[139] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[13] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[140] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[141] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[142] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[143] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[144] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[145] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[146] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[147] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[148] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[149] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[14] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[150] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[151] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[152] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[153] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[154] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[155] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[156] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[157] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[158] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[159] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[15] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[160] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[161] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[162] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[163] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[164] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[165] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[166] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[167] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[168] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[169] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[16] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[170] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[171] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[172] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[173] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[174] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[175] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[176] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[177] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[178] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[179] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[17] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[180] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[181] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[182] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[183] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[184] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[185] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[186] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[187] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[188] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[189] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[18] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[190] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[191] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[192] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[193] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[194] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[195] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[196] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[197] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[198] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[199] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[19] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[1] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[200] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[201] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[202] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[203] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[204] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[205] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[206] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[207] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[208] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[209] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[20] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[210] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[211] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[212] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[213] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[214] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[215] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[216] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[217] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[218] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[219] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[21] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[220] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[221] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[222] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[223] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[224] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[225] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[226] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[227] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[228] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[229] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[22] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[230] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[231] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[232] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[233] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[234] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[235] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[236] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[237] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[238] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[239] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[23] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[240] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[241] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[242] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[243] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[244] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[245] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[246] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[247] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[248] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[249] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[24] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[250] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[251] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[252] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[253] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[254] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[255] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[256] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[257] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[258] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[259] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[25] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[260] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[261] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[262] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[263] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[264] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[265] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[266] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[267] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[268] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[269] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[26] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[270] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[271] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[272] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[273] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[274] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[275] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[276] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[277] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[278] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[279] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[27] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[280] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[281] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[282] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[283] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[284] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[285] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[286] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[287] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[288] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[289] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[28] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[290] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[291] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[292] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[293] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[294] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[295] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[296] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[297] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[298] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[299] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[29] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[2] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[300] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[301] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[302] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[303] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[304] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[305] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[306] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[307] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[308] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[309] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[30] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[310] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[311] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[312] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[313] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[314] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[315] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[316] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[317] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[318] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[319] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[31] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[320] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[321] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[322] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[323] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[324] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[325] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[326] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[327] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[328] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[329] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[32] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[330] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[331] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[332] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[333] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[334] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[335] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[336] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[337] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[338] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[339] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[33] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[340] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[341] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[342] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[343] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[344] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[345] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[346] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[347] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[348] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[349] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[34] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[350] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[351] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[352] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[353] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[354] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[355] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[356] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[357] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[358] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[359] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[35] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[360] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[361] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[362] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[363] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[364] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[365] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[366] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[367] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[368] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[369] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[36] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[370] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[371] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[372] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[373] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[374] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[375] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[376] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[377] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[378] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[379] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[37] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[380] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[381] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[382] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[383] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[384] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[385] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[386] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[387] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[388] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[389] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[38] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[390] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[391] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[392] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[393] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[394] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[395] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[396] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[397] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[398] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[399] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[39] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[3] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[400] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[401] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[402] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[403] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[404] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[405] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[406] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[407] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[408] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[409] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[40] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[410] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[411] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[412] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[413] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[414] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[415] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[416] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[417] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[418] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[419] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[41] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[420] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[421] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[422] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[423] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[424] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[425] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[426] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[427] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[428] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[429] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[42] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[430] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[431] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[432] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[433] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[434] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[435] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[436] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[437] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[438] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[439] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[43] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[440] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[441] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[442] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[443] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[444] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[445] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[446] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[447] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[448] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[449] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[44] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[450] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[451] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[452] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[453] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[454] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[455] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[456] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[457] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[458] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[459] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[45] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[460] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[461] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[462] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[463] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[464] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[465] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[466] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[467] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[468] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[469] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[46] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[470] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[471] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[472] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[473] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[474] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[475] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[476] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[477] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[478] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[479] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[47] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[480] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[481] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[482] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[483] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[484] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[485] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[486] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[487] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[488] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[489] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[48] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[490] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[491] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[492] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[493] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[494] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[495] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[496] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[497] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[498] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[499] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[49] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[4] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[500] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[501] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[502] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[503] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[504] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[505] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[506] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[507] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[508] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[509] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[50] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[510] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[511] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[512] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[513] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[514] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[515] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[516] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[517] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[518] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[519] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[51] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[520] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[521] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[522] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[523] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[524] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[525] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[526] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[527] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[528] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[529] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[52] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[530] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[531] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[532] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[533] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[534] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[535] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[536] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[537] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[538] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[539] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[53] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[540] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[541] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[542] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[543] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[544] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[545] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[546] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[547] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[548] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[549] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[54] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[550] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[551] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[552] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[553] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[554] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[555] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[556] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[557] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[558] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[559] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[55] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[560] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[561] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[562] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[563] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[564] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[565] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[566] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[567] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[568] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[569] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[56] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[570] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[571] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[572] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[573] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[574] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[575] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[576] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[577] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[578] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[579] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[57] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[580] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[581] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[582] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[583] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[584] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[585] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[586] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[587] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[588] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[589] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[58] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[590] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[591] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[592] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[593] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[594] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[595] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[596] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[597] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[598] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[599] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[59] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[5] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[600] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[601] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[602] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[603] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[604] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[605] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[606] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[607] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[608] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[609] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[60] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[610] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[611] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[612] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[613] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[614] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[615] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[61] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[62] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[63] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[64] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[65] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[66] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[67] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[68] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[69] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[6] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[70] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[71] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[72] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[73] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[74] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[75] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[76] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[77] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[78] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[79] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[7] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[80] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[81] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[82] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[83] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[84] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[85] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[86] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[87] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[88] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[89] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[8] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[90] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[91] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[92] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[93] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[94] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[95] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[96] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[97] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[98] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[99] ;
 wire \Inst_LUT4AB_ConfigMem.ConfigBits_N[9] ;
 wire \Inst_LUT4AB_switch_matrix.A ;
 wire \Inst_LUT4AB_switch_matrix.B ;
 wire \Inst_LUT4AB_switch_matrix.C ;
 wire \Inst_LUT4AB_switch_matrix.D ;
 wire \Inst_LUT4AB_switch_matrix.E ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb0 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb1 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb2 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb3 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb4 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb5 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb6 ;
 wire \Inst_LUT4AB_switch_matrix.E2BEGb7 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.E6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.EE4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.F ;
 wire \Inst_LUT4AB_switch_matrix.G ;
 wire \Inst_LUT4AB_switch_matrix.H ;
 wire \Inst_LUT4AB_switch_matrix.J2END_AB_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_CD_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_CD_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_CD_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_CD_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_EF_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_EF_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_GH_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_GH_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_GH_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2END_GH_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JE2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JN2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JS2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.JW2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.J_EN_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J_SR_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.M_AB ;
 wire \Inst_LUT4AB_switch_matrix.M_AD ;
 wire \Inst_LUT4AB_switch_matrix.M_AH ;
 wire \Inst_LUT4AB_switch_matrix.M_EF ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb0 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb1 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb2 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb3 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb4 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb5 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb6 ;
 wire \Inst_LUT4AB_switch_matrix.N2BEGb7 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.N4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.NN4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S0 ;
 wire \Inst_LUT4AB_switch_matrix.S1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S2 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb0 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb1 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb2 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb3 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb4 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb5 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb6 ;
 wire \Inst_LUT4AB_switch_matrix.S2BEGb7 ;
 wire \Inst_LUT4AB_switch_matrix.S3 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.S4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.SS4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W1BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG4 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG5 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG6 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEG7 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb0 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb1 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb2 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb3 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb4 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb5 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb6 ;
 wire \Inst_LUT4AB_switch_matrix.W2BEGb7 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.W6BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG0 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG1 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG2 ;
 wire \Inst_LUT4AB_switch_matrix.WW4BEG3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._1_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A0 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A1 ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN[0] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN[1] ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._0_ ;
 wire \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.AD ;
 wire \Inst_MUX8LUT_frame_config_mux.AH ;
 wire \Inst_MUX8LUT_frame_config_mux.CD ;
 wire \Inst_MUX8LUT_frame_config_mux.EH ;
 wire \Inst_MUX8LUT_frame_config_mux.EH_GH ;
 wire \Inst_MUX8LUT_frame_config_mux.GH ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._1_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN[0] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN[1] ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._0_ ;
 wire \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._1_ ;
 wire \N4BEG_outbuf_0.A ;
 wire \N4BEG_outbuf_0.X ;
 wire \N4BEG_outbuf_1.A ;
 wire \N4BEG_outbuf_1.X ;
 wire \N4BEG_outbuf_10.A ;
 wire \N4BEG_outbuf_10.X ;
 wire \N4BEG_outbuf_11.A ;
 wire \N4BEG_outbuf_11.X ;
 wire \N4BEG_outbuf_2.A ;
 wire \N4BEG_outbuf_2.X ;
 wire \N4BEG_outbuf_3.A ;
 wire \N4BEG_outbuf_3.X ;
 wire \N4BEG_outbuf_4.A ;
 wire \N4BEG_outbuf_4.X ;
 wire \N4BEG_outbuf_5.A ;
 wire \N4BEG_outbuf_5.X ;
 wire \N4BEG_outbuf_6.A ;
 wire \N4BEG_outbuf_6.X ;
 wire \N4BEG_outbuf_7.A ;
 wire \N4BEG_outbuf_7.X ;
 wire \N4BEG_outbuf_8.A ;
 wire \N4BEG_outbuf_8.X ;
 wire \N4BEG_outbuf_9.A ;
 wire \N4BEG_outbuf_9.X ;
 wire \NN4BEG_outbuf_0.A ;
 wire \NN4BEG_outbuf_0.X ;
 wire \NN4BEG_outbuf_1.A ;
 wire \NN4BEG_outbuf_1.X ;
 wire \NN4BEG_outbuf_10.A ;
 wire \NN4BEG_outbuf_10.X ;
 wire \NN4BEG_outbuf_11.A ;
 wire \NN4BEG_outbuf_11.X ;
 wire \NN4BEG_outbuf_2.A ;
 wire \NN4BEG_outbuf_2.X ;
 wire \NN4BEG_outbuf_3.A ;
 wire \NN4BEG_outbuf_3.X ;
 wire \NN4BEG_outbuf_4.A ;
 wire \NN4BEG_outbuf_4.X ;
 wire \NN4BEG_outbuf_5.A ;
 wire \NN4BEG_outbuf_5.X ;
 wire \NN4BEG_outbuf_6.A ;
 wire \NN4BEG_outbuf_6.X ;
 wire \NN4BEG_outbuf_7.A ;
 wire \NN4BEG_outbuf_7.X ;
 wire \NN4BEG_outbuf_8.A ;
 wire \NN4BEG_outbuf_8.X ;
 wire \NN4BEG_outbuf_9.A ;
 wire \NN4BEG_outbuf_9.X ;
 wire \S4BEG_outbuf_0.A ;
 wire \S4BEG_outbuf_0.X ;
 wire \S4BEG_outbuf_1.A ;
 wire \S4BEG_outbuf_1.X ;
 wire \S4BEG_outbuf_10.A ;
 wire \S4BEG_outbuf_10.X ;
 wire \S4BEG_outbuf_11.A ;
 wire \S4BEG_outbuf_11.X ;
 wire \S4BEG_outbuf_2.A ;
 wire \S4BEG_outbuf_2.X ;
 wire \S4BEG_outbuf_3.A ;
 wire \S4BEG_outbuf_3.X ;
 wire \S4BEG_outbuf_4.A ;
 wire \S4BEG_outbuf_4.X ;
 wire \S4BEG_outbuf_5.A ;
 wire \S4BEG_outbuf_5.X ;
 wire \S4BEG_outbuf_6.A ;
 wire \S4BEG_outbuf_6.X ;
 wire \S4BEG_outbuf_7.A ;
 wire \S4BEG_outbuf_7.X ;
 wire \S4BEG_outbuf_8.A ;
 wire \S4BEG_outbuf_8.X ;
 wire \S4BEG_outbuf_9.A ;
 wire \S4BEG_outbuf_9.X ;
 wire \SS4BEG_outbuf_0.A ;
 wire \SS4BEG_outbuf_0.X ;
 wire \SS4BEG_outbuf_1.A ;
 wire \SS4BEG_outbuf_1.X ;
 wire \SS4BEG_outbuf_10.A ;
 wire \SS4BEG_outbuf_10.X ;
 wire \SS4BEG_outbuf_11.A ;
 wire \SS4BEG_outbuf_11.X ;
 wire \SS4BEG_outbuf_2.A ;
 wire \SS4BEG_outbuf_2.X ;
 wire \SS4BEG_outbuf_3.A ;
 wire \SS4BEG_outbuf_3.X ;
 wire \SS4BEG_outbuf_4.A ;
 wire \SS4BEG_outbuf_4.X ;
 wire \SS4BEG_outbuf_5.A ;
 wire \SS4BEG_outbuf_5.X ;
 wire \SS4BEG_outbuf_6.A ;
 wire \SS4BEG_outbuf_6.X ;
 wire \SS4BEG_outbuf_7.A ;
 wire \SS4BEG_outbuf_7.X ;
 wire \SS4BEG_outbuf_8.A ;
 wire \SS4BEG_outbuf_8.X ;
 wire \SS4BEG_outbuf_9.A ;
 wire \SS4BEG_outbuf_9.X ;
 wire \W6BEG_outbuf_0.A ;
 wire \W6BEG_outbuf_0.X ;
 wire \W6BEG_outbuf_1.A ;
 wire \W6BEG_outbuf_1.X ;
 wire \W6BEG_outbuf_2.A ;
 wire \W6BEG_outbuf_2.X ;
 wire \W6BEG_outbuf_3.A ;
 wire \W6BEG_outbuf_3.X ;
 wire \W6BEG_outbuf_4.A ;
 wire \W6BEG_outbuf_4.X ;
 wire \W6BEG_outbuf_5.A ;
 wire \W6BEG_outbuf_5.X ;
 wire \W6BEG_outbuf_6.A ;
 wire \W6BEG_outbuf_6.X ;
 wire \W6BEG_outbuf_7.A ;
 wire \W6BEG_outbuf_7.X ;
 wire \W6BEG_outbuf_8.A ;
 wire \W6BEG_outbuf_8.X ;
 wire \W6BEG_outbuf_9.A ;
 wire \W6BEG_outbuf_9.X ;
 wire \WW4BEG_outbuf_0.A ;
 wire \WW4BEG_outbuf_0.X ;
 wire \WW4BEG_outbuf_1.A ;
 wire \WW4BEG_outbuf_1.X ;
 wire \WW4BEG_outbuf_10.A ;
 wire \WW4BEG_outbuf_10.X ;
 wire \WW4BEG_outbuf_11.A ;
 wire \WW4BEG_outbuf_11.X ;
 wire \WW4BEG_outbuf_2.A ;
 wire \WW4BEG_outbuf_2.X ;
 wire \WW4BEG_outbuf_3.A ;
 wire \WW4BEG_outbuf_3.X ;
 wire \WW4BEG_outbuf_4.A ;
 wire \WW4BEG_outbuf_4.X ;
 wire \WW4BEG_outbuf_5.A ;
 wire \WW4BEG_outbuf_5.X ;
 wire \WW4BEG_outbuf_6.A ;
 wire \WW4BEG_outbuf_6.X ;
 wire \WW4BEG_outbuf_7.A ;
 wire \WW4BEG_outbuf_7.X ;
 wire \WW4BEG_outbuf_8.A ;
 wire \WW4BEG_outbuf_8.X ;
 wire \WW4BEG_outbuf_9.A ;
 wire \WW4BEG_outbuf_9.X ;
 wire \data_inbuf_0.X ;
 wire \data_inbuf_1.X ;
 wire \data_inbuf_10.X ;
 wire \data_inbuf_11.X ;
 wire \data_inbuf_12.X ;
 wire \data_inbuf_13.X ;
 wire \data_inbuf_14.X ;
 wire \data_inbuf_15.X ;
 wire \data_inbuf_16.X ;
 wire \data_inbuf_17.X ;
 wire \data_inbuf_18.X ;
 wire \data_inbuf_19.X ;
 wire \data_inbuf_2.X ;
 wire \data_inbuf_20.X ;
 wire \data_inbuf_21.X ;
 wire \data_inbuf_22.X ;
 wire \data_inbuf_23.X ;
 wire \data_inbuf_24.X ;
 wire \data_inbuf_25.X ;
 wire \data_inbuf_26.X ;
 wire \data_inbuf_27.X ;
 wire \data_inbuf_28.X ;
 wire \data_inbuf_29.X ;
 wire \data_inbuf_3.X ;
 wire \data_inbuf_30.X ;
 wire \data_inbuf_31.X ;
 wire \data_inbuf_4.X ;
 wire \data_inbuf_5.X ;
 wire \data_inbuf_6.X ;
 wire \data_inbuf_7.X ;
 wire \data_inbuf_8.X ;
 wire \data_inbuf_9.X ;
 wire \data_outbuf_0.X ;
 wire \data_outbuf_1.X ;
 wire \data_outbuf_10.X ;
 wire \data_outbuf_11.X ;
 wire \data_outbuf_12.X ;
 wire \data_outbuf_13.X ;
 wire \data_outbuf_14.X ;
 wire \data_outbuf_15.X ;
 wire \data_outbuf_16.X ;
 wire \data_outbuf_17.X ;
 wire \data_outbuf_18.X ;
 wire \data_outbuf_19.X ;
 wire \data_outbuf_2.X ;
 wire \data_outbuf_20.X ;
 wire \data_outbuf_21.X ;
 wire \data_outbuf_22.X ;
 wire \data_outbuf_23.X ;
 wire \data_outbuf_24.X ;
 wire \data_outbuf_25.X ;
 wire \data_outbuf_26.X ;
 wire \data_outbuf_27.X ;
 wire \data_outbuf_28.X ;
 wire \data_outbuf_29.X ;
 wire \data_outbuf_3.X ;
 wire \data_outbuf_30.X ;
 wire \data_outbuf_31.X ;
 wire \data_outbuf_4.X ;
 wire \data_outbuf_5.X ;
 wire \data_outbuf_6.X ;
 wire \data_outbuf_7.X ;
 wire \data_outbuf_8.X ;
 wire \data_outbuf_9.X ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \strobe_inbuf_0.X ;
 wire \strobe_inbuf_1.X ;
 wire \strobe_inbuf_10.X ;
 wire \strobe_inbuf_11.X ;
 wire \strobe_inbuf_12.X ;
 wire \strobe_inbuf_13.X ;
 wire \strobe_inbuf_14.X ;
 wire \strobe_inbuf_15.X ;
 wire \strobe_inbuf_16.X ;
 wire \strobe_inbuf_17.X ;
 wire \strobe_inbuf_18.X ;
 wire \strobe_inbuf_19.X ;
 wire \strobe_inbuf_2.X ;
 wire \strobe_inbuf_3.X ;
 wire \strobe_inbuf_4.X ;
 wire \strobe_inbuf_5.X ;
 wire \strobe_inbuf_6.X ;
 wire \strobe_inbuf_7.X ;
 wire \strobe_inbuf_8.X ;
 wire \strobe_inbuf_9.X ;
 wire \strobe_outbuf_0.X ;
 wire \strobe_outbuf_1.X ;
 wire \strobe_outbuf_10.X ;
 wire \strobe_outbuf_11.X ;
 wire \strobe_outbuf_12.X ;
 wire \strobe_outbuf_13.X ;
 wire \strobe_outbuf_14.X ;
 wire \strobe_outbuf_15.X ;
 wire \strobe_outbuf_16.X ;
 wire \strobe_outbuf_17.X ;
 wire \strobe_outbuf_18.X ;
 wire \strobe_outbuf_19.X ;
 wire \strobe_outbuf_2.X ;
 wire \strobe_outbuf_3.X ;
 wire \strobe_outbuf_4.X ;
 wire \strobe_outbuf_5.X ;
 wire \strobe_outbuf_6.X ;
 wire \strobe_outbuf_7.X ;
 wire \strobe_outbuf_8.X ;
 wire \strobe_outbuf_9.X ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\E6BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\EE4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\EE4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\SS4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\W6BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\EE4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\EE4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(\EE4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\W6BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\WW4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\E6BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\E6BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\Inst_LUT4AB_switch_matrix.N2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\Inst_LUT4AB_switch_matrix.N2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\N4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\N4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\N4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\N4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\E6BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\N4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\NN4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\NN4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\NN4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\NN4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\NN4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\NN4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\NN4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\S4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\S4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\EE4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\S4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\S4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\S4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\SS4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\SS4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\SS4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\SS4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\SS4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\W6BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\W6BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\EE4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\W6BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\WW4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\WW4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\WW4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\WW4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net6),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net539),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\E6BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\EE4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\EE4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\Inst_LUT4AB_switch_matrix.W2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\NN4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\NN4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\NN4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\S4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\SS4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\W6BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_0._0_  (.A(\E6BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_1._0_  (.A(\E6BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_2._0_  (.A(\E6BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_3._0_  (.A(\E6BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_4._0_  (.A(\E6BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_5._0_  (.A(\E6BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_6._0_  (.A(\E6BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_7._0_  (.A(\E6BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_8._0_  (.A(\E6BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_9._0_  (.A(\E6BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_0._0_  (.A(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_1._0_  (.A(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_2._0_  (.A(net28),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_3._0_  (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_4._0_  (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_5._0_  (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_6._0_  (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_7._0_  (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_8._0_  (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_9._0_  (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\E6BEG_outbuf_9.A ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_0._0_  (.A(\EE4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_1._0_  (.A(\EE4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_10._0_  (.A(\EE4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_11._0_  (.A(\EE4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_2._0_  (.A(\EE4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_3._0_  (.A(\EE4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_4._0_  (.A(\EE4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_5._0_  (.A(\EE4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_6._0_  (.A(\EE4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_7._0_  (.A(\EE4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_8._0_  (.A(\EE4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_9._0_  (.A(\EE4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_0._0_  (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_1._0_  (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_10._0_  (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_11._0_  (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_2._0_  (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_3._0_  (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_4._0_  (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_5._0_  (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_6._0_  (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_7._0_  (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_8._0_  (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_9._0_  (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\EE4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_34_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_34_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_34_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_452 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_35_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_35_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_36_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_37_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_38_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_39_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_39_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_40_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_40_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_41_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_203 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_44_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_45_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_45_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_373 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_256 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_48_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_49_348 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_49_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_383 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_50_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_403 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_50_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_51_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_368 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_52_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_369 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_52_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_438 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_53_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_198 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_53_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_54_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_55_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_55_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_56_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_57_263 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_57_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_57_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_58_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_59_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_59_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_60_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_61_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_61_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_62_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_62_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_430 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_254 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_63_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_63_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_63_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_258 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_310 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_69_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_69_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_70_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_71_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_246 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_72_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_408 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_216 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_358 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_370 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_352 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_439 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_450 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_247 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_424 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_77_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LA_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LA_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LA_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LA_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LA_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LA_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LA_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LA_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LA_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LA_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LA_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LA_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LA_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LA_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LA_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LA_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LB_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LB_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LB_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LB_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LB_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LB_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LB_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LB_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LB_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LB_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LB_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LB_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LB_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LB_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LB_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LB_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LC_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LC_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LC_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LC_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LC_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LC_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LC_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LC_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LC_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LC_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LC_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LC_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LC_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LC_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LC_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LC_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LD_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LD_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LD_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LD_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LD_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LD_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LD_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LD_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LD_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LD_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LD_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LD_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LD_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LD_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LD_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LD_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LE_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LE_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LE_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LE_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LE_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LE_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LE_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LE_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LE_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LE_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LE_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LE_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LE_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LF_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_2 \Inst_LF_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LF_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LF_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LF_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LF_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LF_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LF_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LF_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LF_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LF_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LF_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LF_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LG_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LG_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LG_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LG_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LG_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LG_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LG_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LG_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LG_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LG_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LG_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LG_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LG_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LG_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LG_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LG_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr._11_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr._12_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.I[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._02_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LH_LUT4c_frame_config_dffesr._14_  (.A1(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.I[2] ),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._05_ ));
 sky130_fd_sc_hd__a21oi_1 \Inst_LH_LUT4c_frame_config_dffesr._15_  (.A1(\Inst_LH_LUT4c_frame_config_dffesr._01_ ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr._02_ ),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr._05_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.Co ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr._16_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._06_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr._17_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._07_ ));
 sky130_fd_sc_hd__or2b_1 \Inst_LH_LUT4c_frame_config_dffesr._18_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.SR ),
    .B_N(\Inst_LH_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr._08_ ));
 sky130_fd_sc_hd__a21boi_1 \Inst_LH_LUT4c_frame_config_dffesr._19_  (.A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.SR ),
    .B1_N(\Inst_LH_LUT4c_frame_config_dffesr.EN ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._09_ ));
 sky130_fd_sc_hd__a22oi_1 \Inst_LH_LUT4c_frame_config_dffesr._20_  (.A1(\Inst_LH_LUT4c_frame_config_dffesr._06_ ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr._07_ ),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr._08_ ),
    .B2(\Inst_LH_LUT4c_frame_config_dffesr._09_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr._04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LH_LUT4c_frame_config_dffesr._21_  (.CLK(UserCLK),
    .D(\Inst_LH_LUT4c_frame_config_dffesr._04_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ),
    .B(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_  (.A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ ),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.I0mux ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.I[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.Ci ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._2_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._3_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ),
    .B(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._4_  (.A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._0_ ),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_out ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.LUT_flop ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr.I0mux ),
    .S1(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr.I[2] ),
    .S1(\Inst_LH_LUT4c_frame_config_dffesr.I[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.LUT_out ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit0  (.D(net50),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[389] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit1  (.D(net61),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[397] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit10  (.D(net51),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[577] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[577] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit11  (.D(net52),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[576] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[576] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit12  (.D(net53),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[568] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[568] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit13  (.D(net54),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[159] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit14  (.D(net55),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[158] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit15  (.D(net56),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[157] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit16  (.D(net57),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[241] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit17  (.D(net58),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[240] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit18  (.D(net59),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[263] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit19  (.D(net60),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[261] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit20  (.D(net62),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[259] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit21  (.D(net63),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[248] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit22  (.D(net64),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[247] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit23  (.D(net65),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[243] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit24  (.D(net66),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[242] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit3  (.D(net75),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[413] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[413] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit4  (.D(net76),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[462] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[462] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit5  (.D(net77),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[481] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[481] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit6  (.D(net78),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[473] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[473] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit7  (.D(net79),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[472] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[472] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit8  (.D(net80),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[502] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[502] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame0_bit9  (.D(net81),
    .GATE(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[558] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[558] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit0  (.D(net50),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[330] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit1  (.D(net61),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[338] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit10  (.D(net51),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[395] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit11  (.D(net52),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[411] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[411] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit12  (.D(net53),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[557] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[557] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit13  (.D(net54),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[581] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[581] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit14  (.D(net55),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit15  (.D(net56),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit16  (.D(net57),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit17  (.D(net58),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit18  (.D(net59),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit19  (.D(net60),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit2  (.D(net72),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[391] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit20  (.D(net62),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit21  (.D(net63),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[199] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit22  (.D(net64),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[196] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit23  (.D(net65),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[222] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit24  (.D(net66),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[221] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit25  (.D(net67),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[220] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit26  (.D(net68),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[200] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit27  (.D(net69),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[232] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit28  (.D(net70),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[271] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit29  (.D(net71),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[270] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit3  (.D(net75),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[390] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit30  (.D(net73),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[615] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[615] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit31  (.D(net74),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[601] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[601] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit4  (.D(net76),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[381] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit5  (.D(net77),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[380] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit6  (.D(net78),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[377] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit7  (.D(net79),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[376] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit8  (.D(net80),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[360] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame10_bit9  (.D(net81),
    .GATE(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[398] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit0  (.D(net50),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[322] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit1  (.D(net61),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[318] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit10  (.D(net51),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[416] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[416] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit11  (.D(net52),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[394] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit12  (.D(net53),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[410] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[410] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit13  (.D(net54),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[403] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit14  (.D(net55),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[521] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[521] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit15  (.D(net56),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit16  (.D(net57),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit17  (.D(net58),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit18  (.D(net59),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit19  (.D(net60),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit2  (.D(net72),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[296] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit20  (.D(net62),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit21  (.D(net63),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit22  (.D(net64),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[198] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit23  (.D(net65),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[188] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit24  (.D(net66),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[187] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit25  (.D(net67),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[201] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit26  (.D(net68),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[234] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit27  (.D(net69),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[233] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit28  (.D(net70),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[610] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[610] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit29  (.D(net71),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[602] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[602] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit3  (.D(net75),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[332] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit30  (.D(net73),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[585] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[585] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit31  (.D(net74),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[584] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[584] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit4  (.D(net76),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[331] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit5  (.D(net77),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[355] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit6  (.D(net78),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[339] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit7  (.D(net79),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[387] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit8  (.D(net80),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[400] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame11_bit9  (.D(net81),
    .GATE(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[417] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[417] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit0  (.D(net50),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[327] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit1  (.D(net61),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[297] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit10  (.D(net51),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit11  (.D(net52),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit12  (.D(net53),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit13  (.D(net54),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit14  (.D(net55),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit15  (.D(net56),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit16  (.D(net57),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit17  (.D(net58),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit18  (.D(net59),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit19  (.D(net60),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit2  (.D(net72),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[337] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit20  (.D(net62),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[191] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit21  (.D(net63),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[227] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit22  (.D(net64),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[225] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit23  (.D(net65),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[224] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit24  (.D(net66),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[223] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit25  (.D(net67),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[269] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit26  (.D(net68),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[266] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit27  (.D(net69),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[593] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[593] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit28  (.D(net70),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[587] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[587] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit29  (.D(net71),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[612] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[612] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit3  (.D(net75),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[333] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit30  (.D(net73),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[586] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[586] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit31  (.D(net74),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[594] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[594] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit4  (.D(net76),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[342] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit5  (.D(net77),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[362] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit6  (.D(net78),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[372] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit7  (.D(net79),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[401] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit8  (.D(net80),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[408] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[408] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame12_bit9  (.D(net81),
    .GATE(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[392] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit0  (.D(net50),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[302] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit1  (.D(net61),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[326] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit10  (.D(net51),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[406] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[406] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit11  (.D(net52),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[393] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit12  (.D(net53),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit13  (.D(net54),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit14  (.D(net55),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit15  (.D(net56),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit16  (.D(net57),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit17  (.D(net58),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit18  (.D(net59),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit19  (.D(net60),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit2  (.D(net72),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[321] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit20  (.D(net62),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[190] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit21  (.D(net63),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[189] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit22  (.D(net64),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[226] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit23  (.D(net65),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[267] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit24  (.D(net66),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[288] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit25  (.D(net67),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[287] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit26  (.D(net68),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[277] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit27  (.D(net69),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[276] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit28  (.D(net70),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[592] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[592] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit29  (.D(net71),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[613] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[613] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit3  (.D(net75),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[313] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit30  (.D(net73),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[611] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[611] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit31  (.D(net74),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[595] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[595] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit4  (.D(net76),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[306] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit5  (.D(net77),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[343] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit6  (.D(net78),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[365] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit7  (.D(net79),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[373] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit8  (.D(net80),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[409] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[409] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame13_bit9  (.D(net81),
    .GATE(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[407] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[407] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit0  (.D(net50),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[305] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit1  (.D(net61),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[303] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit10  (.D(net51),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[357] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit11  (.D(net52),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[356] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit12  (.D(net53),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[344] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit13  (.D(net54),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[364] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit14  (.D(net55),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[399] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit15  (.D(net56),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit16  (.D(net57),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit17  (.D(net58),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit18  (.D(net59),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit19  (.D(net60),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit2  (.D(net72),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[323] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit20  (.D(net62),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit21  (.D(net63),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit22  (.D(net64),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit23  (.D(net65),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[192] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit24  (.D(net66),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[183] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit25  (.D(net67),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[182] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit26  (.D(net68),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[228] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit27  (.D(net69),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[272] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit28  (.D(net70),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[293] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit29  (.D(net71),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[291] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit3  (.D(net75),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[320] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit30  (.D(net73),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[278] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit31  (.D(net74),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[614] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[614] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit4  (.D(net76),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[316] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit5  (.D(net77),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[312] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit6  (.D(net78),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[310] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit7  (.D(net79),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[308] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit8  (.D(net80),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[307] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame14_bit9  (.D(net81),
    .GATE(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[334] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit0  (.D(net50),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[301] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit1  (.D(net61),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[300] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit10  (.D(net51),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit11  (.D(net52),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit12  (.D(net53),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit13  (.D(net54),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit14  (.D(net55),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit15  (.D(net56),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit16  (.D(net57),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit17  (.D(net58),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit18  (.D(net59),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit19  (.D(net60),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit2  (.D(net72),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[319] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit20  (.D(net62),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit21  (.D(net63),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit22  (.D(net64),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit23  (.D(net65),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit24  (.D(net66),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit25  (.D(net67),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit26  (.D(net68),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[273] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit27  (.D(net69),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[268] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit28  (.D(net70),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[289] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit29  (.D(net71),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[282] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit3  (.D(net75),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[317] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit30  (.D(net73),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[279] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit31  (.D(net74),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[275] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit4  (.D(net76),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[298] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit5  (.D(net77),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[309] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit6  (.D(net78),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit7  (.D(net79),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit8  (.D(net80),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame15_bit9  (.D(net81),
    .GATE(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit0  (.D(net50),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[335] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit1  (.D(net61),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[345] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit10  (.D(net51),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit11  (.D(net52),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit12  (.D(net53),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit13  (.D(net54),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit14  (.D(net55),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit15  (.D(net56),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit16  (.D(net57),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit17  (.D(net58),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit18  (.D(net59),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit19  (.D(net60),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit2  (.D(net72),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit20  (.D(net62),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit21  (.D(net63),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit22  (.D(net64),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit23  (.D(net65),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit24  (.D(net66),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit25  (.D(net67),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit26  (.D(net68),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit27  (.D(net69),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit28  (.D(net70),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit29  (.D(net71),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit3  (.D(net75),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[17] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit30  (.D(net73),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[283] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit31  (.D(net74),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[274] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit4  (.D(net76),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit5  (.D(net77),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit6  (.D(net78),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit7  (.D(net79),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit8  (.D(net80),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame16_bit9  (.D(net81),
    .GATE(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit0  (.D(net50),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[304] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit1  (.D(net61),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[299] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit10  (.D(net51),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit11  (.D(net52),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit12  (.D(net53),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit13  (.D(net54),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit14  (.D(net55),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit15  (.D(net56),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit16  (.D(net57),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit17  (.D(net58),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit18  (.D(net59),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit19  (.D(net60),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit2  (.D(net72),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[325] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit20  (.D(net62),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit21  (.D(net63),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit22  (.D(net64),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit23  (.D(net65),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit24  (.D(net66),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit25  (.D(net67),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit26  (.D(net68),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[6] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit27  (.D(net69),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit28  (.D(net70),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit29  (.D(net71),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit3  (.D(net75),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit30  (.D(net73),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[295] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit31  (.D(net74),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[285] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit4  (.D(net76),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit5  (.D(net77),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[2] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit6  (.D(net78),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[1] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit7  (.D(net79),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[0] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit8  (.D(net80),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame17_bit9  (.D(net81),
    .GATE(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit0  (.D(net50),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[324] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit1  (.D(net61),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[315] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit10  (.D(net51),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit11  (.D(net52),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit12  (.D(net53),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit13  (.D(net54),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit14  (.D(net55),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit15  (.D(net56),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit16  (.D(net57),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit17  (.D(net58),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit18  (.D(net59),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit19  (.D(net60),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit2  (.D(net72),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[314] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit20  (.D(net62),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit21  (.D(net63),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit22  (.D(net64),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit23  (.D(net65),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit24  (.D(net66),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit25  (.D(net67),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit26  (.D(net68),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit27  (.D(net69),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[9] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit28  (.D(net70),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr.ConfigBits[8] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit29  (.D(net71),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[16] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit3  (.D(net75),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit30  (.D(net73),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[294] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit31  (.D(net74),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[284] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit4  (.D(net76),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[14] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit5  (.D(net77),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit6  (.D(net78),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit7  (.D(net79),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit8  (.D(net80),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[18] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame18_bit9  (.D(net81),
    .GATE(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit10  (.D(net51),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[467] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[467] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit11  (.D(net52),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[575] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[575] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit12  (.D(net53),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[574] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[574] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit13  (.D(net54),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[567] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[567] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit14  (.D(net55),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[566] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[566] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit15  (.D(net56),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[562] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[562] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit16  (.D(net57),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[156] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit17  (.D(net58),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[155] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit18  (.D(net59),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[154] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit19  (.D(net60),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[239] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit2  (.D(net72),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[396] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit20  (.D(net62),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[238] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit21  (.D(net63),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[258] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit22  (.D(net64),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[254] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit23  (.D(net65),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[253] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit24  (.D(net66),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[252] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit25  (.D(net67),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[246] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit3  (.D(net75),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[412] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[412] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit4  (.D(net76),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[405] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit5  (.D(net77),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[404] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit6  (.D(net78),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[479] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[479] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit7  (.D(net79),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[478] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[478] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit8  (.D(net80),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[471] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[471] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame19_bit9  (.D(net81),
    .GATE(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[470] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[470] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit10  (.D(net51),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[526] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[526] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit11  (.D(net52),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[543] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[543] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit12  (.D(net53),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[542] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[542] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit13  (.D(net54),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[537] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[537] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit14  (.D(net55),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[534] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[534] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit15  (.D(net56),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[530] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[530] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit16  (.D(net57),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[560] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[560] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit17  (.D(net58),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[559] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[559] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit18  (.D(net59),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[578] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[578] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit19  (.D(net60),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[573] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[573] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit2  (.D(net72),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[388] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit20  (.D(net62),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[572] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[572] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit21  (.D(net63),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[571] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[571] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit22  (.D(net64),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[570] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[570] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit23  (.D(net65),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[569] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[569] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit24  (.D(net66),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[565] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[565] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit25  (.D(net67),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[563] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[563] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit26  (.D(net68),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[262] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit27  (.D(net69),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[260] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit28  (.D(net70),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[256] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit29  (.D(net71),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[255] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit3  (.D(net75),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[386] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit30  (.D(net73),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[250] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit31  (.D(net74),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[249] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit4  (.D(net76),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[422] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[422] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit5  (.D(net77),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[463] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[463] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit7  (.D(net79),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[480] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[480] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit8  (.D(net80),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[504] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[504] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame1_bit9  (.D(net81),
    .GATE(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[527] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[527] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit1  (.D(net61),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[348] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit10  (.D(net51),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[483] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[483] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit11  (.D(net52),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[475] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[475] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit12  (.D(net53),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[474] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[474] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit13  (.D(net54),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[494] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[494] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit14  (.D(net55),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[503] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[503] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit15  (.D(net56),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[499] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[499] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit16  (.D(net57),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[498] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[498] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit17  (.D(net58),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[529] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[529] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit18  (.D(net59),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[528] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[528] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit19  (.D(net60),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[544] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[544] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit20  (.D(net62),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[536] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[536] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit21  (.D(net63),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[535] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[535] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit22  (.D(net64),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[531] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[531] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit23  (.D(net65),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[561] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[561] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit24  (.D(net66),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[564] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[564] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit25  (.D(net67),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[167] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit26  (.D(net68),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[163] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit27  (.D(net69),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[257] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit28  (.D(net70),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[251] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit30  (.D(net73),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[265] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit31  (.D(net74),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[264] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit4  (.D(net76),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[366] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit5  (.D(net77),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[374] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit6  (.D(net78),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[423] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[423] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit7  (.D(net79),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[439] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[439] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit8  (.D(net80),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[464] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[464] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame2_bit9  (.D(net81),
    .GATE(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[461] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[461] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit1  (.D(net61),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[336] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit10  (.D(net51),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[438] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[438] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit11  (.D(net52),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[465] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[465] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit12  (.D(net53),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[477] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[477] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit13  (.D(net54),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[476] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[476] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit14  (.D(net55),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[497] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[497] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit15  (.D(net56),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[496] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[496] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit16  (.D(net57),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[495] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[495] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit17  (.D(net58),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[491] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[491] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit18  (.D(net59),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[505] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[505] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit19  (.D(net60),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[501] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[501] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit2  (.D(net72),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[353] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit20  (.D(net62),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[500] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[500] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit21  (.D(net63),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[547] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[547] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit22  (.D(net64),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[546] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[546] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit23  (.D(net65),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[545] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[545] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit24  (.D(net66),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[533] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[533] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit25  (.D(net67),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[10] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit26  (.D(net68),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[166] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit27  (.D(net69),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[164] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit28  (.D(net70),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[162] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit29  (.D(net71),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit3  (.D(net75),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[349] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit30  (.D(net73),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[186] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit31  (.D(net74),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[168] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit4  (.D(net76),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[367] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit5  (.D(net77),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[431] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[431] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit6  (.D(net78),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[430] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[430] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit7  (.D(net79),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[451] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[451] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit8  (.D(net80),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[450] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[450] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame3_bit9  (.D(net81),
    .GATE(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[446] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[446] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit0  (.D(net50),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[358] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit1  (.D(net61),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[352] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit10  (.D(net51),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[486] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[486] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit11  (.D(net52),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[482] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[482] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit12  (.D(net53),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[469] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[469] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit13  (.D(net54),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[468] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[468] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit14  (.D(net55),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[466] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[466] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit15  (.D(net56),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[517] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[517] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit16  (.D(net57),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[515] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[515] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit17  (.D(net58),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[514] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[514] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit18  (.D(net59),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[509] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[509] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit19  (.D(net60),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[489] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[489] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit2  (.D(net72),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[363] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit20  (.D(net62),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[550] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[550] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit21  (.D(net63),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[549] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[549] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit22  (.D(net64),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[532] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[532] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit23  (.D(net65),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[165] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit24  (.D(net66),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit25  (.D(net67),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[176] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit26  (.D(net68),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[184] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit27  (.D(net69),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[179] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit28  (.D(net70),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[169] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit29  (.D(net71),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[203] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit3  (.D(net75),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[375] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit30  (.D(net73),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[216] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit31  (.D(net74),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[604] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[604] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit4  (.D(net76),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[371] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit5  (.D(net77),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[370] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit6  (.D(net78),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[428] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[428] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit7  (.D(net79),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[455] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[455] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit8  (.D(net80),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[452] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[452] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame4_bit9  (.D(net81),
    .GATE(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[447] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[447] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit0  (.D(net50),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[359] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit1  (.D(net61),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[346] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit10  (.D(net51),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[437] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[437] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit11  (.D(net52),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[436] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[436] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit12  (.D(net53),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[458] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[458] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit13  (.D(net54),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[457] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[457] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit14  (.D(net55),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[516] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[516] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit15  (.D(net56),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[511] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[511] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit16  (.D(net57),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[510] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[510] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit17  (.D(net58),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[506] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[506] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit18  (.D(net59),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[551] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[551] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit19  (.D(net60),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[548] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[548] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit2  (.D(net72),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[421] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[421] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit20  (.D(net62),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[12] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit21  (.D(net63),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[177] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit22  (.D(net64),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[175] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit23  (.D(net65),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[174] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit24  (.D(net66),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[173] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit25  (.D(net67),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[185] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit26  (.D(net68),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[178] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit27  (.D(net69),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[205] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit28  (.D(net70),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[229] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit29  (.D(net71),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[202] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit3  (.D(net75),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[429] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[429] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit30  (.D(net73),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[210] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit31  (.D(net74),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[589] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[589] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit4  (.D(net76),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[454] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[454] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit5  (.D(net77),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[453] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[453] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit6  (.D(net78),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[448] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[448] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit7  (.D(net79),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[444] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[444] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit8  (.D(net80),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[441] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[441] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame5_bit9  (.D(net81),
    .GATE(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[440] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[440] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit0  (.D(net50),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[311] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit1  (.D(net61),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[347] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit10  (.D(net51),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[484] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[484] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit11  (.D(net52),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[456] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[456] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit12  (.D(net53),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[492] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[492] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit13  (.D(net54),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[513] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[513] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit14  (.D(net55),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[490] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[490] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit15  (.D(net56),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[507] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[507] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit16  (.D(net57),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[553] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[553] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit17  (.D(net58),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr.ConfigBits[11] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit18  (.D(net59),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit19  (.D(net60),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[5] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit2  (.D(net72),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[420] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[420] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit20  (.D(net62),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[170] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit21  (.D(net63),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[181] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit22  (.D(net64),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[208] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit23  (.D(net65),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[206] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit24  (.D(net66),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[204] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit25  (.D(net67),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[231] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit26  (.D(net68),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[214] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit27  (.D(net69),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[213] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit28  (.D(net70),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[212] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit29  (.D(net71),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[211] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit3  (.D(net75),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[433] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[433] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit30  (.D(net73),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[606] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[606] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit31  (.D(net74),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[605] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[605] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit4  (.D(net76),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[449] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[449] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit5  (.D(net77),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[425] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[425] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit6  (.D(net78),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[424] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[424] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit7  (.D(net79),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[487] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[487] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit8  (.D(net80),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[459] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[459] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame6_bit9  (.D(net81),
    .GATE(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[485] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[485] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit0  (.D(net50),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[340] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit1  (.D(net61),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[385] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit10  (.D(net51),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[512] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[512] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit11  (.D(net52),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[508] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[508] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit12  (.D(net53),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[488] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[488] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit13  (.D(net54),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[540] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[540] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit14  (.D(net55),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[522] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[522] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit15  (.D(net56),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[582] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[582] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit16  (.D(net57),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[555] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[555] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit17  (.D(net58),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[552] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[552] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit18  (.D(net59),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[7] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit19  (.D(net60),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[160] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit2  (.D(net72),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[415] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[415] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit20  (.D(net62),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[13] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit21  (.D(net63),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[172] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit22  (.D(net64),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[171] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit23  (.D(net65),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[180] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit24  (.D(net66),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[217] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit25  (.D(net67),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[236] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit26  (.D(net68),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[280] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit27  (.D(net69),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[590] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[590] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit28  (.D(net70),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[588] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[588] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit29  (.D(net71),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[609] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[609] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit3  (.D(net75),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[402] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit30  (.D(net73),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[608] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[608] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit31  (.D(net74),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[596] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[596] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit4  (.D(net76),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[442] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[442] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit5  (.D(net77),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[435] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[435] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit6  (.D(net78),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[434] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[434] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit7  (.D(net79),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[460] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[460] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit8  (.D(net80),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[493] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[493] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame7_bit9  (.D(net81),
    .GATE(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[519] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[519] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit0  (.D(net50),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[351] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit1  (.D(net61),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[329] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit10  (.D(net51),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[538] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[538] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit11  (.D(net52),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[520] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[520] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit12  (.D(net53),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[580] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[580] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit13  (.D(net54),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[554] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[554] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit14  (.D(net55),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr.ConfigBits[15] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit15  (.D(net56),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[161] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit16  (.D(net57),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[4] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit17  (.D(net58),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[194] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit18  (.D(net59),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[193] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit19  (.D(net60),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[209] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit2  (.D(net72),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[369] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit20  (.D(net62),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[207] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit21  (.D(net63),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[230] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit22  (.D(net64),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[219] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit23  (.D(net65),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[215] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit24  (.D(net66),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[235] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit25  (.D(net67),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[244] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit26  (.D(net68),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[290] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit27  (.D(net69),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[286] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit28  (.D(net70),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[607] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[607] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit29  (.D(net71),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[600] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[600] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit3  (.D(net75),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[432] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[432] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit30  (.D(net73),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[598] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[598] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit31  (.D(net74),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[597] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[597] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit4  (.D(net76),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[427] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[427] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit5  (.D(net77),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[426] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[426] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit6  (.D(net78),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[443] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[443] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit7  (.D(net79),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[518] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[518] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit8  (.D(net80),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[523] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[523] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame8_bit9  (.D(net81),
    .GATE(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[539] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[539] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit0  (.D(net50),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[354] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit1  (.D(net61),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[350] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit10  (.D(net51),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[361] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit11  (.D(net52),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[419] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[419] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit12  (.D(net53),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[418] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[418] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit13  (.D(net54),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[414] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[414] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit14  (.D(net55),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[445] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[445] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit15  (.D(net56),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[525] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[525] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit16  (.D(net57),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[524] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[524] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit17  (.D(net58),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[541] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[541] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit18  (.D(net59),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[556] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[556] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit19  (.D(net60),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[583] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[583] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit2  (.D(net72),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[341] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit20  (.D(net62),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[579] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[579] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit21  (.D(net63),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr.ConfigBits[3] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit22  (.D(net64),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[197] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit23  (.D(net65),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[195] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit24  (.D(net66),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[218] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit25  (.D(net67),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[237] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit26  (.D(net68),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[245] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit27  (.D(net69),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[292] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit28  (.D(net70),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[281] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit29  (.D(net71),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[591] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[591] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit3  (.D(net75),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[328] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit30  (.D(net73),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[603] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[603] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit31  (.D(net74),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[599] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[599] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit4  (.D(net76),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[368] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit5  (.D(net77),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[384] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit6  (.D(net78),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[383] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit7  (.D(net79),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[382] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit8  (.D(net80),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[379] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem.Inst_Frame9_bit9  (.D(net81),
    .GATE(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\Inst_LUT4AB_ConfigMem.ConfigBits[378] ),
    .Q_N(\Inst_LUT4AB_ConfigMem.ConfigBits_N[378] ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._032_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._033_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._034_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._035_  (.A(net14),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb0 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._036_  (.A(net15),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._037_  (.A(net16),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb2 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._038_  (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._039_  (.A(net18),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb4 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._040_  (.A(net19),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._041_  (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._042_  (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEGb7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._043_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.F ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._044_  (.A(net540),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.G ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._045_  (.A(net515),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.H ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._046_  (.A(net1),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._047_  (.A(\Inst_LA_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._048_  (.A(\Inst_LB_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._049_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._050_  (.A(\Inst_LD_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._051_  (.A(\Inst_LE_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._052_  (.A(\Inst_LF_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._053_  (.A(\Inst_LG_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.Ci ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._054_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG0 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._055_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG1 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._056_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG2 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._057_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._058_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG4 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._059_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._060_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._061_  (.A(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEG7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._062_  (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb0 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._063_  (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._064_  (.A(net116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb2 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._065_  (.A(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._066_  (.A(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb4 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._067_  (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._068_  (.A(net120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._069_  (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N2BEGb7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._070_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._071_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._072_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG2 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._073_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG3 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._074_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG4 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._075_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG5 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._076_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._077_  (.A(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEG7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._078_  (.A(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._079_  (.A(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._080_  (.A(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._081_  (.A(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._082_  (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb4 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._083_  (.A(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._084_  (.A(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._085_  (.A(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2BEGb7 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._086_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._087_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG1 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._088_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._089_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._090_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG4 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._091_  (.A(net533),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._092_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG6 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._093_  (.A(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEG7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._094_  (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb0 ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._095_  (.A(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._096_  (.A(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._097_  (.A(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._098_  (.A(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb4 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._099_  (.A(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb5 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._100_  (.A(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb6 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._101_  (.A(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W2BEGb7 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._102_  (.A(net514),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.A ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._103_  (.A(net513),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.B ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._104_  (.A(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.C ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._105_  (.A(\Inst_LH_LUT4c_frame_config_dffesr.Co ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._106_  (.A(net510),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.D ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix._107_  (.A(net509),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E ));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix._108_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._109_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._110_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._111_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix._112_  (.A(\Inst_LUT4AB_switch_matrix.JE2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst0  (.A0(net5),
    .A1(net209),
    .A2(net514),
    .A3(net513),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[202] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst1  (.A0(net537),
    .A1(net510),
    .A2(net509),
    .A3(net541),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[202] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst2  (.A0(net540),
    .A1(net515),
    .A2(net542),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[202] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[202] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[203] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[204] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[205] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst0  (.A0(net4),
    .A1(net208),
    .A2(net514),
    .A3(net513),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[206] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst1  (.A0(net537),
    .A1(net510),
    .A2(net509),
    .A3(net541),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[206] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst2  (.A0(net511),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[206] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A3(net538),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[206] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[207] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[208] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[209] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net107),
    .A2(net129),
    .A3(net41),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[482] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst1  (.A0(net25),
    .A1(net159),
    .A2(net211),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[482] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst2  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A1(net512),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[482] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[482] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[483] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[484] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[485] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net108),
    .A2(net130),
    .A3(net8),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[486] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst1  (.A0(net22),
    .A1(net160),
    .A2(net212),
    .A3(net247),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[486] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst2  (.A0(net543),
    .A1(net512),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .A3(net535),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[486] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A3(net542),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[486] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[487] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[488] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[489] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net109),
    .A2(net131),
    .A3(net9),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[490] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst1  (.A0(net25),
    .A1(net161),
    .A2(net213),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[490] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .A1(net532),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .A3(net535),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[490] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[490] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[491] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[492] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[493] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net110),
    .A2(net122),
    .A3(net10),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[494] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst1  (.A0(net22),
    .A1(net162),
    .A2(net214),
    .A3(net226),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[494] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .A1(net513),
    .A2(net512),
    .A3(net535),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[494] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[494] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[495] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[496] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[497] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[498] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net163),
    .A3(net207),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[498] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst2  (.A0(net514),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[498] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst3  (.A0(net508),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[498] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[499] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[500] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[501] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[502] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net164),
    .A3(net208),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[502] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[502] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[502] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[503] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[504] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[505] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[506] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net165),
    .A3(net209),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[506] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[506] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[506] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[507] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[508] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[509] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net106),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[510] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net190),
    .A3(net238),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[510] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(net512),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[510] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst3  (.A0(net509),
    .A1(net508),
    .A2(net511),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[510] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[511] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[512] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[513] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JE2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst0  (.A0(net107),
    .A1(net129),
    .A2(net5),
    .A3(net7),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[450] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst1  (.A0(net25),
    .A1(net197),
    .A2(net211),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[450] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst2  (.A0(net513),
    .A1(net537),
    .A2(net510),
    .A3(net509),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[450] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst3  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[450] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[451] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[452] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[453] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst0  (.A0(net108),
    .A1(net130),
    .A2(net2),
    .A3(net8),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[454] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst1  (.A0(net22),
    .A1(net160),
    .A2(net212),
    .A3(net226),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[454] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net512),
    .A2(net510),
    .A3(net509),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[454] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[454] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[455] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[456] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[457] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst0  (.A0(net109),
    .A1(net131),
    .A2(net3),
    .A3(net9),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[458] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst1  (.A0(net25),
    .A1(net161),
    .A2(net213),
    .A3(net245),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[458] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(net510),
    .A3(net509),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[458] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[458] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[459] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[460] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[461] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst0  (.A0(net110),
    .A1(net122),
    .A2(net4),
    .A3(net10),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[462] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst1  (.A0(net22),
    .A1(net162),
    .A2(net214),
    .A3(net226),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[462] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst2  (.A0(net514),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(net512),
    .A3(net509),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[462] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[462] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[463] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[464] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[465] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[466] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst1  (.A0(net155),
    .A1(net163),
    .A2(net207),
    .A3(net209),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[466] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst2  (.A0(net514),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(net537),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[466] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst3  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[466] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[467] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[468] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[469] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[470] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst1  (.A0(net156),
    .A1(net164),
    .A2(net206),
    .A3(net208),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[470] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net532),
    .A2(net537),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[470] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[470] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[471] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[472] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[473] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[474] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst1  (.A0(net157),
    .A1(net165),
    .A2(net207),
    .A3(net209),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[474] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(net537),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[474] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[474] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[475] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[476] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[477] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net106),
    .A2(net2),
    .A3(net34),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[478] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst1  (.A0(net154),
    .A1(net158),
    .A2(net206),
    .A3(net208),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[478] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net532),
    .A2(net537),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[478] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst3  (.A0(net509),
    .A1(net541),
    .A2(net540),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[478] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[479] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[480] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[481] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JN2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst0  (.A0(net145),
    .A1(net5),
    .A2(net7),
    .A3(net25),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[514] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst1  (.A0(net159),
    .A1(net181),
    .A2(net211),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[514] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst2  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A1(net512),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[514] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[514] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[515] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[516] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[517] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst0  (.A0(net146),
    .A1(net2),
    .A2(net42),
    .A3(net22),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[518] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst1  (.A0(net182),
    .A1(net198),
    .A2(net212),
    .A3(net226),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[518] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net512),
    .A2(net510),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[518] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[518] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[519] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[520] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[521] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst0  (.A0(net147),
    .A1(net3),
    .A2(net9),
    .A3(net25),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[522] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst1  (.A0(net161),
    .A1(net183),
    .A2(net213),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[522] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[522] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[522] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[523] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[524] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[525] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst0  (.A0(net110),
    .A1(net4),
    .A2(net10),
    .A3(net22),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[526] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst1  (.A0(net162),
    .A1(net174),
    .A2(net214),
    .A3(net246),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[526] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(net512),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[526] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[526] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[527] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[528] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[529] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[530] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst1  (.A0(net155),
    .A1(net163),
    .A2(net207),
    .A3(net209),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[530] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[530] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst3  (.A0(net508),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[530] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[531] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[532] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[533] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[534] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst1  (.A0(net156),
    .A1(net164),
    .A2(net206),
    .A3(net208),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[534] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[534] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[534] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[535] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[536] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[537] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[538] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst1  (.A0(net157),
    .A1(net165),
    .A2(net207),
    .A3(net209),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[538] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[538] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst3  (.A0(net509),
    .A1(net541),
    .A2(net515),
    .A3(net542),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[538] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[539] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[540] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[541] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net106),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[542] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst1  (.A0(net154),
    .A1(net158),
    .A2(net206),
    .A3(net208),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[542] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .A1(net532),
    .A2(net512),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[542] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst3  (.A0(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .A1(net508),
    .A2(net511),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[542] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[543] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[544] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[545] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JS2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net107),
    .A2(net7),
    .A3(net25),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[546] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst1  (.A0(net159),
    .A1(net181),
    .A2(net211),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[546] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst2  (.A0(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A1(net537),
    .A2(net510),
    .A3(net509),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[546] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst3  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[546] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[547] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[548] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[549] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net108),
    .A2(net8),
    .A3(net22),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[550] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst1  (.A0(net160),
    .A1(net182),
    .A2(net212),
    .A3(net226),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[550] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net512),
    .A2(net510),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[550] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[550] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[551] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[552] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[553] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net109),
    .A2(net43),
    .A3(net25),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[554] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst1  (.A0(net183),
    .A1(net199),
    .A2(net213),
    .A3(net229),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[554] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(net510),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[554] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst3  (.A0(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A1(net511),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[554] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[555] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[556] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[557] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net110),
    .A2(net10),
    .A3(net22),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[558] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst1  (.A0(net162),
    .A1(net174),
    .A2(net214),
    .A3(net246),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[558] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst2  (.A0(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(net512),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[558] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst3  (.A0(net508),
    .A1(net511),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[558] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[559] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[560] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[561] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[562] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net163),
    .A3(net207),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[562] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst2  (.A0(net514),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[562] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst3  (.A0(net508),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AD ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[562] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[563] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[564] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[565] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[566] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net164),
    .A3(net208),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[566] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net532),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[566] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[566] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[567] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[568] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[569] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[570] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net165),
    .A3(net209),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[570] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst2  (.A0(net514),
    .A1(net513),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[570] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst3  (.A0(net509),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .A2(net515),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[570] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[571] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[572] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[573] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net138),
    .A2(net2),
    .A3(net6),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[574] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net158),
    .A3(net206),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[574] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst2  (.A0(net543),
    .A1(net532),
    .A2(net512),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[574] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst3  (.A0(net535),
    .A1(net508),
    .A2(net511),
    .A3(\Inst_LUT4AB_switch_matrix.M_AB ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[574] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[575] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[576] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[577] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.JW2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst0  (.A0(net5),
    .A1(net209),
    .A2(net514),
    .A3(net532),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[258] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst1  (.A0(net537),
    .A1(net510),
    .A2(net509),
    .A3(net508),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[258] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst2  (.A0(net540),
    .A1(net515),
    .A2(net542),
    .A3(\Inst_LUT4AB_switch_matrix.M_AH ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[258] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[258] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[259] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[260] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[261] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst0  (.A0(net4),
    .A1(net208),
    .A2(net514),
    .A3(net532),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[262] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst1  (.A0(net512),
    .A1(net510),
    .A2(net509),
    .A3(net508),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[262] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst2  (.A0(net511),
    .A1(net515),
    .A2(\Inst_LUT4AB_switch_matrix.M_AD ),
    .A3(\Inst_LUT4AB_switch_matrix.M_EF ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[262] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A3(net539),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[262] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[263] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[264] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[265] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W6BEG1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[266] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[266] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst0._0_  (.A(net524),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst0._0__524  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net524));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[275] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[275] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst0._0_  (.A(net516),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst0._0__516  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net516));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[276] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[276] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst0._0_  (.A(net525),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst0._0__525  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net525));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[285] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[285] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst0._0_  (.A(net517),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst0._0__517  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net517));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[286] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[286] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst0._0_  (.A(net526),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst0._0__526  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net526));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[295] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[295] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst0._0_  (.A(net518),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst0._0__518  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net518));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[296] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[296] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst0._0_  (.A(net527),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst0._0__527  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net527));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[305] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[305] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst0._0_  (.A(net519),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst0._0__519  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net519));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[306] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[306] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst0._0_  (.A(net528),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst0._0__528  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net528));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[315] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[315] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst0._0_  (.A(net520),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst0._0__520  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net520));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[316] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[316] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst0._0_  (.A(net529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst0._0__529  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net529));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[325] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[325] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst0._0_  (.A(net521),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst0._0__521  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net521));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[326] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[326] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst0._0_  (.A(net530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst0._0__530  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net530));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[335] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[335] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst0._0_  (.A(net522),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst0._0__522  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net522));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[336] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[336] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.EN ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst0._0_  (.A(net531),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst0._0__531  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net531));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[345] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[345] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr.SR ));
 sky130_fd_sc_hd__buf_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst0._0_  (.A(net523),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst0._0__523  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net523));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG0  (.A0(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[182] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[183] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG1  (.A0(net535),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[184] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[185] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG2  (.A0(net541),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[186] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[187] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG3  (.A0(net540),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[188] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[189] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(net112),
    .A1(net12),
    .A2(net199),
    .A3(net216),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[418] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[419] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(net138),
    .A1(net8),
    .A2(net160),
    .A3(net212),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[420] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[421] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(net110),
    .A1(net34),
    .A2(net162),
    .A3(net214),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[422] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[423] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(net106),
    .A1(net6),
    .A2(net158),
    .A3(net247),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[424] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[425] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(net147),
    .A1(net12),
    .A2(net164),
    .A3(net216),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[426] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[427] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(net108),
    .A1(net8),
    .A2(net160),
    .A3(net246),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[428] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[429] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(net110),
    .A1(net10),
    .A2(net198),
    .A3(net214),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[430] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[431] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(net106),
    .A1(net41),
    .A2(net158),
    .A3(net210),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[432] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[433] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(net113),
    .A1(net42),
    .A2(net165),
    .A3(net217),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[434] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[435] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(net109),
    .A1(net9),
    .A2(net161),
    .A3(net245),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[436] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[437] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(net111),
    .A1(net11),
    .A2(net197),
    .A3(net215),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[438] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[439] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(net146),
    .A1(net7),
    .A2(net159),
    .A3(net211),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[440] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[441] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(net113),
    .A1(net13),
    .A2(net165),
    .A3(net238),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[442] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[443] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(net109),
    .A1(net9),
    .A2(net190),
    .A3(net213),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[444] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[445] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(net145),
    .A1(net11),
    .A2(net163),
    .A3(net215),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[446] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[447] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(net107),
    .A1(net43),
    .A2(net159),
    .A3(net211),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[448] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[449] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(net120),
    .A1(net172),
    .A2(net224),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[354] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[355] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net16),
    .A1(net168),
    .A2(net220),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[356] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[357] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net222),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[358] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[359] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net166),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[360] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[361] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[386] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[387] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[388] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[389] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[390] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[391] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[392] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[393] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net20),
    .A1(net172),
    .A2(net224),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[362] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[363] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net220),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[364] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[365] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net170),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[366] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[367] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(net114),
    .A1(net166),
    .A2(net218),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[368] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[369] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[394] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[395] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[396] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[397] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[398] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[399] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[400] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[401] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net224),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[370] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[371] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net168),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[372] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[373] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(net118),
    .A1(net170),
    .A2(net222),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[374] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[375] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net14),
    .A1(net166),
    .A2(net218),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[376] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[377] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[402] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[403] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[404] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[405] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[406] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[407] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[408] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[409] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net172),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[378] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[379] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(net116),
    .A1(net168),
    .A2(net220),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[380] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[381] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net18),
    .A1(net170),
    .A2(net222),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[382] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[383] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net218),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[384] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[385] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[410] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[411] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[412] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[413] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[414] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[415] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[416] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[417] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(net147),
    .A1(net183),
    .A2(net238),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[578] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[579] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net42),
    .A1(net182),
    .A2(net217),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[580] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[581] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(net129),
    .A1(net25),
    .A2(net229),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[582] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[583] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(net122),
    .A1(net22),
    .A2(net174),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[584] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[585] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net9),
    .A1(net199),
    .A2(net246),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[586] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[587] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(net130),
    .A1(net8),
    .A2(net217),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[588] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[589] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(net145),
    .A1(net41),
    .A2(net181),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[590] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[591] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(net122),
    .A1(net190),
    .A2(net226),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[592] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[593] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(net131),
    .A1(net9),
    .A2(net213),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[594] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[595] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(net146),
    .A1(net8),
    .A2(net182),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[596] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[597] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(net129),
    .A1(net197),
    .A2(net214),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[598] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[599] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net43),
    .A1(net174),
    .A2(net245),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[600] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[601] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(net131),
    .A1(net34),
    .A2(net183),
    .A3(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[602] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[603] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(net130),
    .A1(net198),
    .A2(net212),
    .A3(\Inst_LUT4AB_switch_matrix.JE2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[604] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[605] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net25),
    .A1(net181),
    .A2(net247),
    .A3(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[606] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[607] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(net138),
    .A1(net22),
    .A2(net210),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[608] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[609] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[267] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[268] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[269] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[270] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[271] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[272] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[273] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[274] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LA_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[277] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[278] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[279] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[280] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[281] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[282] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[283] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[284] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LB_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[287] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[288] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[289] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[290] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[291] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[292] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[293] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[294] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LC_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[297] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[298] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[299] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[300] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[301] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[302] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[303] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[304] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LD_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[307] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[308] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[309] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[310] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[311] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[312] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[313] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[314] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LE_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[317] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[318] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[319] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[320] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[321] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[322] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[323] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[324] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LF_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[327] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[328] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[329] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[330] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[331] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[332] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[333] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[334] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LG_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[337] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[338] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.I[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I1  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[339] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[340] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.I[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I2  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[341] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[342] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.I[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I3  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[343] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[344] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LH_LUT4c_frame_config_dffesr.I[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG0  (.A0(net512),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[154] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[155] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG1  (.A0(net510),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[156] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[157] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG1 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG2  (.A0(net509),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[158] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[159] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG3  (.A0(net541),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[160] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[161] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N1BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG0  (.A0(net108),
    .A1(net129),
    .A2(net25),
    .A3(net509),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[162] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[163] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG1  (.A0(net109),
    .A1(net130),
    .A2(net22),
    .A3(net508),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[164] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[165] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG2  (.A0(net106),
    .A1(net131),
    .A2(net229),
    .A3(net540),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[166] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[167] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG3  (.A0(net107),
    .A1(net122),
    .A2(net226),
    .A3(net515),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[168] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[169] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.N4BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S0  (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG4 ),
    .A1(\Inst_LUT4AB_switch_matrix.JE2BEG4 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG4 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG4 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[346] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[347] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S0 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1  (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG5 ),
    .A1(\Inst_LUT4AB_switch_matrix.JE2BEG5 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG5 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[348] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[349] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG0  (.A0(net535),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.JE2BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[210] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[211] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG1  (.A0(net508),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.JE2BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[212] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[213] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG2  (.A0(net511),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.JE2BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[214] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[215] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG3  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.JE2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[216] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[217] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S1BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S2  (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG6 ),
    .A1(\Inst_LUT4AB_switch_matrix.JE2BEG6 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG6 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG6 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[350] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[351] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S3  (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG7 ),
    .A1(\Inst_LUT4AB_switch_matrix.JE2BEG7 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG7 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG7 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[352] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[353] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG0  (.A0(net25),
    .A1(net160),
    .A2(net181),
    .A3(net543),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[218] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[219] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG1  (.A0(net22),
    .A1(net161),
    .A2(net182),
    .A3(net532),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[220] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[221] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG2  (.A0(net158),
    .A1(net183),
    .A2(net229),
    .A3(net512),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[222] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[223] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG3  (.A0(net159),
    .A1(net174),
    .A2(net226),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[224] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[225] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.S4BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG0  (.A0(net508),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[238] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[239] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG1  (.A0(net511),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[240] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[241] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG2  (.A0(net515),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[242] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[243] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG2 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG3  (.A0(net543),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[244] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[245] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.W1BEG3 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[192] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[192] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net156),
    .A3(net541),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[190] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst1  (.A0(net540),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[190] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[191] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[195] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[195] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net5),
    .A2(net157),
    .A3(net543),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[193] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst1  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[193] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[194] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[198] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[198] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net154),
    .A3(net513),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[196] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst1  (.A0(net512),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[196] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[197] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[201] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[201] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net155),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[199] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst1  (.A0(net535),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[199] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[200] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[615] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[615] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.J_EN_BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux41_buf_inst0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[613] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[614] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux41_buf_inst1  (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG2 ),
    .A1(\Inst_LUT4AB_switch_matrix.JE2BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[613] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[614] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[612] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[612] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.J_SR_BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux41_buf_inst0  (.A0(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0 ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[610] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[611] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux41_buf_inst1  (.A0(\Inst_LUT4AB_switch_matrix.JN2BEG1 ),
    .A1(\Inst_LUT4AB_switch_matrix.JE2BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.JS2BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.JW2BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[610] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[611] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[172] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[172] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net208),
    .A3(net541),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[170] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst1  (.A0(net540),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[170] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[171] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[175] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[175] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net5),
    .A2(net209),
    .A3(net514),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[173] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst1  (.A0(net515),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[173] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[174] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[178] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[178] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net206),
    .A3(net513),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[176] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst1  (.A0(net537),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[176] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[177] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[181] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[181] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.NN4BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net207),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[179] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst1  (.A0(net509),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A2(net538),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[179] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[180] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[228] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[228] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net208),
    .A3(net541),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[226] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst1  (.A0(net540),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[226] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[227] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[231] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[231] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net5),
    .A2(net209),
    .A3(net543),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[229] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst1  (.A0(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[229] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[230] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[234] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[234] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net206),
    .A3(net532),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[232] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst1  (.A0(net512),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[232] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[233] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[237] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[237] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.SS4BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net207),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[235] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst1  (.A0(net535),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A2(net539),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[235] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[236] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[248] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[248] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst0  (.A0(net104),
    .A1(net156),
    .A2(net208),
    .A3(net508),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[246] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst1  (.A0(net540),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_GH_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[246] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[247] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[251] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[251] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst0  (.A0(net105),
    .A1(net157),
    .A2(net209),
    .A3(net514),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[249] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst1  (.A0(net515),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_EF_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[249] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[250] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[254] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[254] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst0  (.A0(net102),
    .A1(net154),
    .A2(net206),
    .A3(net532),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[252] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst1  (.A0(net512),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 ),
    .A2(\Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 ),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_CD_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[252] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[253] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._2_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._3_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[257] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[257] ),
    .A2(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._0_ ),
    .B1(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.WW4BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst0  (.A0(net103),
    .A1(net155),
    .A2(net207),
    .A3(net510),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[255] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[256] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst1  (.A0(net535),
    .A1(\Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 ),
    .A2(net539),
    .A3(\Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 ),
    .S0(\Inst_LUT4AB_ConfigMem.ConfigBits[255] ),
    .S1(\Inst_LUT4AB_ConfigMem.ConfigBits[256] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN[1] ),
    .B(\Inst_LUT4AB_switch_matrix.S0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._4_  (.A1(net534),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.M_AB ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.B ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN[1] ),
    .B(\Inst_LUT4AB_switch_matrix.S1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._4_  (.A1(\Inst_LUT4AB_switch_matrix.S1 ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.AD ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.break_comb_loop_inst0._0_  (.A(net542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.CD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN[1] ),
    .B(\Inst_LUT4AB_switch_matrix.S3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._4_  (.A1(\Inst_LUT4AB_switch_matrix.S3 ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.AH ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.break_comb_loop_inst0._0_  (.A(\Inst_MUX8LUT_frame_config_mux.AD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.EH ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN[1] ),
    .B(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._4_  (.A1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.CD ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.C ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.D ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN[1] ),
    .B(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._4_  (.A1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.M_EF ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.E ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.F ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN[1] ),
    .B(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._4_  (.A1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.EH ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.M_EF ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.GH ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.EH_GH ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.break_comb_loop_inst0._0_  (.A(\Inst_MUX8LUT_frame_config_mux.GH ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.EH ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN[1] ),
    .B(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._4_  (.A1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.GH ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.G ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.H ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.M_AD ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.break_comb_loop_inst0._0_  (.A(\Inst_MUX8LUT_frame_config_mux.CD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.AD ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_LUT4AB_switch_matrix.M_AH ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.break_comb_loop_inst0._0_  (.A(\Inst_MUX8LUT_frame_config_mux.EH_GH ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.AH ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.S1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.S0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.S2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.S0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[153] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.break_comb_loop_inst0._0_  (.A(\Inst_LUT4AB_switch_matrix.S3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.break_comb_loop_inst1._0_  (.A(\Inst_LUT4AB_switch_matrix.S1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._2_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._3_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN[1] ),
    .B(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._4_  (.A1(\Inst_LUT4AB_ConfigMem.ConfigBits[152] ),
    .A2(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._0_ ),
    .B1(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._1_ ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(\Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.break_comb_loop_inst0._0_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.break_comb_loop_inst1._0_  (.A(\Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN[1] ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_0._0_  (.A(\N4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_1._0_  (.A(\N4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_10._0_  (.A(\N4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_11._0_  (.A(\N4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_2._0_  (.A(\N4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_3._0_  (.A(\N4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_4._0_  (.A(\N4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_5._0_  (.A(\N4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_6._0_  (.A(\N4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_7._0_  (.A(\N4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_8._0_  (.A(\N4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_9._0_  (.A(\N4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_4 \N4END_inbuf_0._0_  (.A(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_1._0_  (.A(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_4 \N4END_inbuf_10._0_  (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_11._0_  (.A(net128),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_2._0_  (.A(net134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_3._0_  (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_4._0_  (.A(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_5._0_  (.A(net137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_6._0_  (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_7._0_  (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_8._0_  (.A(net125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_9._0_  (.A(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\N4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_0._0_  (.A(\NN4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_1._0_  (.A(\NN4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_10._0_  (.A(\NN4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_11._0_  (.A(\NN4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_2._0_  (.A(\NN4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_3._0_  (.A(\NN4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_4._0_  (.A(\NN4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_5._0_  (.A(\NN4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_6._0_  (.A(\NN4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_7._0_  (.A(\NN4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_8._0_  (.A(\NN4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_9._0_  (.A(\NN4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_0._0_  (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_1._0_  (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_10._0_  (.A(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_11._0_  (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_2._0_  (.A(net150),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_3._0_  (.A(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_4._0_  (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_5._0_  (.A(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_6._0_  (.A(net139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_7._0_  (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_8._0_  (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_9._0_  (.A(net142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\NN4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_0._0_  (.A(\S4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_1._0_  (.A(\S4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_10._0_  (.A(\S4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_11._0_  (.A(\S4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_2._0_  (.A(\S4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_3._0_  (.A(\S4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_4 \S4BEG_outbuf_4._0_  (.A(\S4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_5._0_  (.A(\S4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__buf_2 \S4BEG_outbuf_6._0_  (.A(\S4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_7._0_  (.A(\S4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_8._0_  (.A(\S4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_2 \S4BEG_outbuf_9._0_  (.A(\S4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_0._0_  (.A(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_1._0_  (.A(net185),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_10._0_  (.A(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_11._0_  (.A(net180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_2._0_  (.A(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_3._0_  (.A(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_4._0_  (.A(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_5._0_  (.A(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_6._0_  (.A(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_7._0_  (.A(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_8._0_  (.A(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_1 \S4END_inbuf_9._0_  (.A(net178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\S4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__buf_2 \SS4BEG_outbuf_0._0_  (.A(\SS4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_1._0_  (.A(\SS4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__buf_2 \SS4BEG_outbuf_10._0_  (.A(\SS4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_11._0_  (.A(\SS4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__buf_2 \SS4BEG_outbuf_2._0_  (.A(\SS4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_3._0_  (.A(\SS4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__buf_2 \SS4BEG_outbuf_4._0_  (.A(\SS4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_5._0_  (.A(\SS4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__buf_2 \SS4BEG_outbuf_6._0_  (.A(\SS4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_7._0_  (.A(\SS4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_8._0_  (.A(\SS4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_2 \SS4BEG_outbuf_9._0_  (.A(\SS4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_0._0_  (.A(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_1._0_  (.A(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_10._0_  (.A(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_11._0_  (.A(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_2._0_  (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_3._0_  (.A(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_4._0_  (.A(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_5._0_  (.A(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_6._0_  (.A(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_7._0_  (.A(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_8._0_  (.A(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_1 \SS4END_inbuf_9._0_  (.A(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\SS4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_0._0_  (.A(\W6BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_1._0_  (.A(\W6BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_2._0_  (.A(\W6BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_3._0_  (.A(\W6BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_4._0_  (.A(\W6BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_5._0_  (.A(\W6BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_6._0_  (.A(\W6BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_7._0_  (.A(\W6BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_8._0_  (.A(\W6BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_2 \W6BEG_outbuf_9._0_  (.A(\W6BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_0._0_  (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_1._0_  (.A(net231),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_2._0_  (.A(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_3._0_  (.A(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_4._0_  (.A(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_5._0_  (.A(net235),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_6._0_  (.A(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_7._0_  (.A(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_8._0_  (.A(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_1 \W6END_inbuf_9._0_  (.A(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\W6BEG_outbuf_9.A ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_0._0_  (.A(\WW4BEG_outbuf_0.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_1._0_  (.A(\WW4BEG_outbuf_1.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_10._0_  (.A(\WW4BEG_outbuf_10.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_11._0_  (.A(\WW4BEG_outbuf_11.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_2._0_  (.A(\WW4BEG_outbuf_2.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_3._0_  (.A(\WW4BEG_outbuf_3.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_4._0_  (.A(\WW4BEG_outbuf_4.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_5._0_  (.A(\WW4BEG_outbuf_5.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_6._0_  (.A(\WW4BEG_outbuf_6.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_7._0_  (.A(\WW4BEG_outbuf_7.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_8._0_  (.A(\WW4BEG_outbuf_8.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_2 \WW4BEG_outbuf_9._0_  (.A(\WW4BEG_outbuf_9.A ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_0._0_  (.A(net248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_0.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_1._0_  (.A(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_1.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_10._0_  (.A(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_10.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_11._0_  (.A(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_11.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_2._0_  (.A(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_2.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_3._0_  (.A(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_3.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_4._0_  (.A(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_4.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_5._0_  (.A(net253),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_5.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_6._0_  (.A(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_6.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_7._0_  (.A(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_7.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_8._0_  (.A(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_8.A ));
 sky130_fd_sc_hd__clkbuf_1 \WW4END_inbuf_9._0_  (.A(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\WW4BEG_outbuf_9.A ));
 sky130_fd_sc_hd__clkbuf_1 _000_ (.A(\data_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 _001_ (.A(\data_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 _002_ (.A(\data_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 _003_ (.A(\data_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 _004_ (.A(\data_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 _005_ (.A(\data_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 _006_ (.A(\data_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 _007_ (.A(\data_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 _008_ (.A(\data_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 _009_ (.A(\data_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_1 _010_ (.A(\data_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 _011_ (.A(\data_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 _012_ (.A(\data_outbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 _013_ (.A(\data_outbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 _014_ (.A(\data_outbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 _015_ (.A(\data_outbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 _016_ (.A(\data_outbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 _017_ (.A(\data_outbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 _018_ (.A(\data_outbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 _019_ (.A(\data_outbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 _020_ (.A(\data_outbuf_20.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 _021_ (.A(\data_outbuf_21.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 _022_ (.A(\data_outbuf_22.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 _023_ (.A(\data_outbuf_23.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 _024_ (.A(\data_outbuf_24.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 _025_ (.A(\data_outbuf_25.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 _026_ (.A(\data_outbuf_26.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 _027_ (.A(\data_outbuf_27.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 _028_ (.A(\data_outbuf_28.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 _029_ (.A(\data_outbuf_29.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 _030_ (.A(\data_outbuf_30.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 _031_ (.A(\data_outbuf_31.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 _032_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 _033_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 _034_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 _035_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 _036_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 _037_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 _038_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _039_ (.A(\Inst_LUT4AB_switch_matrix.E2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 _040_ (.A(\E6BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 _041_ (.A(\E6BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 _042_ (.A(\E6BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 _043_ (.A(\E6BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 _044_ (.A(\E6BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 _045_ (.A(\E6BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 _046_ (.A(\E6BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 _047_ (.A(\E6BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 _048_ (.A(\E6BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 _049_ (.A(\E6BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_1 _050_ (.A(\Inst_LUT4AB_switch_matrix.E6BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 _051_ (.A(\Inst_LUT4AB_switch_matrix.E6BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 _052_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__buf_1 _053_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 _054_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 _055_ (.A(\Inst_LUT4AB_switch_matrix.E1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__buf_1 _056_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 _057_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 _058_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 _059_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 _060_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 _061_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__buf_1 _062_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 _063_ (.A(\Inst_LUT4AB_switch_matrix.E2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 _064_ (.A(\strobe_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(\strobe_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 _066_ (.A(\strobe_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(\strobe_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 _068_ (.A(\strobe_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 _069_ (.A(\strobe_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 _070_ (.A(\strobe_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(\strobe_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(\strobe_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(\strobe_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(\strobe_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(\strobe_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(\strobe_outbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(\strobe_outbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(\strobe_outbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(\strobe_outbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 _080_ (.A(\strobe_outbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 _081_ (.A(\strobe_outbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 _082_ (.A(\strobe_outbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 _083_ (.A(\strobe_outbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(\EE4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(\EE4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 _086_ (.A(\EE4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 _087_ (.A(\EE4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(\EE4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(\EE4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(\EE4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(\EE4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(\EE4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(\EE4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(\EE4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(\EE4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(\Inst_LUT4AB_switch_matrix.EE4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(\Inst_LUT4AB_switch_matrix.N1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_1 _104_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_1 _106_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 _107_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 _108_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 _109_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 _110_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(\Inst_LUT4AB_switch_matrix.N2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 _112_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 _113_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 _114_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 _115_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 _118_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(\Inst_LUT4AB_switch_matrix.N2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 _120_ (.A(\N4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 _121_ (.A(\N4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(\N4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(\N4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 _124_ (.A(\N4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 _125_ (.A(\N4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 _126_ (.A(\N4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(\N4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 _128_ (.A(\N4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 _129_ (.A(\N4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 _130_ (.A(\N4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(\N4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 _134_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(\Inst_LUT4AB_switch_matrix.N4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 _136_ (.A(\NN4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 _137_ (.A(\NN4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 _138_ (.A(\NN4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 _139_ (.A(\NN4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 _140_ (.A(\NN4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 _141_ (.A(\NN4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 _142_ (.A(\NN4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 _143_ (.A(\NN4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 _144_ (.A(\NN4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 _145_ (.A(\NN4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 _146_ (.A(\NN4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 _147_ (.A(\NN4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 _148_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 _149_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 _150_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 _151_ (.A(\Inst_LUT4AB_switch_matrix.NN4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 _152_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_1 _153_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 _154_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 _155_ (.A(\Inst_LUT4AB_switch_matrix.S1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net410));
 sky130_fd_sc_hd__buf_1 _156_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 _157_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 _158_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 _159_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 _160_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 _161_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 _162_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net417));
 sky130_fd_sc_hd__buf_1 _163_ (.A(\Inst_LUT4AB_switch_matrix.S2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 _164_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 _165_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_1 _166_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 _167_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 _168_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 _169_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 _170_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 _171_ (.A(\Inst_LUT4AB_switch_matrix.S2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 _172_ (.A(\S4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 _173_ (.A(\S4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 _174_ (.A(\S4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 _175_ (.A(\S4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 _176_ (.A(\S4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 _177_ (.A(\S4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 _178_ (.A(\S4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 _179_ (.A(\S4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 _180_ (.A(\S4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 _181_ (.A(\S4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_1 _182_ (.A(\S4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 _183_ (.A(\S4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 _184_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_1 _185_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 _186_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_1 _187_ (.A(\Inst_LUT4AB_switch_matrix.S4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_1 _188_ (.A(\SS4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 _189_ (.A(\SS4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 _190_ (.A(\SS4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 _191_ (.A(\SS4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 _192_ (.A(\SS4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 _193_ (.A(\SS4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(\SS4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 _195_ (.A(\SS4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 _196_ (.A(\SS4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 _197_ (.A(\SS4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 _198_ (.A(\SS4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 _199_ (.A(\SS4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 _200_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_1 _201_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_1 _202_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_1 _203_ (.A(\Inst_LUT4AB_switch_matrix.SS4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_1 _205_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_1 _206_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_1 _207_ (.A(\Inst_LUT4AB_switch_matrix.W1BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_1 _208_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 _209_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 _210_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 _211_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 _212_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 _213_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 _214_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 _215_ (.A(\Inst_LUT4AB_switch_matrix.W2BEG7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 _216_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_1 _217_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 _218_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 _219_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_1 _220_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb4 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_1 _221_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_1 _222_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb6 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_1 _223_ (.A(\Inst_LUT4AB_switch_matrix.W2BEGb7 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_1 _224_ (.A(\W6BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 _225_ (.A(\W6BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_1 _226_ (.A(\W6BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 _227_ (.A(\W6BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 _228_ (.A(\W6BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 _229_ (.A(\W6BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 _230_ (.A(\W6BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 _231_ (.A(\W6BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 _232_ (.A(\W6BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_1 _233_ (.A(\W6BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_1 _234_ (.A(\Inst_LUT4AB_switch_matrix.W6BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_1 _235_ (.A(\Inst_LUT4AB_switch_matrix.W6BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_1 _236_ (.A(\WW4BEG_outbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 _237_ (.A(\WW4BEG_outbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 _238_ (.A(\WW4BEG_outbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 _239_ (.A(\WW4BEG_outbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 _240_ (.A(\WW4BEG_outbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_1 _241_ (.A(\WW4BEG_outbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 _242_ (.A(\WW4BEG_outbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 _243_ (.A(\WW4BEG_outbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 _244_ (.A(\WW4BEG_outbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_1 _245_ (.A(\WW4BEG_outbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_1 _246_ (.A(\WW4BEG_outbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 _247_ (.A(\WW4BEG_outbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_1 _248_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net495));
 sky130_fd_sc_hd__clkbuf_1 _249_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG1 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_1 _250_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 _251_ (.A(\Inst_LUT4AB_switch_matrix.WW4BEG3 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_0._0_  (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_1._0_  (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_10._0_  (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11._0_  (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_12._0_  (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_13._0_  (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14._0_  (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_15._0_  (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_16._0_  (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_17._0_  (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18._0_  (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19._0_  (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_2._0_  (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20._0_  (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_20.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_21._0_  (.A(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_21.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22._0_  (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_22.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23._0_  (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_23.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24._0_  (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_24.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25._0_  (.A(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_25.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26._0_  (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_26.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_27._0_  (.A(net69),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_27.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_28._0_  (.A(net70),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_28.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_29._0_  (.A(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_29.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_3._0_  (.A(net75),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_30._0_  (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_30.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31._0_  (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_31.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_4._0_  (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_5._0_  (.A(net77),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_6._0_  (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_7._0_  (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_8._0_  (.A(net80),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_9._0_  (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_inbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0._0_  (.A(\data_inbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1._0_  (.A(\data_inbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10._0_  (.A(\data_inbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11._0_  (.A(\data_inbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12._0_  (.A(\data_inbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13._0_  (.A(\data_inbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14._0_  (.A(\data_inbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15._0_  (.A(\data_inbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16._0_  (.A(\data_inbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17._0_  (.A(\data_inbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18._0_  (.A(\data_inbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19._0_  (.A(\data_inbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2._0_  (.A(\data_inbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20._0_  (.A(\data_inbuf_20.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_20.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21._0_  (.A(\data_inbuf_21.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_21.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22._0_  (.A(\data_inbuf_22.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_22.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23._0_  (.A(\data_inbuf_23.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_23.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24._0_  (.A(\data_inbuf_24.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_24.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25._0_  (.A(\data_inbuf_25.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_25.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26._0_  (.A(\data_inbuf_26.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_26.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27._0_  (.A(\data_inbuf_27.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_27.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28._0_  (.A(\data_inbuf_28.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_28.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29._0_  (.A(\data_inbuf_29.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_29.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3._0_  (.A(\data_inbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30._0_  (.A(\data_inbuf_30.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_30.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31._0_  (.A(\data_inbuf_31.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_31.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4._0_  (.A(\data_inbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5._0_  (.A(\data_inbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6._0_  (.A(\data_inbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7._0_  (.A(\data_inbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8._0_  (.A(\data_inbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9._0_  (.A(\data_inbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\data_outbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(Ci),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(E2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_16 input100 (.A(FrameStrobe[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_16 input101 (.A(FrameStrobe[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__buf_4 input102 (.A(N1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__buf_4 input103 (.A(N1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__buf_4 input104 (.A(N1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__buf_4 input105 (.A(N1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(N2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__buf_2 input107 (.A(N2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(N2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__buf_2 input109 (.A(N2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(E2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(N2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(N2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(N2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(N2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(N2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(N2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(N2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_2 input117 (.A(N2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(N2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(N2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(E2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(N2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(N2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(N4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(N4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(N4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(N4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(N4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(N4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(N4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__buf_2 input129 (.A(N4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input13 (.A(E2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input130 (.A(N4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 input131 (.A(N4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(N4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(N4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(N4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(N4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(N4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(N4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(NN4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(NN4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(E2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(NN4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(NN4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(NN4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(NN4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(NN4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 input145 (.A(NN4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(NN4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(NN4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(NN4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(NN4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__buf_2 input15 (.A(E2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(NN4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(NN4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(NN4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(NN4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(S1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(S1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__buf_4 input156 (.A(S1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(S1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__buf_4 input158 (.A(S2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(S2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input16 (.A(E2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input160 (.A(S2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__buf_2 input161 (.A(S2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(S2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(S2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(S2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(S2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(S2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 input167 (.A(S2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__buf_2 input168 (.A(S2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 input169 (.A(S2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(E2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input170 (.A(S2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(S2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(S2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(S2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__buf_2 input174 (.A(S4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(S4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(S4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(S4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(S4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(S4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__buf_2 input18 (.A(E2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(S4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_4 input181 (.A(S4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(S4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__buf_2 input183 (.A(S4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(S4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(S4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(S4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(S4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(S4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(S4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(E2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(SS4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(SS4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(SS4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(SS4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(SS4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(SS4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(SS4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(SS4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(SS4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input199 (.A(SS4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__buf_4 input2 (.A(E1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(E2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(SS4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(SS4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(SS4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(SS4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(SS4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(SS4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__buf_4 input206 (.A(W1END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__buf_4 input207 (.A(W1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 input208 (.A(W1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 input209 (.A(W1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__buf_2 input21 (.A(E2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__dlymetal6s2s_1 input210 (.A(W2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 input211 (.A(W2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__buf_2 input212 (.A(W2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 input213 (.A(W2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(W2END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 input215 (.A(W2END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 input216 (.A(W2END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(W2END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__buf_2 input218 (.A(W2MID[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 input219 (.A(W2MID[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__buf_4 input22 (.A(E6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input220 (.A(W2MID[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__buf_2 input221 (.A(W2MID[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 input222 (.A(W2MID[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 input223 (.A(W2MID[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 input224 (.A(W2MID[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__buf_2 input225 (.A(W2MID[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 input226 (.A(W6END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(W6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(W6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__buf_4 input229 (.A(W6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(E6END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(W6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(W6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(W6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(W6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(W6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(W6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(W6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(W6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__buf_2 input238 (.A(WW4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(WW4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(E6END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(WW4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(WW4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(WW4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(WW4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(WW4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 input245 (.A(WW4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__buf_2 input246 (.A(WW4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 input247 (.A(WW4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(WW4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(WW4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__buf_4 input25 (.A(E6END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(WW4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(WW4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(WW4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(WW4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(E6END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(E6END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(E6END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(E6END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(E1END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(E6END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(E6END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(E6END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(E6END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(EE4END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(EE4END[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(EE4END[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(EE4END[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(EE4END[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(EE4END[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(E1END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(EE4END[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(EE4END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(EE4END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(EE4END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(EE4END[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(EE4END[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(EE4END[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(EE4END[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(EE4END[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(EE4END[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(E1END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input50 (.A(FrameData[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__buf_8 input51 (.A(FrameData[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(FrameData[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__buf_8 input53 (.A(FrameData[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_8 input54 (.A(FrameData[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__buf_8 input55 (.A(FrameData[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__buf_8 input56 (.A(FrameData[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net56));
 sky130_fd_sc_hd__buf_8 input57 (.A(FrameData[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net57));
 sky130_fd_sc_hd__buf_8 input58 (.A(FrameData[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__buf_8 input59 (.A(FrameData[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__buf_2 input6 (.A(E2END[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input60 (.A(FrameData[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net60));
 sky130_fd_sc_hd__buf_8 input61 (.A(FrameData[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net61));
 sky130_fd_sc_hd__buf_8 input62 (.A(FrameData[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net62));
 sky130_fd_sc_hd__buf_8 input63 (.A(FrameData[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net63));
 sky130_fd_sc_hd__buf_8 input64 (.A(FrameData[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net64));
 sky130_fd_sc_hd__buf_8 input65 (.A(FrameData[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net65));
 sky130_fd_sc_hd__buf_8 input66 (.A(FrameData[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net66));
 sky130_fd_sc_hd__buf_8 input67 (.A(FrameData[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net67));
 sky130_fd_sc_hd__buf_8 input68 (.A(FrameData[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net68));
 sky130_fd_sc_hd__buf_8 input69 (.A(FrameData[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net69));
 sky130_fd_sc_hd__buf_2 input7 (.A(E2END[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_8 input70 (.A(FrameData[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net70));
 sky130_fd_sc_hd__buf_8 input71 (.A(FrameData[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__buf_8 input72 (.A(FrameData[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__buf_8 input73 (.A(FrameData[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__buf_8 input74 (.A(FrameData[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__buf_8 input75 (.A(FrameData[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__buf_8 input76 (.A(FrameData[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_16 input77 (.A(FrameData[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__buf_8 input78 (.A(FrameData[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__buf_8 input79 (.A(FrameData[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(E2END[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input80 (.A(FrameData[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__buf_8 input81 (.A(FrameData[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__buf_8 input82 (.A(FrameStrobe[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_16 input83 (.A(FrameStrobe[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_16 input84 (.A(FrameStrobe[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_16 input85 (.A(FrameStrobe[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__buf_8 input86 (.A(FrameStrobe[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__buf_8 input87 (.A(FrameStrobe[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__buf_8 input88 (.A(FrameStrobe[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__buf_8 input89 (.A(FrameStrobe[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input9 (.A(E2END[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_8 input90 (.A(FrameStrobe[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__buf_8 input91 (.A(FrameStrobe[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__buf_8 input92 (.A(FrameStrobe[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_16 input93 (.A(FrameStrobe[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_16 input94 (.A(FrameStrobe[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_16 input95 (.A(FrameStrobe[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__buf_12 input96 (.A(FrameStrobe[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_16 input97 (.A(FrameStrobe[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_16 input98 (.A(FrameStrobe[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__buf_12 input99 (.A(FrameStrobe[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 inst_clk_buf (.A(UserCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net459));
 sky130_fd_sc_hd__buf_6 max_cap508 (.A(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net508));
 sky130_fd_sc_hd__buf_6 max_cap509 (.A(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net509));
 sky130_fd_sc_hd__buf_12 max_cap510 (.A(\Inst_LD_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_8 max_cap511 (.A(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net511));
 sky130_fd_sc_hd__buf_8 max_cap512 (.A(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_8 max_cap513 (.A(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net513));
 sky130_fd_sc_hd__buf_12 max_cap514 (.A(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net514));
 sky130_fd_sc_hd__buf_8 max_cap515 (.A(\Inst_LH_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net515));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(Co));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net257),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output266 (.A(net266),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output272 (.A(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output274 (.A(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output287 (.A(net287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output288 (.A(net288),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output292 (.A(net292),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output298 (.A(net298),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output301 (.A(net301),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output302 (.A(net302),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output305 (.A(net305),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output308 (.A(net308),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output312 (.A(net312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output314 (.A(net314),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output315 (.A(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__clkbuf_4 output317 (.A(net317),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output322 (.A(net322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output325 (.A(net325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output329 (.A(net329),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output345 (.A(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output357 (.A(net357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__buf_2 output366 (.A(net366),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output367 (.A(net367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output379 (.A(net379),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output393 (.A(net393),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output394 (.A(net394),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output395 (.A(net395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output397 (.A(net397),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output398 (.A(net398),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output399 (.A(net399),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net401),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output402 (.A(net402),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output403 (.A(net403),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output404 (.A(net404),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output407 (.A(net407),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output408 (.A(net408),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output410 (.A(net410),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output413 (.A(net413),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output414 (.A(net414),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output416 (.A(net416),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output417 (.A(net417),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output418 (.A(net418),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output420 (.A(net420),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output421 (.A(net421),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output424 (.A(net424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output425 (.A(net425),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output427 (.A(net427),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output428 (.A(net428),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output429 (.A(net429),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output430 (.A(net430),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output431 (.A(net431),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output432 (.A(net432),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output433 (.A(net433),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__buf_2 output434 (.A(net434),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output435 (.A(net435),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output436 (.A(net436),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output437 (.A(net437),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__buf_2 output438 (.A(net438),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output440 (.A(net440),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output441 (.A(net441),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output442 (.A(net442),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output443 (.A(net443),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output444 (.A(net444),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output445 (.A(net445),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output446 (.A(net446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output448 (.A(net448),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output449 (.A(net449),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output450 (.A(net450),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output451 (.A(net451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output452 (.A(net452),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output453 (.A(net453),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output454 (.A(net454),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output455 (.A(net455),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output456 (.A(net456),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output457 (.A(net457),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output458 (.A(net458),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output459 (.A(net459),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output460 (.A(net460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output461 (.A(net461),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output462 (.A(net462),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output463 (.A(net463),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output464 (.A(net464),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output465 (.A(net465),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output466 (.A(net466),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output467 (.A(net467),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output468 (.A(net468),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output469 (.A(net469),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output470 (.A(net470),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output471 (.A(net471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output472 (.A(net472),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output473 (.A(net473),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output474 (.A(net474),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output475 (.A(net475),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output476 (.A(net476),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output477 (.A(net477),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output478 (.A(net478),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output479 (.A(net479),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output480 (.A(net480),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output481 (.A(net481),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output482 (.A(net482),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output483 (.A(net483),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output484 (.A(net484),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output485 (.A(net485),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output486 (.A(net486),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output487 (.A(net487),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output488 (.A(net488),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output489 (.A(net489),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output490 (.A(net490),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output491 (.A(net491),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output492 (.A(net492),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output493 (.A(net493),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output494 (.A(net494),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output495 (.A(net495),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output496 (.A(net496),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output497 (.A(net497),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output498 (.A(net498),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output499 (.A(net499),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output500 (.A(net500),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output501 (.A(net501),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output502 (.A(net502),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output503 (.A(net503),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output504 (.A(net504),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output505 (.A(net505),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output506 (.A(net506),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output507 (.A(net507),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net538));
 sky130_fd_sc_hd__buf_1 rebuffer2 (.A(\Inst_LUT4AB_switch_matrix.JW2BEG5 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net533));
 sky130_fd_sc_hd__buf_6 rebuffer3 (.A(net536),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net534));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(\Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(\Inst_LUT4AB_switch_matrix.S0 ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net536));
 sky130_fd_sc_hd__buf_6 split1 (.A(\Inst_LB_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net532));
 sky130_fd_sc_hd__buf_6 split4 (.A(\Inst_LE_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net535));
 sky130_fd_sc_hd__buf_4 split5 (.A(\Inst_LG_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net540));
 sky130_fd_sc_hd__buf_6 split6 (.A(\Inst_LC_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net537));
 sky130_fd_sc_hd__buf_6 split7 (.A(\Inst_LF_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net541));
 sky130_fd_sc_hd__buf_4 split8 (.A(\Inst_LUT4AB_switch_matrix.M_AB ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net542));
 sky130_fd_sc_hd__buf_4 split9 (.A(\Inst_LA_LUT4c_frame_config_dffesr.O ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0._0_  (.A(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_1._0_  (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_10._0_  (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_11._0_  (.A(net84),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_12._0_  (.A(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_13._0_  (.A(net86),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_14._0_  (.A(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_15._0_  (.A(net88),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_16._0_  (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_17._0_  (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_18._0_  (.A(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_19._0_  (.A(net92),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2._0_  (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_3._0_  (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4._0_  (.A(net96),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_5._0_  (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_6._0_  (.A(net98),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_7._0_  (.A(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_8._0_  (.A(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_9._0_  (.A(net101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_inbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0._0_  (.A(\strobe_inbuf_0.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1._0_  (.A(\strobe_inbuf_1.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10._0_  (.A(\strobe_inbuf_10.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11._0_  (.A(\strobe_inbuf_11.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12._0_  (.A(\strobe_inbuf_12.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13._0_  (.A(\strobe_inbuf_13.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14._0_  (.A(\strobe_inbuf_14.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15._0_  (.A(\strobe_inbuf_15.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16._0_  (.A(\strobe_inbuf_16.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17._0_  (.A(\strobe_inbuf_17.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_18._0_  (.A(\strobe_inbuf_18.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19._0_  (.A(\strobe_inbuf_19.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_2._0_  (.A(\strobe_inbuf_2.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_3._0_  (.A(\strobe_inbuf_3.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_4._0_  (.A(\strobe_inbuf_4.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5._0_  (.A(\strobe_inbuf_5.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6._0_  (.A(\strobe_inbuf_6.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7._0_  (.A(\strobe_inbuf_7.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8._0_  (.A(\strobe_inbuf_8.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9._0_  (.A(\strobe_inbuf_9.X ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(\strobe_outbuf_9.X ));
endmodule
