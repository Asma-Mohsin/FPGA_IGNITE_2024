// This is the unpowered netlist.
module W_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire \Inst_A_IO_1_bidirectional_frame_config_pass.I ;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.O ;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_A_IO_1_bidirectional_frame_config_pass.T ;
 wire \Inst_A_config_Config_access.ConfigBits[0] ;
 wire \Inst_A_config_Config_access.ConfigBits[1] ;
 wire \Inst_A_config_Config_access.ConfigBits[2] ;
 wire \Inst_A_config_Config_access.ConfigBits[3] ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.I ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.O ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.T ;
 wire \Inst_B_config_Config_access.ConfigBits[0] ;
 wire \Inst_B_config_Config_access.ConfigBits[1] ;
 wire \Inst_B_config_Config_access.ConfigBits[2] ;
 wire \Inst_B_config_Config_access.ConfigBits[3] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[100] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[101] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[102] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[103] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[104] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[105] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[106] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[107] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[108] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[109] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[10] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[110] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[111] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[112] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[113] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[11] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[12] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[13] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[14] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[15] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[16] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[17] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[18] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[19] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[20] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[21] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[22] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[23] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[24] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[25] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[26] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[27] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[28] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[29] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[30] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[31] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[32] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[33] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[34] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[35] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[36] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[37] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[38] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[39] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[40] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[41] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[42] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[43] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[44] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[45] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[46] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[47] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[48] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[49] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[50] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[51] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[52] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[53] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[54] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[55] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[56] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[57] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[58] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[59] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[60] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[61] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[62] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[63] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[64] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[65] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[66] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[67] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[68] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[69] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[70] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[71] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[72] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[73] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[74] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[75] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[76] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[77] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[78] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[79] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[80] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[81] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[82] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[83] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[84] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[85] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[86] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[87] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[88] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[89] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[8] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[90] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[91] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[92] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[93] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[94] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[95] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[96] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[97] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[98] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[99] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits[9] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[0] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[100] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[101] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[102] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[103] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[104] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[105] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[106] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[107] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[108] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[109] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[10] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[110] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[111] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[112] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[113] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[11] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[12] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[13] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[14] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[15] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[16] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[17] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[18] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[19] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[1] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[20] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[21] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[22] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[23] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[24] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[25] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[26] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[27] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[28] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[29] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[2] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[30] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[31] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[32] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[33] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[34] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[35] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[36] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[37] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[38] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[39] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[3] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[40] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[41] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[42] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[43] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[44] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[45] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[46] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[47] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[48] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[49] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[4] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[50] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[51] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[52] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[53] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[54] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[55] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[56] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[57] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[58] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[59] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[5] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[60] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[61] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[62] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[63] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[64] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[65] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[66] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[67] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[68] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[69] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[6] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[70] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[71] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[72] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[73] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[74] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[75] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[76] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[77] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[78] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[79] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[7] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[80] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[81] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[82] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[83] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[84] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[85] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[86] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[87] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[88] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[89] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[8] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[90] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[91] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[92] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[93] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[94] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[95] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[96] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[97] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[98] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[99] ;
 wire \Inst_W_IO_ConfigMem.ConfigBits_N[9] ;
 wire \Inst_W_IO_switch_matrix.E1BEG0 ;
 wire \Inst_W_IO_switch_matrix.E1BEG1 ;
 wire \Inst_W_IO_switch_matrix.E1BEG2 ;
 wire \Inst_W_IO_switch_matrix.E1BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG0 ;
 wire \Inst_W_IO_switch_matrix.E2BEG1 ;
 wire \Inst_W_IO_switch_matrix.E2BEG2 ;
 wire \Inst_W_IO_switch_matrix.E2BEG3 ;
 wire \Inst_W_IO_switch_matrix.E2BEG4 ;
 wire \Inst_W_IO_switch_matrix.E2BEG5 ;
 wire \Inst_W_IO_switch_matrix.E2BEG6 ;
 wire \Inst_W_IO_switch_matrix.E2BEG7 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb0 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb1 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb2 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb3 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb4 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb5 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb6 ;
 wire \Inst_W_IO_switch_matrix.E2BEGb7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG0 ;
 wire \Inst_W_IO_switch_matrix.E6BEG1 ;
 wire \Inst_W_IO_switch_matrix.E6BEG10 ;
 wire \Inst_W_IO_switch_matrix.E6BEG11 ;
 wire \Inst_W_IO_switch_matrix.E6BEG2 ;
 wire \Inst_W_IO_switch_matrix.E6BEG3 ;
 wire \Inst_W_IO_switch_matrix.E6BEG4 ;
 wire \Inst_W_IO_switch_matrix.E6BEG5 ;
 wire \Inst_W_IO_switch_matrix.E6BEG6 ;
 wire \Inst_W_IO_switch_matrix.E6BEG7 ;
 wire \Inst_W_IO_switch_matrix.E6BEG8 ;
 wire \Inst_W_IO_switch_matrix.E6BEG9 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG0 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG1 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG10 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG11 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG12 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG13 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG14 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG15 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG2 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG3 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG4 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG5 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG6 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG7 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG8 ;
 wire \Inst_W_IO_switch_matrix.EE4BEG9 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out0 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out1 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out2 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out3 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out0 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out1 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out2 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out3 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN[0] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN[1] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._0_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._1_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN[0] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN[1] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._0_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._1_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN[0] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN[1] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._0_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._1_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN[0] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN[1] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._0_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._1_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A0 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A1 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN[0] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN[1] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._0_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._1_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A0 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A1 ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN[0] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN[1] ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._0_ ;
 wire \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._1_ ;
 wire \data_inbuf_0.X ;
 wire \data_inbuf_1.X ;
 wire \data_inbuf_10.X ;
 wire \data_inbuf_11.X ;
 wire \data_inbuf_12.X ;
 wire \data_inbuf_13.X ;
 wire \data_inbuf_14.X ;
 wire \data_inbuf_15.X ;
 wire \data_inbuf_16.X ;
 wire \data_inbuf_17.X ;
 wire \data_inbuf_18.X ;
 wire \data_inbuf_19.X ;
 wire \data_inbuf_2.X ;
 wire \data_inbuf_20.X ;
 wire \data_inbuf_21.X ;
 wire \data_inbuf_22.X ;
 wire \data_inbuf_23.X ;
 wire \data_inbuf_24.X ;
 wire \data_inbuf_25.X ;
 wire \data_inbuf_26.X ;
 wire \data_inbuf_27.X ;
 wire \data_inbuf_28.X ;
 wire \data_inbuf_29.X ;
 wire \data_inbuf_3.X ;
 wire \data_inbuf_30.X ;
 wire \data_inbuf_31.X ;
 wire \data_inbuf_4.X ;
 wire \data_inbuf_5.X ;
 wire \data_inbuf_6.X ;
 wire \data_inbuf_7.X ;
 wire \data_inbuf_8.X ;
 wire \data_inbuf_9.X ;
 wire \data_outbuf_0.X ;
 wire \data_outbuf_1.X ;
 wire \data_outbuf_10.X ;
 wire \data_outbuf_11.X ;
 wire \data_outbuf_12.X ;
 wire \data_outbuf_13.X ;
 wire \data_outbuf_14.X ;
 wire \data_outbuf_15.X ;
 wire \data_outbuf_16.X ;
 wire \data_outbuf_17.X ;
 wire \data_outbuf_18.X ;
 wire \data_outbuf_19.X ;
 wire \data_outbuf_2.X ;
 wire \data_outbuf_20.X ;
 wire \data_outbuf_21.X ;
 wire \data_outbuf_22.X ;
 wire \data_outbuf_23.X ;
 wire \data_outbuf_24.X ;
 wire \data_outbuf_25.X ;
 wire \data_outbuf_26.X ;
 wire \data_outbuf_27.X ;
 wire \data_outbuf_28.X ;
 wire \data_outbuf_29.X ;
 wire \data_outbuf_3.X ;
 wire \data_outbuf_30.X ;
 wire \data_outbuf_31.X ;
 wire \data_outbuf_4.X ;
 wire \data_outbuf_5.X ;
 wire \data_outbuf_6.X ;
 wire \data_outbuf_7.X ;
 wire \data_outbuf_8.X ;
 wire \data_outbuf_9.X ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \strobe_inbuf_0.X ;
 wire \strobe_inbuf_1.X ;
 wire \strobe_inbuf_10.X ;
 wire \strobe_inbuf_11.X ;
 wire \strobe_inbuf_12.X ;
 wire \strobe_inbuf_13.X ;
 wire \strobe_inbuf_14.X ;
 wire \strobe_inbuf_15.X ;
 wire \strobe_inbuf_16.X ;
 wire \strobe_inbuf_17.X ;
 wire \strobe_inbuf_18.X ;
 wire \strobe_inbuf_19.X ;
 wire \strobe_inbuf_2.X ;
 wire \strobe_inbuf_3.X ;
 wire \strobe_inbuf_4.X ;
 wire \strobe_inbuf_5.X ;
 wire \strobe_inbuf_6.X ;
 wire \strobe_inbuf_7.X ;
 wire \strobe_inbuf_8.X ;
 wire \strobe_inbuf_9.X ;
 wire \strobe_outbuf_0.X ;
 wire \strobe_outbuf_1.X ;
 wire \strobe_outbuf_10.X ;
 wire \strobe_outbuf_11.X ;
 wire \strobe_outbuf_12.X ;
 wire \strobe_outbuf_13.X ;
 wire \strobe_outbuf_14.X ;
 wire \strobe_outbuf_15.X ;
 wire \strobe_outbuf_16.X ;
 wire \strobe_outbuf_17.X ;
 wire \strobe_outbuf_18.X ;
 wire \strobe_outbuf_19.X ;
 wire \strobe_outbuf_2.X ;
 wire \strobe_outbuf_3.X ;
 wire \strobe_outbuf_4.X ;
 wire \strobe_outbuf_5.X ;
 wire \strobe_outbuf_6.X ;
 wire \strobe_outbuf_7.X ;
 wire \strobe_outbuf_8.X ;
 wire \strobe_outbuf_9.X ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\strobe_inbuf_17.X ));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_9 ();
 sky130_fd_sc_hd__inv_2 \Inst_A_IO_1_bidirectional_frame_config_pass._0_  (.A(\Inst_A_IO_1_bidirectional_frame_config_pass.T ),
    .Y(net104));
 sky130_fd_sc_hd__dfxtp_1 \Inst_A_IO_1_bidirectional_frame_config_pass._1_  (.CLK(UserCLK),
    .D(net1),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_IO_1_bidirectional_frame_config_pass._2_  (.A(\Inst_A_IO_1_bidirectional_frame_config_pass.I ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_2 \Inst_A_IO_1_bidirectional_frame_config_pass._3_  (.A(net1),
    .X(\Inst_A_IO_1_bidirectional_frame_config_pass.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access._0_  (.A(\Inst_A_config_Config_access.ConfigBits[0] ),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access._1_  (.A(\Inst_A_config_Config_access.ConfigBits[1] ),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access._2_  (.A(\Inst_A_config_Config_access.ConfigBits[2] ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 \Inst_A_config_Config_access._3_  (.A(\Inst_A_config_Config_access.ConfigBits[3] ),
    .X(net108));
 sky130_fd_sc_hd__inv_2 \Inst_B_IO_1_bidirectional_frame_config_pass._0_  (.A(\Inst_B_IO_1_bidirectional_frame_config_pass.T ),
    .Y(net110));
 sky130_fd_sc_hd__dfxtp_1 \Inst_B_IO_1_bidirectional_frame_config_pass._1_  (.CLK(UserCLK),
    .D(net2),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_IO_1_bidirectional_frame_config_pass._2_  (.A(\Inst_B_IO_1_bidirectional_frame_config_pass.I ),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 \Inst_B_IO_1_bidirectional_frame_config_pass._3_  (.A(net2),
    .X(\Inst_B_IO_1_bidirectional_frame_config_pass.O ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access._0_  (.A(\Inst_B_config_Config_access.ConfigBits[0] ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access._1_  (.A(\Inst_B_config_Config_access.ConfigBits[1] ),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access._2_  (.A(\Inst_B_config_Config_access.ConfigBits[2] ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 \Inst_B_config_Config_access._3_  (.A(\Inst_B_config_Config_access.ConfigBits[3] ),
    .X(net114));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit0  (.D(net3),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[82] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit1  (.D(net14),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[83] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit10  (.D(net4),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[92] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit11  (.D(net5),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[93] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit12  (.D(net6),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[94] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit13  (.D(net7),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[95] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit14  (.D(net8),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[96] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit15  (.D(net9),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[97] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit16  (.D(net10),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[98] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit17  (.D(net11),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[99] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit18  (.D(net12),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[100] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit19  (.D(net13),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[101] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit2  (.D(net25),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[84] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit20  (.D(net15),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[102] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit21  (.D(net16),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[103] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit22  (.D(net17),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[104] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit23  (.D(net18),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[105] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit24  (.D(net19),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[106] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit25  (.D(net20),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[107] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit26  (.D(net21),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[108] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit27  (.D(net22),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[109] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit28  (.D(net23),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[110] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit29  (.D(net24),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[111] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit3  (.D(net28),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[85] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit30  (.D(net26),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[112] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit31  (.D(net27),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[113] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit4  (.D(net29),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[86] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit5  (.D(net30),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[87] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit6  (.D(net31),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[88] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit7  (.D(net32),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[89] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit8  (.D(net33),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[90] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame0_bit9  (.D(net34),
    .GATE(net35),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[91] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit0  (.D(net3),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[50] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit1  (.D(net14),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[51] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit10  (.D(net4),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[60] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit11  (.D(net5),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[61] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit12  (.D(net6),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[62] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit13  (.D(net7),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[63] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit14  (.D(net8),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[64] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit15  (.D(net9),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[65] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit16  (.D(net10),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[66] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit17  (.D(net11),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[67] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit18  (.D(net12),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[68] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit19  (.D(net13),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[69] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit2  (.D(net25),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[52] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit20  (.D(net15),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[70] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit21  (.D(net16),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[71] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit22  (.D(net17),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[72] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit23  (.D(net18),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[73] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit24  (.D(net19),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[74] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit25  (.D(net20),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[75] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit26  (.D(net21),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[76] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit27  (.D(net22),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[77] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit28  (.D(net23),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[78] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit29  (.D(net24),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[79] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit3  (.D(net28),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[53] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit30  (.D(net26),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[80] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit31  (.D(net27),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[81] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit4  (.D(net29),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[54] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit5  (.D(net30),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[55] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit6  (.D(net31),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[56] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit7  (.D(net32),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[57] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit8  (.D(net33),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[58] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame1_bit9  (.D(net34),
    .GATE(net46),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[59] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit0  (.D(net3),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[18] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit1  (.D(net14),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[19] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit10  (.D(net4),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[28] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit11  (.D(net5),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[29] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit12  (.D(net6),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[30] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit13  (.D(net7),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[31] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit14  (.D(net8),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[32] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit15  (.D(net9),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[33] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit16  (.D(net10),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[34] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit17  (.D(net11),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[35] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit18  (.D(net12),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[36] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit19  (.D(net13),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[37] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit2  (.D(net25),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[20] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit20  (.D(net15),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[38] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit21  (.D(net16),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[39] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit22  (.D(net17),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[40] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit23  (.D(net18),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[41] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit24  (.D(net19),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[42] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit25  (.D(net20),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[43] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit26  (.D(net21),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[44] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit27  (.D(net22),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[45] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit28  (.D(net23),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[46] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit29  (.D(net24),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[47] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit3  (.D(net28),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[21] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit30  (.D(net26),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[48] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit31  (.D(net27),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[49] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit4  (.D(net29),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[22] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit5  (.D(net30),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[23] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit6  (.D(net31),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[24] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit7  (.D(net32),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[25] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit8  (.D(net33),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[26] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame2_bit9  (.D(net34),
    .GATE(net47),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[27] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit14  (.D(net8),
    .GATE(net48),
    .Q(\Inst_A_config_Config_access.ConfigBits[0] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit15  (.D(net9),
    .GATE(net48),
    .Q(\Inst_A_config_Config_access.ConfigBits[1] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit16  (.D(net10),
    .GATE(net48),
    .Q(\Inst_A_config_Config_access.ConfigBits[2] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit17  (.D(net11),
    .GATE(net48),
    .Q(\Inst_A_config_Config_access.ConfigBits[3] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit18  (.D(net12),
    .GATE(net48),
    .Q(\Inst_B_config_Config_access.ConfigBits[0] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit19  (.D(net13),
    .GATE(net48),
    .Q(\Inst_B_config_Config_access.ConfigBits[1] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit20  (.D(net15),
    .GATE(net48),
    .Q(\Inst_B_config_Config_access.ConfigBits[2] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit21  (.D(net16),
    .GATE(net48),
    .Q(\Inst_B_config_Config_access.ConfigBits[3] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit22  (.D(net17),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[8] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit23  (.D(net18),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[9] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit24  (.D(net19),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[10] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit25  (.D(net20),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[11] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit26  (.D(net21),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[12] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit27  (.D(net22),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[13] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit28  (.D(net23),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[14] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit29  (.D(net24),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[15] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit30  (.D(net26),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[16] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_W_IO_ConfigMem.Inst_frame3_bit31  (.D(net27),
    .GATE(net48),
    .Q(\Inst_W_IO_ConfigMem.ConfigBits[17] ),
    .Q_N(\Inst_W_IO_ConfigMem.ConfigBits_N[17] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst0  (.A0(net67),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[100] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst1  (.A0(net71),
    .A1(net72),
    .A2(net73),
    .A3(net74),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[100] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst2  (.A0(net59),
    .A1(net60),
    .A2(net61),
    .A3(net62),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[100] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst3  (.A0(net63),
    .A1(net64),
    .A2(net65),
    .A3(net66),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[100] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[101] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst4  (.A0(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out0 ),
    .A1(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out1 ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out2 ),
    .A3(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out3 ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[102] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[103] ),
    .X(\Inst_A_IO_1_bidirectional_frame_config_pass.I ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst0  (.A0(net67),
    .A1(net68),
    .A2(net69),
    .A3(net70),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[107] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst1  (.A0(net71),
    .A1(net72),
    .A2(net73),
    .A3(net74),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[107] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst2  (.A0(net59),
    .A1(net60),
    .A2(net61),
    .A3(net62),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[107] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst3  (.A0(net63),
    .A1(net64),
    .A2(net65),
    .A3(net66),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[107] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[108] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst4  (.A0(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out0 ),
    .A1(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out1 ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out2 ),
    .A3(\Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out3 ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[109] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[110] ),
    .X(\Inst_B_IO_1_bidirectional_frame_config_pass.I ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._2_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._3_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN[1] ),
    .B(\Inst_W_IO_ConfigMem.ConfigBits[8] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._4_  (.A1(\Inst_W_IO_ConfigMem.ConfigBits[8] ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._0_ ),
    .B1(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._1_ ),
    .Y(\Inst_W_IO_switch_matrix.E1BEG0 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.break_comb_loop_inst0._0_  (.A(net58),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.break_comb_loop_inst1._0_  (.A(\Inst_A_IO_1_bidirectional_frame_config_pass.O ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._2_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._3_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN[1] ),
    .B(\Inst_W_IO_ConfigMem.ConfigBits[9] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._4_  (.A1(\Inst_W_IO_ConfigMem.ConfigBits[9] ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._0_ ),
    .B1(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._1_ ),
    .Y(\Inst_W_IO_switch_matrix.E1BEG1 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.break_comb_loop_inst0._0_  (.A(net57),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.break_comb_loop_inst1._0_  (.A(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._2_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._3_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN[1] ),
    .B(\Inst_W_IO_ConfigMem.ConfigBits[10] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._4_  (.A1(\Inst_W_IO_ConfigMem.ConfigBits[10] ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._0_ ),
    .B1(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._1_ ),
    .Y(\Inst_W_IO_switch_matrix.E1BEG2 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.break_comb_loop_inst0._0_  (.A(net56),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.break_comb_loop_inst1._0_  (.A(\Inst_B_IO_1_bidirectional_frame_config_pass.O ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._2_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._3_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN[1] ),
    .B(\Inst_W_IO_ConfigMem.ConfigBits[11] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._4_  (.A1(\Inst_W_IO_ConfigMem.ConfigBits[11] ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._0_ ),
    .B1(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._1_ ),
    .Y(\Inst_W_IO_switch_matrix.E1BEG3 ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.break_comb_loop_inst0._0_  (.A(net55),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.break_comb_loop_inst1._0_  (.A(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG0  (.A0(net74),
    .A1(net100),
    .A2(net93),
    .A3(net84),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[12] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[13] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG1  (.A0(net73),
    .A1(net99),
    .A2(net92),
    .A3(net83),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[14] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[15] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG2  (.A0(net72),
    .A1(net98),
    .A2(net91),
    .A3(net82),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[16] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[17] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG3  (.A0(net71),
    .A1(net97),
    .A2(net90),
    .A3(net81),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[18] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[19] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG4  (.A0(net70),
    .A1(net96),
    .A2(net89),
    .A3(net80),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[20] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[21] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG5  (.A0(net69),
    .A1(net95),
    .A2(net88),
    .A3(net79),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[22] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[23] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG6  (.A0(net68),
    .A1(net94),
    .A2(net102),
    .A3(net78),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[24] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[25] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG7  (.A0(net67),
    .A1(net87),
    .A2(net101),
    .A3(net75),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[26] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[27] ),
    .X(\Inst_W_IO_switch_matrix.E2BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb0  (.A0(net66),
    .A1(net100),
    .A2(net93),
    .A3(net84),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[28] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[29] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb1  (.A0(net65),
    .A1(net99),
    .A2(net92),
    .A3(net83),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[30] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[31] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb2  (.A0(net64),
    .A1(net98),
    .A2(net91),
    .A3(net82),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[32] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[33] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb3  (.A0(net63),
    .A1(net97),
    .A2(net90),
    .A3(net81),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[34] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[35] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb4  (.A0(net62),
    .A1(net96),
    .A2(net89),
    .A3(net80),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[36] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[37] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb5  (.A0(net61),
    .A1(net95),
    .A2(net88),
    .A3(net79),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[38] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[39] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb6  (.A0(net60),
    .A1(net94),
    .A2(net102),
    .A3(net78),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[40] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[41] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb7  (.A0(net59),
    .A1(net87),
    .A2(net101),
    .A3(net75),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[42] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[43] ),
    .X(\Inst_W_IO_switch_matrix.E2BEGb7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG0  (.A0(net57),
    .A1(net89),
    .A2(net77),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[76] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[77] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG1  (.A0(net58),
    .A1(net88),
    .A2(net76),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[78] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[79] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG10  (.A0(net56),
    .A1(net94),
    .A2(net78),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[96] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[97] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG10 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG11  (.A0(net55),
    .A1(net87),
    .A2(net75),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[98] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[99] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG11 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG2  (.A0(net100),
    .A1(net93),
    .A2(net84),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[80] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[81] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG3  (.A0(net99),
    .A1(net92),
    .A2(net83),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[82] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[83] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG4  (.A0(net57),
    .A1(net96),
    .A2(net80),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[84] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[85] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG5  (.A0(net58),
    .A1(net95),
    .A2(net79),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[86] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[87] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG6  (.A0(net56),
    .A1(net102),
    .A2(net86),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[88] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[89] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG7  (.A0(net55),
    .A1(net101),
    .A2(net85),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[90] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[91] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG8  (.A0(net98),
    .A1(net91),
    .A2(net82),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[92] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[93] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG8 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG9  (.A0(net97),
    .A1(net90),
    .A2(net81),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[94] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[95] ),
    .X(\Inst_W_IO_switch_matrix.E6BEG9 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG0  (.A0(net75),
    .A1(net79),
    .A2(net81),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[44] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[45] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG1  (.A0(net83),
    .A1(net85),
    .A2(net76),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[46] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[47] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG10  (.A0(net75),
    .A1(net79),
    .A2(net81),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[64] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[65] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG10 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG11  (.A0(net83),
    .A1(net85),
    .A2(net76),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.O ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[66] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[67] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG11 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG12  (.A0(net78),
    .A1(net80),
    .A2(net82),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[68] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[69] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG12 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG13  (.A0(net84),
    .A1(net86),
    .A2(net77),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[70] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[71] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG13 ));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG14  (.A0(net67),
    .A1(net69),
    .A2(net71),
    .A3(net73),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[72] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[73] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG14 ));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG15  (.A0(net68),
    .A1(net70),
    .A2(net72),
    .A3(net74),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[74] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[75] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG15 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG2  (.A0(net78),
    .A1(net80),
    .A2(net82),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[48] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[49] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG3  (.A0(net84),
    .A1(net86),
    .A2(net77),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[50] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[51] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG4  (.A0(net59),
    .A1(net61),
    .A2(net63),
    .A3(net65),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[52] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[53] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG4 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG5  (.A0(net60),
    .A1(net62),
    .A2(net64),
    .A3(net66),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[54] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[55] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG5 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG6  (.A0(net67),
    .A1(net69),
    .A2(net71),
    .A3(net73),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[56] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[57] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG6 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG7  (.A0(net68),
    .A1(net70),
    .A2(net72),
    .A3(net74),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[58] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[59] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG7 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG8  (.A0(net81),
    .A1(net83),
    .A2(net85),
    .A3(net76),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[60] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[61] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG8 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG9  (.A0(net78),
    .A1(net80),
    .A2(net82),
    .A3(net84),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[62] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[63] ),
    .X(\Inst_W_IO_switch_matrix.EE4BEG9 ));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._2_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._3_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN[1] ),
    .B(\Inst_W_IO_ConfigMem.ConfigBits[106] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._4_  (.A1(\Inst_W_IO_ConfigMem.ConfigBits[106] ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._0_ ),
    .B1(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._1_ ),
    .Y(\Inst_A_IO_1_bidirectional_frame_config_pass.T ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A0 ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A1 ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst0  (.A0(net74),
    .A1(net59),
    .A2(net60),
    .A3(net61),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[104] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[105] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst1  (.A0(net62),
    .A1(net63),
    .A2(net216),
    .A3(net218),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[104] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[105] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst1_216  (.LO(net216));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst1_218  (.HI(net218));
 sky130_fd_sc_hd__inv_2 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._2_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN[0] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._3_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN[1] ),
    .B(\Inst_W_IO_ConfigMem.ConfigBits[113] ),
    .Y(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._4_  (.A1(\Inst_W_IO_ConfigMem.ConfigBits[113] ),
    .A2(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._0_ ),
    .B1(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._1_ ),
    .Y(\Inst_B_IO_1_bidirectional_frame_config_pass.T ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.break_comb_loop_inst0._0_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A0 ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.break_comb_loop_inst1._0_  (.A(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A1 ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst0  (.A0(net73),
    .A1(net74),
    .A2(net59),
    .A3(net63),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[111] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[112] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst1  (.A0(net64),
    .A1(net65),
    .A2(net217),
    .A3(net219),
    .S0(\Inst_W_IO_ConfigMem.ConfigBits[111] ),
    .S1(\Inst_W_IO_ConfigMem.ConfigBits[112] ),
    .X(\Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A1 ));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst1_217  (.LO(net217));
 sky130_fd_sc_hd__conb_1 \Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst1_219  (.HI(net219));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__clkbuf_1 _00_ (.A(\Inst_W_IO_switch_matrix.E1BEG0 ),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 _01_ (.A(\Inst_W_IO_switch_matrix.E1BEG1 ),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 _02_ (.A(\Inst_W_IO_switch_matrix.E1BEG2 ),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 _03_ (.A(\Inst_W_IO_switch_matrix.E1BEG3 ),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 _04_ (.A(\Inst_W_IO_switch_matrix.E2BEG0 ),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 _05_ (.A(\Inst_W_IO_switch_matrix.E2BEG1 ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(\Inst_W_IO_switch_matrix.E2BEG2 ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 _07_ (.A(\Inst_W_IO_switch_matrix.E2BEG3 ),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 _08_ (.A(\Inst_W_IO_switch_matrix.E2BEG4 ),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 _09_ (.A(\Inst_W_IO_switch_matrix.E2BEG5 ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _10_ (.A(\Inst_W_IO_switch_matrix.E2BEG6 ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 _11_ (.A(\Inst_W_IO_switch_matrix.E2BEG7 ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 _12_ (.A(\Inst_W_IO_switch_matrix.E2BEGb0 ),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _13_ (.A(\Inst_W_IO_switch_matrix.E2BEGb1 ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _14_ (.A(\Inst_W_IO_switch_matrix.E2BEGb2 ),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _15_ (.A(\Inst_W_IO_switch_matrix.E2BEGb3 ),
    .X(net130));
 sky130_fd_sc_hd__buf_1 _16_ (.A(\Inst_W_IO_switch_matrix.E2BEGb4 ),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _17_ (.A(\Inst_W_IO_switch_matrix.E2BEGb5 ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _18_ (.A(\Inst_W_IO_switch_matrix.E2BEGb6 ),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _19_ (.A(\Inst_W_IO_switch_matrix.E2BEGb7 ),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 _20_ (.A(\Inst_W_IO_switch_matrix.E6BEG0 ),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _21_ (.A(\Inst_W_IO_switch_matrix.E6BEG1 ),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _22_ (.A(\Inst_W_IO_switch_matrix.E6BEG2 ),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _23_ (.A(\Inst_W_IO_switch_matrix.E6BEG3 ),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _24_ (.A(\Inst_W_IO_switch_matrix.E6BEG4 ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _25_ (.A(\Inst_W_IO_switch_matrix.E6BEG5 ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _26_ (.A(\Inst_W_IO_switch_matrix.E6BEG6 ),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 _27_ (.A(\Inst_W_IO_switch_matrix.E6BEG7 ),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _28_ (.A(\Inst_W_IO_switch_matrix.E6BEG8 ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _29_ (.A(\Inst_W_IO_switch_matrix.E6BEG9 ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _30_ (.A(\Inst_W_IO_switch_matrix.E6BEG10 ),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _31_ (.A(\Inst_W_IO_switch_matrix.E6BEG11 ),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _32_ (.A(\Inst_W_IO_switch_matrix.EE4BEG0 ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _33_ (.A(\Inst_W_IO_switch_matrix.EE4BEG1 ),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _34_ (.A(\Inst_W_IO_switch_matrix.EE4BEG2 ),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _35_ (.A(\Inst_W_IO_switch_matrix.EE4BEG3 ),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _36_ (.A(\Inst_W_IO_switch_matrix.EE4BEG4 ),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _37_ (.A(\Inst_W_IO_switch_matrix.EE4BEG5 ),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _38_ (.A(\Inst_W_IO_switch_matrix.EE4BEG6 ),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _39_ (.A(\Inst_W_IO_switch_matrix.EE4BEG7 ),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _40_ (.A(\Inst_W_IO_switch_matrix.EE4BEG8 ),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _41_ (.A(\Inst_W_IO_switch_matrix.EE4BEG9 ),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _42_ (.A(\Inst_W_IO_switch_matrix.EE4BEG10 ),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _43_ (.A(\Inst_W_IO_switch_matrix.EE4BEG11 ),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _44_ (.A(\Inst_W_IO_switch_matrix.EE4BEG12 ),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _45_ (.A(\Inst_W_IO_switch_matrix.EE4BEG13 ),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _46_ (.A(\Inst_W_IO_switch_matrix.EE4BEG14 ),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _47_ (.A(\Inst_W_IO_switch_matrix.EE4BEG15 ),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _48_ (.A(\data_outbuf_0.X ),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _49_ (.A(\data_outbuf_1.X ),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _50_ (.A(\data_outbuf_2.X ),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _51_ (.A(\data_outbuf_3.X ),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 _52_ (.A(\data_outbuf_4.X ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 _53_ (.A(\data_outbuf_5.X ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 _54_ (.A(\data_outbuf_6.X ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 _55_ (.A(\data_outbuf_7.X ),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 _56_ (.A(\data_outbuf_8.X ),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 _57_ (.A(\data_outbuf_9.X ),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 _58_ (.A(\data_outbuf_10.X ),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _59_ (.A(\data_outbuf_11.X ),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _60_ (.A(\data_outbuf_12.X ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 _61_ (.A(\data_outbuf_13.X ),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 _62_ (.A(\data_outbuf_14.X ),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _63_ (.A(\data_outbuf_15.X ),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 _64_ (.A(\data_outbuf_16.X ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 _65_ (.A(\data_outbuf_17.X ),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 _66_ (.A(\data_outbuf_18.X ),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _67_ (.A(\data_outbuf_19.X ),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 _68_ (.A(\data_outbuf_20.X ),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _69_ (.A(\data_outbuf_21.X ),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 _70_ (.A(\data_outbuf_22.X ),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 _71_ (.A(\data_outbuf_23.X ),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 _72_ (.A(\data_outbuf_24.X ),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 _73_ (.A(\data_outbuf_25.X ),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _74_ (.A(\data_outbuf_26.X ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _75_ (.A(\data_outbuf_27.X ),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _76_ (.A(\data_outbuf_28.X ),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _77_ (.A(\data_outbuf_29.X ),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _78_ (.A(\data_outbuf_30.X ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _79_ (.A(\data_outbuf_31.X ),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 _80_ (.A(\strobe_outbuf_0.X ),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 _81_ (.A(\strobe_outbuf_1.X ),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_1 _82_ (.A(\strobe_outbuf_2.X ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 _83_ (.A(\strobe_outbuf_3.X ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 _84_ (.A(\strobe_outbuf_4.X ),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 _85_ (.A(\strobe_outbuf_5.X ),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 _86_ (.A(\strobe_outbuf_6.X ),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_1 _87_ (.A(\strobe_outbuf_7.X ),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 _88_ (.A(\strobe_outbuf_8.X ),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 _89_ (.A(\strobe_outbuf_9.X ),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 _90_ (.A(\strobe_outbuf_10.X ),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _91_ (.A(\strobe_outbuf_11.X ),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 _92_ (.A(\strobe_outbuf_12.X ),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _93_ (.A(\strobe_outbuf_13.X ),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 _94_ (.A(\strobe_outbuf_14.X ),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 _95_ (.A(\strobe_outbuf_15.X ),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 _96_ (.A(\strobe_outbuf_16.X ),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 _97_ (.A(\strobe_outbuf_17.X ),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 _98_ (.A(\strobe_outbuf_18.X ),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 _99_ (.A(\strobe_outbuf_19.X ),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_0._0_  (.A(net3),
    .X(\data_inbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_1._0_  (.A(net14),
    .X(\data_inbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_10._0_  (.A(net4),
    .X(\data_inbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11._0_  (.A(net5),
    .X(\data_inbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_12._0_  (.A(net6),
    .X(\data_inbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_13._0_  (.A(net7),
    .X(\data_inbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14._0_  (.A(net8),
    .X(\data_inbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_15._0_  (.A(net9),
    .X(\data_inbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_16._0_  (.A(net10),
    .X(\data_inbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_17._0_  (.A(net11),
    .X(\data_inbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18._0_  (.A(net12),
    .X(\data_inbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19._0_  (.A(net13),
    .X(\data_inbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_2._0_  (.A(net25),
    .X(\data_inbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20._0_  (.A(net15),
    .X(\data_inbuf_20.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_21._0_  (.A(net16),
    .X(\data_inbuf_21.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22._0_  (.A(net17),
    .X(\data_inbuf_22.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23._0_  (.A(net18),
    .X(\data_inbuf_23.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24._0_  (.A(net19),
    .X(\data_inbuf_24.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25._0_  (.A(net20),
    .X(\data_inbuf_25.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26._0_  (.A(net21),
    .X(\data_inbuf_26.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_27._0_  (.A(net22),
    .X(\data_inbuf_27.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_28._0_  (.A(net23),
    .X(\data_inbuf_28.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_29._0_  (.A(net24),
    .X(\data_inbuf_29.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_3._0_  (.A(net28),
    .X(\data_inbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_30._0_  (.A(net26),
    .X(\data_inbuf_30.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31._0_  (.A(net27),
    .X(\data_inbuf_31.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_4._0_  (.A(net29),
    .X(\data_inbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_5._0_  (.A(net30),
    .X(\data_inbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_6._0_  (.A(net31),
    .X(\data_inbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_7._0_  (.A(net32),
    .X(\data_inbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_8._0_  (.A(net33),
    .X(\data_inbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_9._0_  (.A(net34),
    .X(\data_inbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0._0_  (.A(\data_inbuf_0.X ),
    .X(\data_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1._0_  (.A(\data_inbuf_1.X ),
    .X(\data_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10._0_  (.A(\data_inbuf_10.X ),
    .X(\data_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11._0_  (.A(\data_inbuf_11.X ),
    .X(\data_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12._0_  (.A(\data_inbuf_12.X ),
    .X(\data_outbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13._0_  (.A(\data_inbuf_13.X ),
    .X(\data_outbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14._0_  (.A(\data_inbuf_14.X ),
    .X(\data_outbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15._0_  (.A(\data_inbuf_15.X ),
    .X(\data_outbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16._0_  (.A(\data_inbuf_16.X ),
    .X(\data_outbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17._0_  (.A(\data_inbuf_17.X ),
    .X(\data_outbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18._0_  (.A(\data_inbuf_18.X ),
    .X(\data_outbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19._0_  (.A(\data_inbuf_19.X ),
    .X(\data_outbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2._0_  (.A(\data_inbuf_2.X ),
    .X(\data_outbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20._0_  (.A(\data_inbuf_20.X ),
    .X(\data_outbuf_20.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21._0_  (.A(\data_inbuf_21.X ),
    .X(\data_outbuf_21.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22._0_  (.A(\data_inbuf_22.X ),
    .X(\data_outbuf_22.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23._0_  (.A(\data_inbuf_23.X ),
    .X(\data_outbuf_23.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24._0_  (.A(\data_inbuf_24.X ),
    .X(\data_outbuf_24.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25._0_  (.A(\data_inbuf_25.X ),
    .X(\data_outbuf_25.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26._0_  (.A(\data_inbuf_26.X ),
    .X(\data_outbuf_26.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27._0_  (.A(\data_inbuf_27.X ),
    .X(\data_outbuf_27.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28._0_  (.A(\data_inbuf_28.X ),
    .X(\data_outbuf_28.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29._0_  (.A(\data_inbuf_29.X ),
    .X(\data_outbuf_29.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3._0_  (.A(\data_inbuf_3.X ),
    .X(\data_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30._0_  (.A(\data_inbuf_30.X ),
    .X(\data_outbuf_30.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31._0_  (.A(\data_inbuf_31.X ),
    .X(\data_outbuf_31.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4._0_  (.A(\data_inbuf_4.X ),
    .X(\data_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5._0_  (.A(\data_inbuf_5.X ),
    .X(\data_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6._0_  (.A(\data_inbuf_6.X ),
    .X(\data_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7._0_  (.A(\data_inbuf_7.X ),
    .X(\data_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8._0_  (.A(\data_inbuf_8.X ),
    .X(\data_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9._0_  (.A(\data_inbuf_9.X ),
    .X(\data_outbuf_9.X ));
 sky130_fd_sc_hd__buf_1 input1 (.A(A_O_top),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(FrameData[16]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input100 (.A(WW4END[7]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(WW4END[8]),
    .X(net101));
 sky130_fd_sc_hd__dlymetal6s2s_1 input102 (.A(WW4END[9]),
    .X(net102));
 sky130_fd_sc_hd__buf_2 input11 (.A(FrameData[17]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(FrameData[18]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(FrameData[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(FrameData[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(FrameData[20]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(FrameData[21]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(FrameData[22]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(FrameData[23]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(FrameData[24]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(B_O_top),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(FrameData[25]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(FrameData[26]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(FrameData[27]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(FrameData[28]),
    .X(net23));
 sky130_fd_sc_hd__buf_2 input24 (.A(FrameData[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(FrameData[2]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(FrameData[30]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 input27 (.A(FrameData[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(FrameData[3]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(FrameData[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(FrameData[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(FrameData[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(FrameData[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(FrameData[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(FrameData[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(FrameData[9]),
    .X(net34));
 sky130_fd_sc_hd__buf_8 input35 (.A(FrameStrobe[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(FrameStrobe[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(FrameStrobe[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(FrameStrobe[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(FrameStrobe[13]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(FrameData[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(FrameStrobe[14]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(FrameStrobe[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(FrameStrobe[16]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(FrameStrobe[17]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(FrameStrobe[18]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(FrameStrobe[19]),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(FrameStrobe[1]),
    .X(net46));
 sky130_fd_sc_hd__buf_8 input47 (.A(FrameStrobe[2]),
    .X(net47));
 sky130_fd_sc_hd__buf_4 input48 (.A(FrameStrobe[3]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(FrameStrobe[4]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(FrameData[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(FrameStrobe[5]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(FrameStrobe[6]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(FrameStrobe[7]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(FrameStrobe[8]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(FrameStrobe[9]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(W1END[0]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(W1END[1]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(W1END[2]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(W1END[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(W2END[0]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(FrameData[12]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input60 (.A(W2END[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(W2END[2]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(W2END[3]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(W2END[4]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(W2END[5]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(W2END[6]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(W2END[7]),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 input67 (.A(W2MID[0]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(W2MID[1]),
    .X(net68));
 sky130_fd_sc_hd__dlymetal6s2s_1 input69 (.A(W2MID[2]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(FrameData[13]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input70 (.A(W2MID[3]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(W2MID[4]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(W2MID[5]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 input73 (.A(W2MID[6]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(W2MID[7]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(W6END[0]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(W6END[10]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(W6END[11]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(W6END[1]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(W6END[2]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(FrameData[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(W6END[3]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 input81 (.A(W6END[4]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(W6END[5]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(W6END[6]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(W6END[7]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(W6END[8]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(W6END[9]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(WW4END[0]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(WW4END[10]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(WW4END[11]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(FrameData[15]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input90 (.A(WW4END[12]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(WW4END[13]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(WW4END[14]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(WW4END[15]),
    .X(net93));
 sky130_fd_sc_hd__dlymetal6s2s_1 input94 (.A(WW4END[1]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(WW4END[2]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(WW4END[3]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(WW4END[4]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(WW4END[5]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(WW4END[6]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 inst_clk_buf (.A(UserCLK),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(A_I_top));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(A_T_top));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(A_config_C_bit0));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(A_config_C_bit1));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(A_config_C_bit2));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(A_config_C_bit3));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(B_I_top));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(B_T_top));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(B_config_C_bit0));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(B_config_C_bit1));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(B_config_C_bit2));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(B_config_C_bit3));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net115),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net116),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net122),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net140),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net142),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net143),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net144),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net146),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net147),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net148),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net157),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net158),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net163),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net164),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net165),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net166),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output167 (.A(net167),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net168),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net169),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net170),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net171),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output173 (.A(net173),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output174 (.A(net174),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output176 (.A(net176),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__clkbuf_4 output177 (.A(net177),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__clkbuf_4 output178 (.A(net178),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output182 (.A(net182),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output184 (.A(net184),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__clkbuf_4 output185 (.A(net185),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output186 (.A(net186),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output187 (.A(net187),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__clkbuf_4 output188 (.A(net188),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output191 (.A(net191),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output192 (.A(net192),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output194 (.A(net194),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output195 (.A(net195),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output197 (.A(net197),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output199 (.A(net199),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output201 (.A(net201),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output205 (.A(net205),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output207 (.A(net207),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_1 output215 (.A(net215),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0._0_  (.A(net35),
    .X(\strobe_inbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_1._0_  (.A(net46),
    .X(\strobe_inbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_10._0_  (.A(net36),
    .X(\strobe_inbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_11._0_  (.A(net37),
    .X(\strobe_inbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_12._0_  (.A(net38),
    .X(\strobe_inbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_13._0_  (.A(net39),
    .X(\strobe_inbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_14._0_  (.A(net40),
    .X(\strobe_inbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_15._0_  (.A(net41),
    .X(\strobe_inbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_16._0_  (.A(net42),
    .X(\strobe_inbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_17._0_  (.A(net43),
    .X(\strobe_inbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_18._0_  (.A(net44),
    .X(\strobe_inbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_19._0_  (.A(net45),
    .X(\strobe_inbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2._0_  (.A(net47),
    .X(\strobe_inbuf_2.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_3._0_  (.A(net48),
    .X(\strobe_inbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4._0_  (.A(net49),
    .X(\strobe_inbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_5._0_  (.A(net50),
    .X(\strobe_inbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_6._0_  (.A(net51),
    .X(\strobe_inbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_7._0_  (.A(net52),
    .X(\strobe_inbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_8._0_  (.A(net53),
    .X(\strobe_inbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_9._0_  (.A(net54),
    .X(\strobe_inbuf_9.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0._0_  (.A(\strobe_inbuf_0.X ),
    .X(\strobe_outbuf_0.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1._0_  (.A(\strobe_inbuf_1.X ),
    .X(\strobe_outbuf_1.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10._0_  (.A(\strobe_inbuf_10.X ),
    .X(\strobe_outbuf_10.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11._0_  (.A(\strobe_inbuf_11.X ),
    .X(\strobe_outbuf_11.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12._0_  (.A(\strobe_inbuf_12.X ),
    .X(\strobe_outbuf_12.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13._0_  (.A(\strobe_inbuf_13.X ),
    .X(\strobe_outbuf_13.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14._0_  (.A(\strobe_inbuf_14.X ),
    .X(\strobe_outbuf_14.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15._0_  (.A(\strobe_inbuf_15.X ),
    .X(\strobe_outbuf_15.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16._0_  (.A(\strobe_inbuf_16.X ),
    .X(\strobe_outbuf_16.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17._0_  (.A(\strobe_inbuf_17.X ),
    .X(\strobe_outbuf_17.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_18._0_  (.A(\strobe_inbuf_18.X ),
    .X(\strobe_outbuf_18.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19._0_  (.A(\strobe_inbuf_19.X ),
    .X(\strobe_outbuf_19.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_2._0_  (.A(\strobe_inbuf_2.X ),
    .X(\strobe_outbuf_2.X ));
 sky130_fd_sc_hd__buf_1 \strobe_outbuf_3._0_  (.A(\strobe_inbuf_3.X ),
    .X(\strobe_outbuf_3.X ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_outbuf_4._0_  (.A(\strobe_inbuf_4.X ),
    .X(\strobe_outbuf_4.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5._0_  (.A(\strobe_inbuf_5.X ),
    .X(\strobe_outbuf_5.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6._0_  (.A(\strobe_inbuf_6.X ),
    .X(\strobe_outbuf_6.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7._0_  (.A(\strobe_inbuf_7.X ),
    .X(\strobe_outbuf_7.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8._0_  (.A(\strobe_inbuf_8.X ),
    .X(\strobe_outbuf_8.X ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9._0_  (.A(\strobe_inbuf_9.X ),
    .X(\strobe_outbuf_9.X ));
endmodule

