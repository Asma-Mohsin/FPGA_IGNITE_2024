VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_IO
  CLASS BLOCK ;
  FOREIGN W_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 181.000 BY 250.000 ;
  PIN A_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.230 0.700 174.610 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.430 0.700 184.810 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.990 0.700 179.370 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.510 0.700 205.890 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.950 0.700 211.330 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.710 0.700 216.090 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.150 0.700 221.530 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.870 0.700 190.250 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.070 0.700 200.450 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.310 0.700 195.690 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.590 0.700 226.970 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.350 0.700 231.730 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.790 0.700 237.170 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.230 0.700 242.610 ;
    END
  END B_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 3.550 181.000 3.930 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 5.590 181.000 5.970 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 6.950 181.000 7.330 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 8.990 181.000 9.370 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 11.030 181.000 11.410 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 13.070 181.000 13.450 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 14.430 181.000 14.810 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 16.470 181.000 16.850 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 18.510 181.000 18.890 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 20.550 181.000 20.930 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 22.590 181.000 22.970 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 23.950 181.000 24.330 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 25.990 181.000 26.370 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 28.030 181.000 28.410 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 30.070 181.000 30.450 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 32.110 181.000 32.490 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 33.470 181.000 33.850 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 35.510 181.000 35.890 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 37.550 181.000 37.930 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 39.590 181.000 39.970 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 71.550 181.000 71.930 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 90.590 181.000 90.970 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 92.630 181.000 93.010 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 73.590 181.000 73.970 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 75.630 181.000 76.010 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 77.670 181.000 78.050 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 79.030 181.000 79.410 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 81.070 181.000 81.450 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 83.110 181.000 83.490 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 85.150 181.000 85.530 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 87.190 181.000 87.570 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 88.550 181.000 88.930 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 41.630 181.000 42.010 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 60.670 181.000 61.050 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 62.030 181.000 62.410 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 64.070 181.000 64.450 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 66.110 181.000 66.490 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 68.150 181.000 68.530 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 69.510 181.000 69.890 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 42.990 181.000 43.370 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 45.030 181.000 45.410 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 47.070 181.000 47.450 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 49.110 181.000 49.490 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 51.150 181.000 51.530 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 52.510 181.000 52.890 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 54.550 181.000 54.930 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 56.590 181.000 56.970 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 58.630 181.000 59.010 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.950 0.700 7.330 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.310 0.700 59.690 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.070 0.700 64.450 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.510 0.700 69.890 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.950 0.700 75.330 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.710 0.700 80.090 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.150 0.700 85.530 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.590 0.700 90.970 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.350 0.700 95.730 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.790 0.700 101.170 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.230 0.700 106.610 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.710 0.700 12.090 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.990 0.700 111.370 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.430 0.700 116.810 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.870 0.700 122.250 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.310 0.700 127.690 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.070 0.700 132.450 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.510 0.700 137.890 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.950 0.700 143.330 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.710 0.700 148.090 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.150 0.700 153.530 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.590 0.700 158.970 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.150 0.700 17.530 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.350 0.700 163.730 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.790 0.700 169.170 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.590 0.700 22.970 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.350 0.700 27.730 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.790 0.700 33.170 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.230 0.700 38.610 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.990 0.700 43.370 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.430 0.700 48.810 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.870 0.700 54.250 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 185.790 181.000 186.170 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 204.830 181.000 205.210 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 206.870 181.000 207.250 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 208.230 181.000 208.610 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 210.270 181.000 210.650 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 212.310 181.000 212.690 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 214.350 181.000 214.730 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 216.390 181.000 216.770 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 217.750 181.000 218.130 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 219.790 181.000 220.170 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 221.830 181.000 222.210 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 187.830 181.000 188.210 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 223.870 181.000 224.250 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 225.230 181.000 225.610 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 227.270 181.000 227.650 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 229.310 181.000 229.690 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 231.350 181.000 231.730 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 233.390 181.000 233.770 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 234.750 181.000 235.130 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 236.790 181.000 237.170 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 238.830 181.000 239.210 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 240.870 181.000 241.250 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 189.190 181.000 189.570 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 242.910 181.000 243.290 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 244.270 181.000 244.650 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 191.230 181.000 191.610 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 193.270 181.000 193.650 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 195.310 181.000 195.690 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 197.350 181.000 197.730 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 198.710 181.000 199.090 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 180.300 200.750 181.000 201.130 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 202.790 181.000 203.170 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 9.700 0.000 10.080 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 90.200 0.000 90.580 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 98.020 0.000 98.400 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 106.300 0.000 106.680 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 114.120 0.000 114.500 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 122.400 0.000 122.780 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 130.220 0.000 130.600 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 138.500 0.000 138.880 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 0.000 146.700 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 154.600 0.000 154.980 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 162.420 0.000 162.800 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.520 0.000 17.900 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 25.800 0.000 26.180 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 33.620 0.000 34.000 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.900 0.000 42.280 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 49.720 0.000 50.100 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 58.000 0.000 58.380 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 65.820 0.000 66.200 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.100 0.000 74.480 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 81.920 0.000 82.300 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.700 249.300 10.080 250.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.200 249.300 90.580 250.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.020 249.300 98.400 250.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.300 249.300 106.680 250.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.120 249.300 114.500 250.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.400 249.300 122.780 250.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.220 249.300 130.600 250.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.500 249.300 138.880 250.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 249.300 146.700 250.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.600 249.300 154.980 250.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.420 249.300 162.800 250.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.520 249.300 17.900 250.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.800 249.300 26.180 250.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 33.620 249.300 34.000 250.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.900 249.300 42.280 250.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 49.720 249.300 50.100 250.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 249.300 58.380 250.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.820 249.300 66.200 250.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.100 249.300 74.480 250.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 81.920 249.300 82.300 250.000 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 170.700 0.000 171.080 0.700 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 170.700 249.300 171.080 250.000 ;
    END
  END UserCLKo
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 94.670 181.000 95.050 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 96.710 181.000 97.090 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 98.070 181.000 98.450 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 100.110 181.000 100.490 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 117.110 181.000 117.490 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 119.150 181.000 119.530 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 121.190 181.000 121.570 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 123.230 181.000 123.610 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 124.590 181.000 124.970 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 126.630 181.000 127.010 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 128.670 181.000 129.050 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 130.710 181.000 131.090 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 102.150 181.000 102.530 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 104.190 181.000 104.570 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 106.230 181.000 106.610 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 107.590 181.000 107.970 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 109.630 181.000 110.010 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 111.670 181.000 112.050 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 113.710 181.000 114.090 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 115.750 181.000 116.130 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 162.670 181.000 163.050 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 181.710 181.000 182.090 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 183.750 181.000 184.130 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 164.710 181.000 165.090 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 166.750 181.000 167.130 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 168.790 181.000 169.170 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 170.150 181.000 170.530 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 172.190 181.000 172.570 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 174.230 181.000 174.610 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 176.270 181.000 176.650 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 178.310 181.000 178.690 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 179.670 181.000 180.050 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 132.750 181.000 133.130 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 151.790 181.000 152.170 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 153.150 181.000 153.530 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 155.190 181.000 155.570 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 157.230 181.000 157.610 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 159.270 181.000 159.650 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 161.310 181.000 161.690 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 134.110 181.000 134.490 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 136.150 181.000 136.530 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 138.190 181.000 138.570 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 140.230 181.000 140.610 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 142.270 181.000 142.650 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 143.630 181.000 144.010 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 145.670 181.000 146.050 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 147.710 181.000 148.090 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 149.750 181.000 150.130 ;
    END
  END WW4END[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.580 5.200 22.180 245.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 5.200 175.780 245.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 21.290 175.960 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 174.470 175.960 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.880 5.200 25.480 245.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 175.720 244.885 ;
      LAYER met1 ;
        RECT 3.750 3.440 177.490 246.120 ;
      LAYER met2 ;
        RECT 3.770 249.020 9.420 249.300 ;
        RECT 10.360 249.020 17.240 249.300 ;
        RECT 18.180 249.020 25.520 249.300 ;
        RECT 26.460 249.020 33.340 249.300 ;
        RECT 34.280 249.020 41.620 249.300 ;
        RECT 42.560 249.020 49.440 249.300 ;
        RECT 50.380 249.020 57.720 249.300 ;
        RECT 58.660 249.020 65.540 249.300 ;
        RECT 66.480 249.020 73.820 249.300 ;
        RECT 74.760 249.020 81.640 249.300 ;
        RECT 82.580 249.020 89.920 249.300 ;
        RECT 90.860 249.020 97.740 249.300 ;
        RECT 98.680 249.020 106.020 249.300 ;
        RECT 106.960 249.020 113.840 249.300 ;
        RECT 114.780 249.020 122.120 249.300 ;
        RECT 123.060 249.020 129.940 249.300 ;
        RECT 130.880 249.020 138.220 249.300 ;
        RECT 139.160 249.020 146.040 249.300 ;
        RECT 146.980 249.020 154.320 249.300 ;
        RECT 155.260 249.020 162.140 249.300 ;
        RECT 163.080 249.020 170.420 249.300 ;
        RECT 171.360 249.020 177.470 249.300 ;
        RECT 3.770 0.980 177.470 249.020 ;
        RECT 3.770 0.700 9.420 0.980 ;
        RECT 10.360 0.700 17.240 0.980 ;
        RECT 18.180 0.700 25.520 0.980 ;
        RECT 26.460 0.700 33.340 0.980 ;
        RECT 34.280 0.700 41.620 0.980 ;
        RECT 42.560 0.700 49.440 0.980 ;
        RECT 50.380 0.700 57.720 0.980 ;
        RECT 58.660 0.700 65.540 0.980 ;
        RECT 66.480 0.700 73.820 0.980 ;
        RECT 74.760 0.700 81.640 0.980 ;
        RECT 82.580 0.700 89.920 0.980 ;
        RECT 90.860 0.700 97.740 0.980 ;
        RECT 98.680 0.700 106.020 0.980 ;
        RECT 106.960 0.700 113.840 0.980 ;
        RECT 114.780 0.700 122.120 0.980 ;
        RECT 123.060 0.700 129.940 0.980 ;
        RECT 130.880 0.700 138.220 0.980 ;
        RECT 139.160 0.700 146.040 0.980 ;
        RECT 146.980 0.700 154.320 0.980 ;
        RECT 155.260 0.700 162.140 0.980 ;
        RECT 163.080 0.700 170.420 0.980 ;
        RECT 171.360 0.700 177.470 0.980 ;
      LAYER met3 ;
        RECT 0.700 243.870 179.900 244.965 ;
        RECT 0.700 243.690 180.300 243.870 ;
        RECT 0.700 243.010 179.900 243.690 ;
        RECT 1.100 242.510 179.900 243.010 ;
        RECT 1.100 241.830 180.300 242.510 ;
        RECT 0.700 241.650 180.300 241.830 ;
        RECT 0.700 240.470 179.900 241.650 ;
        RECT 0.700 239.610 180.300 240.470 ;
        RECT 0.700 238.430 179.900 239.610 ;
        RECT 0.700 237.570 180.300 238.430 ;
        RECT 1.100 236.390 179.900 237.570 ;
        RECT 0.700 235.530 180.300 236.390 ;
        RECT 0.700 234.350 179.900 235.530 ;
        RECT 0.700 234.170 180.300 234.350 ;
        RECT 0.700 232.990 179.900 234.170 ;
        RECT 0.700 232.130 180.300 232.990 ;
        RECT 1.100 230.950 179.900 232.130 ;
        RECT 0.700 230.090 180.300 230.950 ;
        RECT 0.700 228.910 179.900 230.090 ;
        RECT 0.700 228.050 180.300 228.910 ;
        RECT 0.700 227.370 179.900 228.050 ;
        RECT 1.100 226.870 179.900 227.370 ;
        RECT 1.100 226.190 180.300 226.870 ;
        RECT 0.700 226.010 180.300 226.190 ;
        RECT 0.700 224.830 179.900 226.010 ;
        RECT 0.700 224.650 180.300 224.830 ;
        RECT 0.700 223.470 179.900 224.650 ;
        RECT 0.700 222.610 180.300 223.470 ;
        RECT 0.700 221.930 179.900 222.610 ;
        RECT 1.100 221.430 179.900 221.930 ;
        RECT 1.100 220.750 180.300 221.430 ;
        RECT 0.700 220.570 180.300 220.750 ;
        RECT 0.700 219.390 179.900 220.570 ;
        RECT 0.700 218.530 180.300 219.390 ;
        RECT 0.700 217.350 179.900 218.530 ;
        RECT 0.700 217.170 180.300 217.350 ;
        RECT 0.700 216.490 179.900 217.170 ;
        RECT 1.100 215.990 179.900 216.490 ;
        RECT 1.100 215.310 180.300 215.990 ;
        RECT 0.700 215.130 180.300 215.310 ;
        RECT 0.700 213.950 179.900 215.130 ;
        RECT 0.700 213.090 180.300 213.950 ;
        RECT 0.700 211.910 179.900 213.090 ;
        RECT 0.700 211.730 180.300 211.910 ;
        RECT 1.100 211.050 180.300 211.730 ;
        RECT 1.100 210.550 179.900 211.050 ;
        RECT 0.700 209.870 179.900 210.550 ;
        RECT 0.700 209.010 180.300 209.870 ;
        RECT 0.700 207.830 179.900 209.010 ;
        RECT 0.700 207.650 180.300 207.830 ;
        RECT 0.700 206.470 179.900 207.650 ;
        RECT 0.700 206.290 180.300 206.470 ;
        RECT 1.100 205.610 180.300 206.290 ;
        RECT 1.100 205.110 179.900 205.610 ;
        RECT 0.700 204.430 179.900 205.110 ;
        RECT 0.700 203.570 180.300 204.430 ;
        RECT 0.700 202.390 179.900 203.570 ;
        RECT 0.700 201.530 180.300 202.390 ;
        RECT 0.700 200.850 179.900 201.530 ;
        RECT 1.100 200.350 179.900 200.850 ;
        RECT 1.100 199.670 180.300 200.350 ;
        RECT 0.700 199.490 180.300 199.670 ;
        RECT 0.700 198.310 179.900 199.490 ;
        RECT 0.700 198.130 180.300 198.310 ;
        RECT 0.700 196.950 179.900 198.130 ;
        RECT 0.700 196.090 180.300 196.950 ;
        RECT 1.100 194.910 179.900 196.090 ;
        RECT 0.700 194.050 180.300 194.910 ;
        RECT 0.700 192.870 179.900 194.050 ;
        RECT 0.700 192.010 180.300 192.870 ;
        RECT 0.700 190.830 179.900 192.010 ;
        RECT 0.700 190.650 180.300 190.830 ;
        RECT 1.100 189.970 180.300 190.650 ;
        RECT 1.100 189.470 179.900 189.970 ;
        RECT 0.700 188.790 179.900 189.470 ;
        RECT 0.700 188.610 180.300 188.790 ;
        RECT 0.700 187.430 179.900 188.610 ;
        RECT 0.700 186.570 180.300 187.430 ;
        RECT 0.700 185.390 179.900 186.570 ;
        RECT 0.700 185.210 180.300 185.390 ;
        RECT 1.100 184.530 180.300 185.210 ;
        RECT 1.100 184.030 179.900 184.530 ;
        RECT 0.700 183.350 179.900 184.030 ;
        RECT 0.700 182.490 180.300 183.350 ;
        RECT 0.700 181.310 179.900 182.490 ;
        RECT 0.700 180.450 180.300 181.310 ;
        RECT 0.700 179.770 179.900 180.450 ;
        RECT 1.100 179.270 179.900 179.770 ;
        RECT 1.100 179.090 180.300 179.270 ;
        RECT 1.100 178.590 179.900 179.090 ;
        RECT 0.700 177.910 179.900 178.590 ;
        RECT 0.700 177.050 180.300 177.910 ;
        RECT 0.700 175.870 179.900 177.050 ;
        RECT 0.700 175.010 180.300 175.870 ;
        RECT 1.100 173.830 179.900 175.010 ;
        RECT 0.700 172.970 180.300 173.830 ;
        RECT 0.700 171.790 179.900 172.970 ;
        RECT 0.700 170.930 180.300 171.790 ;
        RECT 0.700 169.750 179.900 170.930 ;
        RECT 0.700 169.570 180.300 169.750 ;
        RECT 1.100 168.390 179.900 169.570 ;
        RECT 0.700 167.530 180.300 168.390 ;
        RECT 0.700 166.350 179.900 167.530 ;
        RECT 0.700 165.490 180.300 166.350 ;
        RECT 0.700 164.310 179.900 165.490 ;
        RECT 0.700 164.130 180.300 164.310 ;
        RECT 1.100 163.450 180.300 164.130 ;
        RECT 1.100 162.950 179.900 163.450 ;
        RECT 0.700 162.270 179.900 162.950 ;
        RECT 0.700 162.090 180.300 162.270 ;
        RECT 0.700 160.910 179.900 162.090 ;
        RECT 0.700 160.050 180.300 160.910 ;
        RECT 0.700 159.370 179.900 160.050 ;
        RECT 1.100 158.870 179.900 159.370 ;
        RECT 1.100 158.190 180.300 158.870 ;
        RECT 0.700 158.010 180.300 158.190 ;
        RECT 0.700 156.830 179.900 158.010 ;
        RECT 0.700 155.970 180.300 156.830 ;
        RECT 0.700 154.790 179.900 155.970 ;
        RECT 0.700 153.930 180.300 154.790 ;
        RECT 1.100 152.750 179.900 153.930 ;
        RECT 0.700 152.570 180.300 152.750 ;
        RECT 0.700 151.390 179.900 152.570 ;
        RECT 0.700 150.530 180.300 151.390 ;
        RECT 0.700 149.350 179.900 150.530 ;
        RECT 0.700 148.490 180.300 149.350 ;
        RECT 1.100 147.310 179.900 148.490 ;
        RECT 0.700 146.450 180.300 147.310 ;
        RECT 0.700 145.270 179.900 146.450 ;
        RECT 0.700 144.410 180.300 145.270 ;
        RECT 0.700 143.730 179.900 144.410 ;
        RECT 1.100 143.230 179.900 143.730 ;
        RECT 1.100 143.050 180.300 143.230 ;
        RECT 1.100 142.550 179.900 143.050 ;
        RECT 0.700 141.870 179.900 142.550 ;
        RECT 0.700 141.010 180.300 141.870 ;
        RECT 0.700 139.830 179.900 141.010 ;
        RECT 0.700 138.970 180.300 139.830 ;
        RECT 0.700 138.290 179.900 138.970 ;
        RECT 1.100 137.790 179.900 138.290 ;
        RECT 1.100 137.110 180.300 137.790 ;
        RECT 0.700 136.930 180.300 137.110 ;
        RECT 0.700 135.750 179.900 136.930 ;
        RECT 0.700 134.890 180.300 135.750 ;
        RECT 0.700 133.710 179.900 134.890 ;
        RECT 0.700 133.530 180.300 133.710 ;
        RECT 0.700 132.850 179.900 133.530 ;
        RECT 1.100 132.350 179.900 132.850 ;
        RECT 1.100 131.670 180.300 132.350 ;
        RECT 0.700 131.490 180.300 131.670 ;
        RECT 0.700 130.310 179.900 131.490 ;
        RECT 0.700 129.450 180.300 130.310 ;
        RECT 0.700 128.270 179.900 129.450 ;
        RECT 0.700 128.090 180.300 128.270 ;
        RECT 1.100 127.410 180.300 128.090 ;
        RECT 1.100 126.910 179.900 127.410 ;
        RECT 0.700 126.230 179.900 126.910 ;
        RECT 0.700 125.370 180.300 126.230 ;
        RECT 0.700 124.190 179.900 125.370 ;
        RECT 0.700 124.010 180.300 124.190 ;
        RECT 0.700 122.830 179.900 124.010 ;
        RECT 0.700 122.650 180.300 122.830 ;
        RECT 1.100 121.970 180.300 122.650 ;
        RECT 1.100 121.470 179.900 121.970 ;
        RECT 0.700 120.790 179.900 121.470 ;
        RECT 0.700 119.930 180.300 120.790 ;
        RECT 0.700 118.750 179.900 119.930 ;
        RECT 0.700 117.890 180.300 118.750 ;
        RECT 0.700 117.210 179.900 117.890 ;
        RECT 1.100 116.710 179.900 117.210 ;
        RECT 1.100 116.530 180.300 116.710 ;
        RECT 1.100 116.030 179.900 116.530 ;
        RECT 0.700 115.350 179.900 116.030 ;
        RECT 0.700 114.490 180.300 115.350 ;
        RECT 0.700 113.310 179.900 114.490 ;
        RECT 0.700 112.450 180.300 113.310 ;
        RECT 0.700 111.770 179.900 112.450 ;
        RECT 1.100 111.270 179.900 111.770 ;
        RECT 1.100 110.590 180.300 111.270 ;
        RECT 0.700 110.410 180.300 110.590 ;
        RECT 0.700 109.230 179.900 110.410 ;
        RECT 0.700 108.370 180.300 109.230 ;
        RECT 0.700 107.190 179.900 108.370 ;
        RECT 0.700 107.010 180.300 107.190 ;
        RECT 1.100 105.830 179.900 107.010 ;
        RECT 0.700 104.970 180.300 105.830 ;
        RECT 0.700 103.790 179.900 104.970 ;
        RECT 0.700 102.930 180.300 103.790 ;
        RECT 0.700 101.750 179.900 102.930 ;
        RECT 0.700 101.570 180.300 101.750 ;
        RECT 1.100 100.890 180.300 101.570 ;
        RECT 1.100 100.390 179.900 100.890 ;
        RECT 0.700 99.710 179.900 100.390 ;
        RECT 0.700 98.850 180.300 99.710 ;
        RECT 0.700 97.670 179.900 98.850 ;
        RECT 0.700 97.490 180.300 97.670 ;
        RECT 0.700 96.310 179.900 97.490 ;
        RECT 0.700 96.130 180.300 96.310 ;
        RECT 1.100 95.450 180.300 96.130 ;
        RECT 1.100 94.950 179.900 95.450 ;
        RECT 0.700 94.270 179.900 94.950 ;
        RECT 0.700 93.410 180.300 94.270 ;
        RECT 0.700 92.230 179.900 93.410 ;
        RECT 0.700 91.370 180.300 92.230 ;
        RECT 1.100 90.190 179.900 91.370 ;
        RECT 0.700 89.330 180.300 90.190 ;
        RECT 0.700 88.150 179.900 89.330 ;
        RECT 0.700 87.970 180.300 88.150 ;
        RECT 0.700 86.790 179.900 87.970 ;
        RECT 0.700 85.930 180.300 86.790 ;
        RECT 1.100 84.750 179.900 85.930 ;
        RECT 0.700 83.890 180.300 84.750 ;
        RECT 0.700 82.710 179.900 83.890 ;
        RECT 0.700 81.850 180.300 82.710 ;
        RECT 0.700 80.670 179.900 81.850 ;
        RECT 0.700 80.490 180.300 80.670 ;
        RECT 1.100 79.810 180.300 80.490 ;
        RECT 1.100 79.310 179.900 79.810 ;
        RECT 0.700 78.630 179.900 79.310 ;
        RECT 0.700 78.450 180.300 78.630 ;
        RECT 0.700 77.270 179.900 78.450 ;
        RECT 0.700 76.410 180.300 77.270 ;
        RECT 0.700 75.730 179.900 76.410 ;
        RECT 1.100 75.230 179.900 75.730 ;
        RECT 1.100 74.550 180.300 75.230 ;
        RECT 0.700 74.370 180.300 74.550 ;
        RECT 0.700 73.190 179.900 74.370 ;
        RECT 0.700 72.330 180.300 73.190 ;
        RECT 0.700 71.150 179.900 72.330 ;
        RECT 0.700 70.290 180.300 71.150 ;
        RECT 1.100 69.110 179.900 70.290 ;
        RECT 0.700 68.930 180.300 69.110 ;
        RECT 0.700 67.750 179.900 68.930 ;
        RECT 0.700 66.890 180.300 67.750 ;
        RECT 0.700 65.710 179.900 66.890 ;
        RECT 0.700 64.850 180.300 65.710 ;
        RECT 1.100 63.670 179.900 64.850 ;
        RECT 0.700 62.810 180.300 63.670 ;
        RECT 0.700 61.630 179.900 62.810 ;
        RECT 0.700 61.450 180.300 61.630 ;
        RECT 0.700 60.270 179.900 61.450 ;
        RECT 0.700 60.090 180.300 60.270 ;
        RECT 1.100 59.410 180.300 60.090 ;
        RECT 1.100 58.910 179.900 59.410 ;
        RECT 0.700 58.230 179.900 58.910 ;
        RECT 0.700 57.370 180.300 58.230 ;
        RECT 0.700 56.190 179.900 57.370 ;
        RECT 0.700 55.330 180.300 56.190 ;
        RECT 0.700 54.650 179.900 55.330 ;
        RECT 1.100 54.150 179.900 54.650 ;
        RECT 1.100 53.470 180.300 54.150 ;
        RECT 0.700 53.290 180.300 53.470 ;
        RECT 0.700 52.110 179.900 53.290 ;
        RECT 0.700 51.930 180.300 52.110 ;
        RECT 0.700 50.750 179.900 51.930 ;
        RECT 0.700 49.890 180.300 50.750 ;
        RECT 0.700 49.210 179.900 49.890 ;
        RECT 1.100 48.710 179.900 49.210 ;
        RECT 1.100 48.030 180.300 48.710 ;
        RECT 0.700 47.850 180.300 48.030 ;
        RECT 0.700 46.670 179.900 47.850 ;
        RECT 0.700 45.810 180.300 46.670 ;
        RECT 0.700 44.630 179.900 45.810 ;
        RECT 0.700 43.770 180.300 44.630 ;
        RECT 1.100 42.590 179.900 43.770 ;
        RECT 0.700 42.410 180.300 42.590 ;
        RECT 0.700 41.230 179.900 42.410 ;
        RECT 0.700 40.370 180.300 41.230 ;
        RECT 0.700 39.190 179.900 40.370 ;
        RECT 0.700 39.010 180.300 39.190 ;
        RECT 1.100 38.330 180.300 39.010 ;
        RECT 1.100 37.830 179.900 38.330 ;
        RECT 0.700 37.150 179.900 37.830 ;
        RECT 0.700 36.290 180.300 37.150 ;
        RECT 0.700 35.110 179.900 36.290 ;
        RECT 0.700 34.250 180.300 35.110 ;
        RECT 0.700 33.570 179.900 34.250 ;
        RECT 1.100 33.070 179.900 33.570 ;
        RECT 1.100 32.890 180.300 33.070 ;
        RECT 1.100 32.390 179.900 32.890 ;
        RECT 0.700 31.710 179.900 32.390 ;
        RECT 0.700 30.850 180.300 31.710 ;
        RECT 0.700 29.670 179.900 30.850 ;
        RECT 0.700 28.810 180.300 29.670 ;
        RECT 0.700 28.130 179.900 28.810 ;
        RECT 1.100 27.630 179.900 28.130 ;
        RECT 1.100 26.950 180.300 27.630 ;
        RECT 0.700 26.770 180.300 26.950 ;
        RECT 0.700 25.590 179.900 26.770 ;
        RECT 0.700 24.730 180.300 25.590 ;
        RECT 0.700 23.550 179.900 24.730 ;
        RECT 0.700 23.370 180.300 23.550 ;
        RECT 1.100 22.190 179.900 23.370 ;
        RECT 0.700 21.330 180.300 22.190 ;
        RECT 0.700 20.150 179.900 21.330 ;
        RECT 0.700 19.290 180.300 20.150 ;
        RECT 0.700 18.110 179.900 19.290 ;
        RECT 0.700 17.930 180.300 18.110 ;
        RECT 1.100 17.250 180.300 17.930 ;
        RECT 1.100 16.750 179.900 17.250 ;
        RECT 0.700 16.070 179.900 16.750 ;
        RECT 0.700 15.210 180.300 16.070 ;
        RECT 0.700 14.030 179.900 15.210 ;
        RECT 0.700 13.850 180.300 14.030 ;
        RECT 0.700 12.670 179.900 13.850 ;
        RECT 0.700 12.490 180.300 12.670 ;
        RECT 1.100 11.810 180.300 12.490 ;
        RECT 1.100 11.310 179.900 11.810 ;
        RECT 0.700 10.630 179.900 11.310 ;
        RECT 0.700 9.770 180.300 10.630 ;
        RECT 0.700 8.590 179.900 9.770 ;
        RECT 0.700 7.730 180.300 8.590 ;
        RECT 1.100 6.550 179.900 7.730 ;
        RECT 0.700 6.370 180.300 6.550 ;
        RECT 0.700 5.190 179.900 6.370 ;
        RECT 0.700 4.330 180.300 5.190 ;
        RECT 0.700 3.575 179.900 4.330 ;
      LAYER met4 ;
        RECT 78.495 44.375 106.425 243.945 ;
  END
END W_IO
END LIBRARY

