magic
tech sky130A
magscale 1 2
timestamp 1732487376
<< obsli1 >>
rect 1104 1071 43516 43537
<< obsm1 >>
rect 14 348 44606 44260
<< metal2 >>
rect 4986 44463 5042 44623
rect 5262 44463 5318 44623
rect 5538 44463 5594 44623
rect 5814 44463 5870 44623
rect 6090 44463 6146 44623
rect 6366 44463 6422 44623
rect 6642 44463 6698 44623
rect 6918 44463 6974 44623
rect 7194 44463 7250 44623
rect 7470 44463 7526 44623
rect 7746 44463 7802 44623
rect 8022 44463 8078 44623
rect 8298 44463 8354 44623
rect 8574 44463 8630 44623
rect 8850 44463 8906 44623
rect 9126 44463 9182 44623
rect 9402 44463 9458 44623
rect 9678 44463 9734 44623
rect 9954 44463 10010 44623
rect 10230 44463 10286 44623
rect 10506 44463 10562 44623
rect 10782 44463 10838 44623
rect 11058 44463 11114 44623
rect 11334 44463 11390 44623
rect 11610 44463 11666 44623
rect 11886 44463 11942 44623
rect 12162 44463 12218 44623
rect 12438 44463 12494 44623
rect 12714 44463 12770 44623
rect 12990 44463 13046 44623
rect 13266 44463 13322 44623
rect 13542 44463 13598 44623
rect 13818 44463 13874 44623
rect 14094 44463 14150 44623
rect 14370 44463 14426 44623
rect 14646 44463 14702 44623
rect 14922 44463 14978 44623
rect 15198 44463 15254 44623
rect 15474 44463 15530 44623
rect 15750 44463 15806 44623
rect 16026 44463 16082 44623
rect 16302 44463 16358 44623
rect 16578 44463 16634 44623
rect 16854 44463 16910 44623
rect 17130 44463 17186 44623
rect 17406 44463 17462 44623
rect 17682 44463 17738 44623
rect 17958 44463 18014 44623
rect 18234 44463 18290 44623
rect 18510 44463 18566 44623
rect 18786 44463 18842 44623
rect 19062 44463 19118 44623
rect 19338 44463 19394 44623
rect 19614 44463 19670 44623
rect 19890 44463 19946 44623
rect 20166 44463 20222 44623
rect 20442 44463 20498 44623
rect 20718 44463 20774 44623
rect 20994 44463 21050 44623
rect 21270 44463 21326 44623
rect 21546 44463 21602 44623
rect 21822 44463 21878 44623
rect 22098 44463 22154 44623
rect 22374 44463 22430 44623
rect 22650 44463 22706 44623
rect 22926 44463 22982 44623
rect 23202 44463 23258 44623
rect 23478 44463 23534 44623
rect 23754 44463 23810 44623
rect 24030 44463 24086 44623
rect 24306 44463 24362 44623
rect 24582 44463 24638 44623
rect 24858 44463 24914 44623
rect 25134 44463 25190 44623
rect 25410 44463 25466 44623
rect 25686 44463 25742 44623
rect 25962 44463 26018 44623
rect 26238 44463 26294 44623
rect 26514 44463 26570 44623
rect 26790 44463 26846 44623
rect 27066 44463 27122 44623
rect 27342 44463 27398 44623
rect 27618 44463 27674 44623
rect 27894 44463 27950 44623
rect 28170 44463 28226 44623
rect 28446 44463 28502 44623
rect 28722 44463 28778 44623
rect 28998 44463 29054 44623
rect 29274 44463 29330 44623
rect 29550 44463 29606 44623
rect 29826 44463 29882 44623
rect 30102 44463 30158 44623
rect 30378 44463 30434 44623
rect 30654 44463 30710 44623
rect 30930 44463 30986 44623
rect 31206 44463 31262 44623
rect 31482 44463 31538 44623
rect 31758 44463 31814 44623
rect 32034 44463 32090 44623
rect 32310 44463 32366 44623
rect 32586 44463 32642 44623
rect 32862 44463 32918 44623
rect 33138 44463 33194 44623
rect 33414 44463 33470 44623
rect 33690 44463 33746 44623
rect 33966 44463 34022 44623
rect 34242 44463 34298 44623
rect 34518 44463 34574 44623
rect 34794 44463 34850 44623
rect 35070 44463 35126 44623
rect 35346 44463 35402 44623
rect 35622 44463 35678 44623
rect 35898 44463 35954 44623
rect 36174 44463 36230 44623
rect 36450 44463 36506 44623
rect 36726 44463 36782 44623
rect 37002 44463 37058 44623
rect 37278 44463 37334 44623
rect 37554 44463 37610 44623
rect 37830 44463 37886 44623
rect 38106 44463 38162 44623
rect 38382 44463 38438 44623
rect 38658 44463 38714 44623
rect 38934 44463 38990 44623
rect 39210 44463 39266 44623
rect 39486 44463 39542 44623
rect 4986 0 5042 160
rect 5262 0 5318 160
rect 5538 0 5594 160
rect 5814 0 5870 160
rect 6090 0 6146 160
rect 6366 0 6422 160
rect 6642 0 6698 160
rect 6918 0 6974 160
rect 7194 0 7250 160
rect 7470 0 7526 160
rect 7746 0 7802 160
rect 8022 0 8078 160
rect 8298 0 8354 160
rect 8574 0 8630 160
rect 8850 0 8906 160
rect 9126 0 9182 160
rect 9402 0 9458 160
rect 9678 0 9734 160
rect 9954 0 10010 160
rect 10230 0 10286 160
rect 10506 0 10562 160
rect 10782 0 10838 160
rect 11058 0 11114 160
rect 11334 0 11390 160
rect 11610 0 11666 160
rect 11886 0 11942 160
rect 12162 0 12218 160
rect 12438 0 12494 160
rect 12714 0 12770 160
rect 12990 0 13046 160
rect 13266 0 13322 160
rect 13542 0 13598 160
rect 13818 0 13874 160
rect 14094 0 14150 160
rect 14370 0 14426 160
rect 14646 0 14702 160
rect 14922 0 14978 160
rect 15198 0 15254 160
rect 15474 0 15530 160
rect 15750 0 15806 160
rect 16026 0 16082 160
rect 16302 0 16358 160
rect 16578 0 16634 160
rect 16854 0 16910 160
rect 17130 0 17186 160
rect 17406 0 17462 160
rect 17682 0 17738 160
rect 17958 0 18014 160
rect 18234 0 18290 160
rect 18510 0 18566 160
rect 18786 0 18842 160
rect 19062 0 19118 160
rect 19338 0 19394 160
rect 19614 0 19670 160
rect 19890 0 19946 160
rect 20166 0 20222 160
rect 20442 0 20498 160
rect 20718 0 20774 160
rect 20994 0 21050 160
rect 21270 0 21326 160
rect 21546 0 21602 160
rect 21822 0 21878 160
rect 22098 0 22154 160
rect 22374 0 22430 160
rect 22650 0 22706 160
rect 22926 0 22982 160
rect 23202 0 23258 160
rect 23478 0 23534 160
rect 23754 0 23810 160
rect 24030 0 24086 160
rect 24306 0 24362 160
rect 24582 0 24638 160
rect 24858 0 24914 160
rect 25134 0 25190 160
rect 25410 0 25466 160
rect 25686 0 25742 160
rect 25962 0 26018 160
rect 26238 0 26294 160
rect 26514 0 26570 160
rect 26790 0 26846 160
rect 27066 0 27122 160
rect 27342 0 27398 160
rect 27618 0 27674 160
rect 27894 0 27950 160
rect 28170 0 28226 160
rect 28446 0 28502 160
rect 28722 0 28778 160
rect 28998 0 29054 160
rect 29274 0 29330 160
rect 29550 0 29606 160
rect 29826 0 29882 160
rect 30102 0 30158 160
rect 30378 0 30434 160
rect 30654 0 30710 160
rect 30930 0 30986 160
rect 31206 0 31262 160
rect 31482 0 31538 160
rect 31758 0 31814 160
rect 32034 0 32090 160
rect 32310 0 32366 160
rect 32586 0 32642 160
rect 32862 0 32918 160
rect 33138 0 33194 160
rect 33414 0 33470 160
rect 33690 0 33746 160
rect 33966 0 34022 160
rect 34242 0 34298 160
rect 34518 0 34574 160
rect 34794 0 34850 160
rect 35070 0 35126 160
rect 35346 0 35402 160
rect 35622 0 35678 160
rect 35898 0 35954 160
rect 36174 0 36230 160
rect 36450 0 36506 160
rect 36726 0 36782 160
rect 37002 0 37058 160
rect 37278 0 37334 160
rect 37554 0 37610 160
rect 37830 0 37886 160
rect 38106 0 38162 160
rect 38382 0 38438 160
rect 38658 0 38714 160
rect 38934 0 38990 160
rect 39210 0 39266 160
rect 39486 0 39542 160
<< obsm2 >>
rect 20 44407 4930 44554
rect 5098 44407 5206 44554
rect 5374 44407 5482 44554
rect 5650 44407 5758 44554
rect 5926 44407 6034 44554
rect 6202 44407 6310 44554
rect 6478 44407 6586 44554
rect 6754 44407 6862 44554
rect 7030 44407 7138 44554
rect 7306 44407 7414 44554
rect 7582 44407 7690 44554
rect 7858 44407 7966 44554
rect 8134 44407 8242 44554
rect 8410 44407 8518 44554
rect 8686 44407 8794 44554
rect 8962 44407 9070 44554
rect 9238 44407 9346 44554
rect 9514 44407 9622 44554
rect 9790 44407 9898 44554
rect 10066 44407 10174 44554
rect 10342 44407 10450 44554
rect 10618 44407 10726 44554
rect 10894 44407 11002 44554
rect 11170 44407 11278 44554
rect 11446 44407 11554 44554
rect 11722 44407 11830 44554
rect 11998 44407 12106 44554
rect 12274 44407 12382 44554
rect 12550 44407 12658 44554
rect 12826 44407 12934 44554
rect 13102 44407 13210 44554
rect 13378 44407 13486 44554
rect 13654 44407 13762 44554
rect 13930 44407 14038 44554
rect 14206 44407 14314 44554
rect 14482 44407 14590 44554
rect 14758 44407 14866 44554
rect 15034 44407 15142 44554
rect 15310 44407 15418 44554
rect 15586 44407 15694 44554
rect 15862 44407 15970 44554
rect 16138 44407 16246 44554
rect 16414 44407 16522 44554
rect 16690 44407 16798 44554
rect 16966 44407 17074 44554
rect 17242 44407 17350 44554
rect 17518 44407 17626 44554
rect 17794 44407 17902 44554
rect 18070 44407 18178 44554
rect 18346 44407 18454 44554
rect 18622 44407 18730 44554
rect 18898 44407 19006 44554
rect 19174 44407 19282 44554
rect 19450 44407 19558 44554
rect 19726 44407 19834 44554
rect 20002 44407 20110 44554
rect 20278 44407 20386 44554
rect 20554 44407 20662 44554
rect 20830 44407 20938 44554
rect 21106 44407 21214 44554
rect 21382 44407 21490 44554
rect 21658 44407 21766 44554
rect 21934 44407 22042 44554
rect 22210 44407 22318 44554
rect 22486 44407 22594 44554
rect 22762 44407 22870 44554
rect 23038 44407 23146 44554
rect 23314 44407 23422 44554
rect 23590 44407 23698 44554
rect 23866 44407 23974 44554
rect 24142 44407 24250 44554
rect 24418 44407 24526 44554
rect 24694 44407 24802 44554
rect 24970 44407 25078 44554
rect 25246 44407 25354 44554
rect 25522 44407 25630 44554
rect 25798 44407 25906 44554
rect 26074 44407 26182 44554
rect 26350 44407 26458 44554
rect 26626 44407 26734 44554
rect 26902 44407 27010 44554
rect 27178 44407 27286 44554
rect 27454 44407 27562 44554
rect 27730 44407 27838 44554
rect 28006 44407 28114 44554
rect 28282 44407 28390 44554
rect 28558 44407 28666 44554
rect 28834 44407 28942 44554
rect 29110 44407 29218 44554
rect 29386 44407 29494 44554
rect 29662 44407 29770 44554
rect 29938 44407 30046 44554
rect 30214 44407 30322 44554
rect 30490 44407 30598 44554
rect 30766 44407 30874 44554
rect 31042 44407 31150 44554
rect 31318 44407 31426 44554
rect 31594 44407 31702 44554
rect 31870 44407 31978 44554
rect 32146 44407 32254 44554
rect 32422 44407 32530 44554
rect 32698 44407 32806 44554
rect 32974 44407 33082 44554
rect 33250 44407 33358 44554
rect 33526 44407 33634 44554
rect 33802 44407 33910 44554
rect 34078 44407 34186 44554
rect 34354 44407 34462 44554
rect 34630 44407 34738 44554
rect 34906 44407 35014 44554
rect 35182 44407 35290 44554
rect 35458 44407 35566 44554
rect 35734 44407 35842 44554
rect 36010 44407 36118 44554
rect 36286 44407 36394 44554
rect 36562 44407 36670 44554
rect 36838 44407 36946 44554
rect 37114 44407 37222 44554
rect 37390 44407 37498 44554
rect 37666 44407 37774 44554
rect 37942 44407 38050 44554
rect 38218 44407 38326 44554
rect 38494 44407 38602 44554
rect 38770 44407 38878 44554
rect 39046 44407 39154 44554
rect 39322 44407 39430 44554
rect 39598 44407 44600 44554
rect 20 216 44600 44407
rect 20 31 4930 216
rect 5098 31 5206 216
rect 5374 31 5482 216
rect 5650 31 5758 216
rect 5926 31 6034 216
rect 6202 31 6310 216
rect 6478 31 6586 216
rect 6754 31 6862 216
rect 7030 31 7138 216
rect 7306 31 7414 216
rect 7582 31 7690 216
rect 7858 31 7966 216
rect 8134 31 8242 216
rect 8410 31 8518 216
rect 8686 31 8794 216
rect 8962 31 9070 216
rect 9238 31 9346 216
rect 9514 31 9622 216
rect 9790 31 9898 216
rect 10066 31 10174 216
rect 10342 31 10450 216
rect 10618 31 10726 216
rect 10894 31 11002 216
rect 11170 31 11278 216
rect 11446 31 11554 216
rect 11722 31 11830 216
rect 11998 31 12106 216
rect 12274 31 12382 216
rect 12550 31 12658 216
rect 12826 31 12934 216
rect 13102 31 13210 216
rect 13378 31 13486 216
rect 13654 31 13762 216
rect 13930 31 14038 216
rect 14206 31 14314 216
rect 14482 31 14590 216
rect 14758 31 14866 216
rect 15034 31 15142 216
rect 15310 31 15418 216
rect 15586 31 15694 216
rect 15862 31 15970 216
rect 16138 31 16246 216
rect 16414 31 16522 216
rect 16690 31 16798 216
rect 16966 31 17074 216
rect 17242 31 17350 216
rect 17518 31 17626 216
rect 17794 31 17902 216
rect 18070 31 18178 216
rect 18346 31 18454 216
rect 18622 31 18730 216
rect 18898 31 19006 216
rect 19174 31 19282 216
rect 19450 31 19558 216
rect 19726 31 19834 216
rect 20002 31 20110 216
rect 20278 31 20386 216
rect 20554 31 20662 216
rect 20830 31 20938 216
rect 21106 31 21214 216
rect 21382 31 21490 216
rect 21658 31 21766 216
rect 21934 31 22042 216
rect 22210 31 22318 216
rect 22486 31 22594 216
rect 22762 31 22870 216
rect 23038 31 23146 216
rect 23314 31 23422 216
rect 23590 31 23698 216
rect 23866 31 23974 216
rect 24142 31 24250 216
rect 24418 31 24526 216
rect 24694 31 24802 216
rect 24970 31 25078 216
rect 25246 31 25354 216
rect 25522 31 25630 216
rect 25798 31 25906 216
rect 26074 31 26182 216
rect 26350 31 26458 216
rect 26626 31 26734 216
rect 26902 31 27010 216
rect 27178 31 27286 216
rect 27454 31 27562 216
rect 27730 31 27838 216
rect 28006 31 28114 216
rect 28282 31 28390 216
rect 28558 31 28666 216
rect 28834 31 28942 216
rect 29110 31 29218 216
rect 29386 31 29494 216
rect 29662 31 29770 216
rect 29938 31 30046 216
rect 30214 31 30322 216
rect 30490 31 30598 216
rect 30766 31 30874 216
rect 31042 31 31150 216
rect 31318 31 31426 216
rect 31594 31 31702 216
rect 31870 31 31978 216
rect 32146 31 32254 216
rect 32422 31 32530 216
rect 32698 31 32806 216
rect 32974 31 33082 216
rect 33250 31 33358 216
rect 33526 31 33634 216
rect 33802 31 33910 216
rect 34078 31 34186 216
rect 34354 31 34462 216
rect 34630 31 34738 216
rect 34906 31 35014 216
rect 35182 31 35290 216
rect 35458 31 35566 216
rect 35734 31 35842 216
rect 36010 31 36118 216
rect 36286 31 36394 216
rect 36562 31 36670 216
rect 36838 31 36946 216
rect 37114 31 37222 216
rect 37390 31 37498 216
rect 37666 31 37774 216
rect 37942 31 38050 216
rect 38218 31 38326 216
rect 38494 31 38602 216
rect 38770 31 38878 216
rect 39046 31 39154 216
rect 39322 31 39430 216
rect 39598 31 44600 216
<< metal3 >>
rect 0 39448 160 39568
rect 0 39176 160 39296
rect 0 38904 160 39024
rect 0 38632 160 38752
rect 0 38360 160 38480
rect 0 38088 160 38208
rect 0 37816 160 37936
rect 0 37544 160 37664
rect 0 37272 160 37392
rect 0 37000 160 37120
rect 0 36728 160 36848
rect 0 36456 160 36576
rect 0 36184 160 36304
rect 0 35912 160 36032
rect 0 35640 160 35760
rect 0 35368 160 35488
rect 0 35096 160 35216
rect 0 34824 160 34944
rect 0 34552 160 34672
rect 0 34280 160 34400
rect 0 34008 160 34128
rect 0 33736 160 33856
rect 0 33464 160 33584
rect 0 33192 160 33312
rect 0 32920 160 33040
rect 0 32648 160 32768
rect 0 32376 160 32496
rect 0 32104 160 32224
rect 0 31832 160 31952
rect 0 31560 160 31680
rect 0 31288 160 31408
rect 0 31016 160 31136
rect 0 30744 160 30864
rect 0 30472 160 30592
rect 0 30200 160 30320
rect 0 29928 160 30048
rect 0 29656 160 29776
rect 0 29384 160 29504
rect 0 29112 160 29232
rect 0 28840 160 28960
rect 0 28568 160 28688
rect 0 28296 160 28416
rect 0 28024 160 28144
rect 0 27752 160 27872
rect 0 27480 160 27600
rect 0 27208 160 27328
rect 0 26936 160 27056
rect 0 26664 160 26784
rect 0 26392 160 26512
rect 0 26120 160 26240
rect 0 25848 160 25968
rect 0 25576 160 25696
rect 0 25304 160 25424
rect 0 25032 160 25152
rect 0 24760 160 24880
rect 0 24488 160 24608
rect 0 24216 160 24336
rect 0 23944 160 24064
rect 0 23672 160 23792
rect 0 23400 160 23520
rect 0 23128 160 23248
rect 0 22856 160 22976
rect 0 22584 160 22704
rect 0 22312 160 22432
rect 0 22040 160 22160
rect 0 21768 160 21888
rect 0 21496 160 21616
rect 0 21224 160 21344
rect 0 20952 160 21072
rect 0 20680 160 20800
rect 0 20408 160 20528
rect 0 20136 160 20256
rect 0 19864 160 19984
rect 0 19592 160 19712
rect 0 19320 160 19440
rect 0 19048 160 19168
rect 0 18776 160 18896
rect 0 18504 160 18624
rect 0 18232 160 18352
rect 0 17960 160 18080
rect 0 17688 160 17808
rect 0 17416 160 17536
rect 0 17144 160 17264
rect 0 16872 160 16992
rect 0 16600 160 16720
rect 0 16328 160 16448
rect 0 16056 160 16176
rect 0 15784 160 15904
rect 0 15512 160 15632
rect 0 15240 160 15360
rect 0 14968 160 15088
rect 0 14696 160 14816
rect 0 14424 160 14544
rect 0 14152 160 14272
rect 0 13880 160 14000
rect 0 13608 160 13728
rect 0 13336 160 13456
rect 0 13064 160 13184
rect 0 12792 160 12912
rect 0 12520 160 12640
rect 0 12248 160 12368
rect 0 11976 160 12096
rect 0 11704 160 11824
rect 0 11432 160 11552
rect 0 11160 160 11280
rect 0 10888 160 11008
rect 0 10616 160 10736
rect 0 10344 160 10464
rect 0 10072 160 10192
rect 0 9800 160 9920
rect 0 9528 160 9648
rect 0 9256 160 9376
rect 0 8984 160 9104
rect 0 8712 160 8832
rect 0 8440 160 8560
rect 0 8168 160 8288
rect 0 7896 160 8016
rect 0 7624 160 7744
rect 0 7352 160 7472
rect 0 7080 160 7200
rect 0 6808 160 6928
rect 0 6536 160 6656
rect 0 6264 160 6384
rect 0 5992 160 6112
rect 0 5720 160 5840
rect 0 5448 160 5568
rect 0 5176 160 5296
rect 0 4904 160 5024
rect 44495 39448 44655 39568
rect 44495 39176 44655 39296
rect 44495 38904 44655 39024
rect 44495 38632 44655 38752
rect 44495 38360 44655 38480
rect 44495 38088 44655 38208
rect 44495 37816 44655 37936
rect 44495 37544 44655 37664
rect 44495 37272 44655 37392
rect 44495 37000 44655 37120
rect 44495 36728 44655 36848
rect 44495 36456 44655 36576
rect 44495 36184 44655 36304
rect 44495 35912 44655 36032
rect 44495 35640 44655 35760
rect 44495 35368 44655 35488
rect 44495 35096 44655 35216
rect 44495 34824 44655 34944
rect 44495 34552 44655 34672
rect 44495 34280 44655 34400
rect 44495 34008 44655 34128
rect 44495 33736 44655 33856
rect 44495 33464 44655 33584
rect 44495 33192 44655 33312
rect 44495 32920 44655 33040
rect 44495 32648 44655 32768
rect 44495 32376 44655 32496
rect 44495 32104 44655 32224
rect 44495 31832 44655 31952
rect 44495 31560 44655 31680
rect 44495 31288 44655 31408
rect 44495 31016 44655 31136
rect 44495 30744 44655 30864
rect 44495 30472 44655 30592
rect 44495 30200 44655 30320
rect 44495 29928 44655 30048
rect 44495 29656 44655 29776
rect 44495 29384 44655 29504
rect 44495 29112 44655 29232
rect 44495 28840 44655 28960
rect 44495 28568 44655 28688
rect 44495 28296 44655 28416
rect 44495 28024 44655 28144
rect 44495 27752 44655 27872
rect 44495 27480 44655 27600
rect 44495 27208 44655 27328
rect 44495 26936 44655 27056
rect 44495 26664 44655 26784
rect 44495 26392 44655 26512
rect 44495 26120 44655 26240
rect 44495 25848 44655 25968
rect 44495 25576 44655 25696
rect 44495 25304 44655 25424
rect 44495 25032 44655 25152
rect 44495 24760 44655 24880
rect 44495 24488 44655 24608
rect 44495 24216 44655 24336
rect 44495 23944 44655 24064
rect 44495 23672 44655 23792
rect 44495 23400 44655 23520
rect 44495 23128 44655 23248
rect 44495 22856 44655 22976
rect 44495 22584 44655 22704
rect 44495 22312 44655 22432
rect 44495 22040 44655 22160
rect 44495 21768 44655 21888
rect 44495 21496 44655 21616
rect 44495 21224 44655 21344
rect 44495 20952 44655 21072
rect 44495 20680 44655 20800
rect 44495 20408 44655 20528
rect 44495 20136 44655 20256
rect 44495 19864 44655 19984
rect 44495 19592 44655 19712
rect 44495 19320 44655 19440
rect 44495 19048 44655 19168
rect 44495 18776 44655 18896
rect 44495 18504 44655 18624
rect 44495 18232 44655 18352
rect 44495 17960 44655 18080
rect 44495 17688 44655 17808
rect 44495 17416 44655 17536
rect 44495 17144 44655 17264
rect 44495 16872 44655 16992
rect 44495 16600 44655 16720
rect 44495 16328 44655 16448
rect 44495 16056 44655 16176
rect 44495 15784 44655 15904
rect 44495 15512 44655 15632
rect 44495 15240 44655 15360
rect 44495 14968 44655 15088
rect 44495 14696 44655 14816
rect 44495 14424 44655 14544
rect 44495 14152 44655 14272
rect 44495 13880 44655 14000
rect 44495 13608 44655 13728
rect 44495 13336 44655 13456
rect 44495 13064 44655 13184
rect 44495 12792 44655 12912
rect 44495 12520 44655 12640
rect 44495 12248 44655 12368
rect 44495 11976 44655 12096
rect 44495 11704 44655 11824
rect 44495 11432 44655 11552
rect 44495 11160 44655 11280
rect 44495 10888 44655 11008
rect 44495 10616 44655 10736
rect 44495 10344 44655 10464
rect 44495 10072 44655 10192
rect 44495 9800 44655 9920
rect 44495 9528 44655 9648
rect 44495 9256 44655 9376
rect 44495 8984 44655 9104
rect 44495 8712 44655 8832
rect 44495 8440 44655 8560
rect 44495 8168 44655 8288
rect 44495 7896 44655 8016
rect 44495 7624 44655 7744
rect 44495 7352 44655 7472
rect 44495 7080 44655 7200
rect 44495 6808 44655 6928
rect 44495 6536 44655 6656
rect 44495 6264 44655 6384
rect 44495 5992 44655 6112
rect 44495 5720 44655 5840
rect 44495 5448 44655 5568
rect 44495 5176 44655 5296
rect 44495 4904 44655 5024
<< obsm3 >>
rect 160 39648 44495 43621
rect 240 4824 44415 39648
rect 160 35 44495 4824
<< metal4 >>
rect 4208 1040 4528 43568
rect 19568 1040 19888 43568
rect 34928 1040 35248 43568
<< obsm4 >>
rect 611 960 4128 43621
rect 4608 960 19488 43621
rect 19968 960 34848 43621
rect 35328 960 43365 43621
rect 611 35 43365 960
<< obsm5 >>
rect 2140 860 43308 42660
<< labels >>
rlabel metal2 s 33966 0 34022 160 6 Ci
port 1 nsew signal input
rlabel metal2 s 33966 44463 34022 44623 6 Co
port 2 nsew signal output
rlabel metal3 s 44495 17960 44655 18080 6 E1BEG[0]
port 3 nsew signal output
rlabel metal3 s 44495 18232 44655 18352 6 E1BEG[1]
port 4 nsew signal output
rlabel metal3 s 44495 18504 44655 18624 6 E1BEG[2]
port 5 nsew signal output
rlabel metal3 s 44495 18776 44655 18896 6 E1BEG[3]
port 6 nsew signal output
rlabel metal3 s 0 17960 160 18080 6 E1END[0]
port 7 nsew signal input
rlabel metal3 s 0 18232 160 18352 6 E1END[1]
port 8 nsew signal input
rlabel metal3 s 0 18504 160 18624 6 E1END[2]
port 9 nsew signal input
rlabel metal3 s 0 18776 160 18896 6 E1END[3]
port 10 nsew signal input
rlabel metal3 s 44495 19048 44655 19168 6 E2BEG[0]
port 11 nsew signal output
rlabel metal3 s 44495 19320 44655 19440 6 E2BEG[1]
port 12 nsew signal output
rlabel metal3 s 44495 19592 44655 19712 6 E2BEG[2]
port 13 nsew signal output
rlabel metal3 s 44495 19864 44655 19984 6 E2BEG[3]
port 14 nsew signal output
rlabel metal3 s 44495 20136 44655 20256 6 E2BEG[4]
port 15 nsew signal output
rlabel metal3 s 44495 20408 44655 20528 6 E2BEG[5]
port 16 nsew signal output
rlabel metal3 s 44495 20680 44655 20800 6 E2BEG[6]
port 17 nsew signal output
rlabel metal3 s 44495 20952 44655 21072 6 E2BEG[7]
port 18 nsew signal output
rlabel metal3 s 44495 21224 44655 21344 6 E2BEGb[0]
port 19 nsew signal output
rlabel metal3 s 44495 21496 44655 21616 6 E2BEGb[1]
port 20 nsew signal output
rlabel metal3 s 44495 21768 44655 21888 6 E2BEGb[2]
port 21 nsew signal output
rlabel metal3 s 44495 22040 44655 22160 6 E2BEGb[3]
port 22 nsew signal output
rlabel metal3 s 44495 22312 44655 22432 6 E2BEGb[4]
port 23 nsew signal output
rlabel metal3 s 44495 22584 44655 22704 6 E2BEGb[5]
port 24 nsew signal output
rlabel metal3 s 44495 22856 44655 22976 6 E2BEGb[6]
port 25 nsew signal output
rlabel metal3 s 44495 23128 44655 23248 6 E2BEGb[7]
port 26 nsew signal output
rlabel metal3 s 0 21224 160 21344 6 E2END[0]
port 27 nsew signal input
rlabel metal3 s 0 21496 160 21616 6 E2END[1]
port 28 nsew signal input
rlabel metal3 s 0 21768 160 21888 6 E2END[2]
port 29 nsew signal input
rlabel metal3 s 0 22040 160 22160 6 E2END[3]
port 30 nsew signal input
rlabel metal3 s 0 22312 160 22432 6 E2END[4]
port 31 nsew signal input
rlabel metal3 s 0 22584 160 22704 6 E2END[5]
port 32 nsew signal input
rlabel metal3 s 0 22856 160 22976 6 E2END[6]
port 33 nsew signal input
rlabel metal3 s 0 23128 160 23248 6 E2END[7]
port 34 nsew signal input
rlabel metal3 s 0 19048 160 19168 6 E2MID[0]
port 35 nsew signal input
rlabel metal3 s 0 19320 160 19440 6 E2MID[1]
port 36 nsew signal input
rlabel metal3 s 0 19592 160 19712 6 E2MID[2]
port 37 nsew signal input
rlabel metal3 s 0 19864 160 19984 6 E2MID[3]
port 38 nsew signal input
rlabel metal3 s 0 20136 160 20256 6 E2MID[4]
port 39 nsew signal input
rlabel metal3 s 0 20408 160 20528 6 E2MID[5]
port 40 nsew signal input
rlabel metal3 s 0 20680 160 20800 6 E2MID[6]
port 41 nsew signal input
rlabel metal3 s 0 20952 160 21072 6 E2MID[7]
port 42 nsew signal input
rlabel metal3 s 44495 27752 44655 27872 6 E6BEG[0]
port 43 nsew signal output
rlabel metal3 s 44495 30472 44655 30592 6 E6BEG[10]
port 44 nsew signal output
rlabel metal3 s 44495 30744 44655 30864 6 E6BEG[11]
port 45 nsew signal output
rlabel metal3 s 44495 28024 44655 28144 6 E6BEG[1]
port 46 nsew signal output
rlabel metal3 s 44495 28296 44655 28416 6 E6BEG[2]
port 47 nsew signal output
rlabel metal3 s 44495 28568 44655 28688 6 E6BEG[3]
port 48 nsew signal output
rlabel metal3 s 44495 28840 44655 28960 6 E6BEG[4]
port 49 nsew signal output
rlabel metal3 s 44495 29112 44655 29232 6 E6BEG[5]
port 50 nsew signal output
rlabel metal3 s 44495 29384 44655 29504 6 E6BEG[6]
port 51 nsew signal output
rlabel metal3 s 44495 29656 44655 29776 6 E6BEG[7]
port 52 nsew signal output
rlabel metal3 s 44495 29928 44655 30048 6 E6BEG[8]
port 53 nsew signal output
rlabel metal3 s 44495 30200 44655 30320 6 E6BEG[9]
port 54 nsew signal output
rlabel metal3 s 0 27752 160 27872 6 E6END[0]
port 55 nsew signal input
rlabel metal3 s 0 30472 160 30592 6 E6END[10]
port 56 nsew signal input
rlabel metal3 s 0 30744 160 30864 6 E6END[11]
port 57 nsew signal input
rlabel metal3 s 0 28024 160 28144 6 E6END[1]
port 58 nsew signal input
rlabel metal3 s 0 28296 160 28416 6 E6END[2]
port 59 nsew signal input
rlabel metal3 s 0 28568 160 28688 6 E6END[3]
port 60 nsew signal input
rlabel metal3 s 0 28840 160 28960 6 E6END[4]
port 61 nsew signal input
rlabel metal3 s 0 29112 160 29232 6 E6END[5]
port 62 nsew signal input
rlabel metal3 s 0 29384 160 29504 6 E6END[6]
port 63 nsew signal input
rlabel metal3 s 0 29656 160 29776 6 E6END[7]
port 64 nsew signal input
rlabel metal3 s 0 29928 160 30048 6 E6END[8]
port 65 nsew signal input
rlabel metal3 s 0 30200 160 30320 6 E6END[9]
port 66 nsew signal input
rlabel metal3 s 44495 23400 44655 23520 6 EE4BEG[0]
port 67 nsew signal output
rlabel metal3 s 44495 26120 44655 26240 6 EE4BEG[10]
port 68 nsew signal output
rlabel metal3 s 44495 26392 44655 26512 6 EE4BEG[11]
port 69 nsew signal output
rlabel metal3 s 44495 26664 44655 26784 6 EE4BEG[12]
port 70 nsew signal output
rlabel metal3 s 44495 26936 44655 27056 6 EE4BEG[13]
port 71 nsew signal output
rlabel metal3 s 44495 27208 44655 27328 6 EE4BEG[14]
port 72 nsew signal output
rlabel metal3 s 44495 27480 44655 27600 6 EE4BEG[15]
port 73 nsew signal output
rlabel metal3 s 44495 23672 44655 23792 6 EE4BEG[1]
port 74 nsew signal output
rlabel metal3 s 44495 23944 44655 24064 6 EE4BEG[2]
port 75 nsew signal output
rlabel metal3 s 44495 24216 44655 24336 6 EE4BEG[3]
port 76 nsew signal output
rlabel metal3 s 44495 24488 44655 24608 6 EE4BEG[4]
port 77 nsew signal output
rlabel metal3 s 44495 24760 44655 24880 6 EE4BEG[5]
port 78 nsew signal output
rlabel metal3 s 44495 25032 44655 25152 6 EE4BEG[6]
port 79 nsew signal output
rlabel metal3 s 44495 25304 44655 25424 6 EE4BEG[7]
port 80 nsew signal output
rlabel metal3 s 44495 25576 44655 25696 6 EE4BEG[8]
port 81 nsew signal output
rlabel metal3 s 44495 25848 44655 25968 6 EE4BEG[9]
port 82 nsew signal output
rlabel metal3 s 0 23400 160 23520 6 EE4END[0]
port 83 nsew signal input
rlabel metal3 s 0 26120 160 26240 6 EE4END[10]
port 84 nsew signal input
rlabel metal3 s 0 26392 160 26512 6 EE4END[11]
port 85 nsew signal input
rlabel metal3 s 0 26664 160 26784 6 EE4END[12]
port 86 nsew signal input
rlabel metal3 s 0 26936 160 27056 6 EE4END[13]
port 87 nsew signal input
rlabel metal3 s 0 27208 160 27328 6 EE4END[14]
port 88 nsew signal input
rlabel metal3 s 0 27480 160 27600 6 EE4END[15]
port 89 nsew signal input
rlabel metal3 s 0 23672 160 23792 6 EE4END[1]
port 90 nsew signal input
rlabel metal3 s 0 23944 160 24064 6 EE4END[2]
port 91 nsew signal input
rlabel metal3 s 0 24216 160 24336 6 EE4END[3]
port 92 nsew signal input
rlabel metal3 s 0 24488 160 24608 6 EE4END[4]
port 93 nsew signal input
rlabel metal3 s 0 24760 160 24880 6 EE4END[5]
port 94 nsew signal input
rlabel metal3 s 0 25032 160 25152 6 EE4END[6]
port 95 nsew signal input
rlabel metal3 s 0 25304 160 25424 6 EE4END[7]
port 96 nsew signal input
rlabel metal3 s 0 25576 160 25696 6 EE4END[8]
port 97 nsew signal input
rlabel metal3 s 0 25848 160 25968 6 EE4END[9]
port 98 nsew signal input
rlabel metal3 s 0 31016 160 31136 6 FrameData[0]
port 99 nsew signal input
rlabel metal3 s 0 33736 160 33856 6 FrameData[10]
port 100 nsew signal input
rlabel metal3 s 0 34008 160 34128 6 FrameData[11]
port 101 nsew signal input
rlabel metal3 s 0 34280 160 34400 6 FrameData[12]
port 102 nsew signal input
rlabel metal3 s 0 34552 160 34672 6 FrameData[13]
port 103 nsew signal input
rlabel metal3 s 0 34824 160 34944 6 FrameData[14]
port 104 nsew signal input
rlabel metal3 s 0 35096 160 35216 6 FrameData[15]
port 105 nsew signal input
rlabel metal3 s 0 35368 160 35488 6 FrameData[16]
port 106 nsew signal input
rlabel metal3 s 0 35640 160 35760 6 FrameData[17]
port 107 nsew signal input
rlabel metal3 s 0 35912 160 36032 6 FrameData[18]
port 108 nsew signal input
rlabel metal3 s 0 36184 160 36304 6 FrameData[19]
port 109 nsew signal input
rlabel metal3 s 0 31288 160 31408 6 FrameData[1]
port 110 nsew signal input
rlabel metal3 s 0 36456 160 36576 6 FrameData[20]
port 111 nsew signal input
rlabel metal3 s 0 36728 160 36848 6 FrameData[21]
port 112 nsew signal input
rlabel metal3 s 0 37000 160 37120 6 FrameData[22]
port 113 nsew signal input
rlabel metal3 s 0 37272 160 37392 6 FrameData[23]
port 114 nsew signal input
rlabel metal3 s 0 37544 160 37664 6 FrameData[24]
port 115 nsew signal input
rlabel metal3 s 0 37816 160 37936 6 FrameData[25]
port 116 nsew signal input
rlabel metal3 s 0 38088 160 38208 6 FrameData[26]
port 117 nsew signal input
rlabel metal3 s 0 38360 160 38480 6 FrameData[27]
port 118 nsew signal input
rlabel metal3 s 0 38632 160 38752 6 FrameData[28]
port 119 nsew signal input
rlabel metal3 s 0 38904 160 39024 6 FrameData[29]
port 120 nsew signal input
rlabel metal3 s 0 31560 160 31680 6 FrameData[2]
port 121 nsew signal input
rlabel metal3 s 0 39176 160 39296 6 FrameData[30]
port 122 nsew signal input
rlabel metal3 s 0 39448 160 39568 6 FrameData[31]
port 123 nsew signal input
rlabel metal3 s 0 31832 160 31952 6 FrameData[3]
port 124 nsew signal input
rlabel metal3 s 0 32104 160 32224 6 FrameData[4]
port 125 nsew signal input
rlabel metal3 s 0 32376 160 32496 6 FrameData[5]
port 126 nsew signal input
rlabel metal3 s 0 32648 160 32768 6 FrameData[6]
port 127 nsew signal input
rlabel metal3 s 0 32920 160 33040 6 FrameData[7]
port 128 nsew signal input
rlabel metal3 s 0 33192 160 33312 6 FrameData[8]
port 129 nsew signal input
rlabel metal3 s 0 33464 160 33584 6 FrameData[9]
port 130 nsew signal input
rlabel metal3 s 44495 31016 44655 31136 6 FrameData_O[0]
port 131 nsew signal output
rlabel metal3 s 44495 33736 44655 33856 6 FrameData_O[10]
port 132 nsew signal output
rlabel metal3 s 44495 34008 44655 34128 6 FrameData_O[11]
port 133 nsew signal output
rlabel metal3 s 44495 34280 44655 34400 6 FrameData_O[12]
port 134 nsew signal output
rlabel metal3 s 44495 34552 44655 34672 6 FrameData_O[13]
port 135 nsew signal output
rlabel metal3 s 44495 34824 44655 34944 6 FrameData_O[14]
port 136 nsew signal output
rlabel metal3 s 44495 35096 44655 35216 6 FrameData_O[15]
port 137 nsew signal output
rlabel metal3 s 44495 35368 44655 35488 6 FrameData_O[16]
port 138 nsew signal output
rlabel metal3 s 44495 35640 44655 35760 6 FrameData_O[17]
port 139 nsew signal output
rlabel metal3 s 44495 35912 44655 36032 6 FrameData_O[18]
port 140 nsew signal output
rlabel metal3 s 44495 36184 44655 36304 6 FrameData_O[19]
port 141 nsew signal output
rlabel metal3 s 44495 31288 44655 31408 6 FrameData_O[1]
port 142 nsew signal output
rlabel metal3 s 44495 36456 44655 36576 6 FrameData_O[20]
port 143 nsew signal output
rlabel metal3 s 44495 36728 44655 36848 6 FrameData_O[21]
port 144 nsew signal output
rlabel metal3 s 44495 37000 44655 37120 6 FrameData_O[22]
port 145 nsew signal output
rlabel metal3 s 44495 37272 44655 37392 6 FrameData_O[23]
port 146 nsew signal output
rlabel metal3 s 44495 37544 44655 37664 6 FrameData_O[24]
port 147 nsew signal output
rlabel metal3 s 44495 37816 44655 37936 6 FrameData_O[25]
port 148 nsew signal output
rlabel metal3 s 44495 38088 44655 38208 6 FrameData_O[26]
port 149 nsew signal output
rlabel metal3 s 44495 38360 44655 38480 6 FrameData_O[27]
port 150 nsew signal output
rlabel metal3 s 44495 38632 44655 38752 6 FrameData_O[28]
port 151 nsew signal output
rlabel metal3 s 44495 38904 44655 39024 6 FrameData_O[29]
port 152 nsew signal output
rlabel metal3 s 44495 31560 44655 31680 6 FrameData_O[2]
port 153 nsew signal output
rlabel metal3 s 44495 39176 44655 39296 6 FrameData_O[30]
port 154 nsew signal output
rlabel metal3 s 44495 39448 44655 39568 6 FrameData_O[31]
port 155 nsew signal output
rlabel metal3 s 44495 31832 44655 31952 6 FrameData_O[3]
port 156 nsew signal output
rlabel metal3 s 44495 32104 44655 32224 6 FrameData_O[4]
port 157 nsew signal output
rlabel metal3 s 44495 32376 44655 32496 6 FrameData_O[5]
port 158 nsew signal output
rlabel metal3 s 44495 32648 44655 32768 6 FrameData_O[6]
port 159 nsew signal output
rlabel metal3 s 44495 32920 44655 33040 6 FrameData_O[7]
port 160 nsew signal output
rlabel metal3 s 44495 33192 44655 33312 6 FrameData_O[8]
port 161 nsew signal output
rlabel metal3 s 44495 33464 44655 33584 6 FrameData_O[9]
port 162 nsew signal output
rlabel metal2 s 34242 0 34298 160 6 FrameStrobe[0]
port 163 nsew signal input
rlabel metal2 s 37002 0 37058 160 6 FrameStrobe[10]
port 164 nsew signal input
rlabel metal2 s 37278 0 37334 160 6 FrameStrobe[11]
port 165 nsew signal input
rlabel metal2 s 37554 0 37610 160 6 FrameStrobe[12]
port 166 nsew signal input
rlabel metal2 s 37830 0 37886 160 6 FrameStrobe[13]
port 167 nsew signal input
rlabel metal2 s 38106 0 38162 160 6 FrameStrobe[14]
port 168 nsew signal input
rlabel metal2 s 38382 0 38438 160 6 FrameStrobe[15]
port 169 nsew signal input
rlabel metal2 s 38658 0 38714 160 6 FrameStrobe[16]
port 170 nsew signal input
rlabel metal2 s 38934 0 38990 160 6 FrameStrobe[17]
port 171 nsew signal input
rlabel metal2 s 39210 0 39266 160 6 FrameStrobe[18]
port 172 nsew signal input
rlabel metal2 s 39486 0 39542 160 6 FrameStrobe[19]
port 173 nsew signal input
rlabel metal2 s 34518 0 34574 160 6 FrameStrobe[1]
port 174 nsew signal input
rlabel metal2 s 34794 0 34850 160 6 FrameStrobe[2]
port 175 nsew signal input
rlabel metal2 s 35070 0 35126 160 6 FrameStrobe[3]
port 176 nsew signal input
rlabel metal2 s 35346 0 35402 160 6 FrameStrobe[4]
port 177 nsew signal input
rlabel metal2 s 35622 0 35678 160 6 FrameStrobe[5]
port 178 nsew signal input
rlabel metal2 s 35898 0 35954 160 6 FrameStrobe[6]
port 179 nsew signal input
rlabel metal2 s 36174 0 36230 160 6 FrameStrobe[7]
port 180 nsew signal input
rlabel metal2 s 36450 0 36506 160 6 FrameStrobe[8]
port 181 nsew signal input
rlabel metal2 s 36726 0 36782 160 6 FrameStrobe[9]
port 182 nsew signal input
rlabel metal2 s 34242 44463 34298 44623 6 FrameStrobe_O[0]
port 183 nsew signal output
rlabel metal2 s 37002 44463 37058 44623 6 FrameStrobe_O[10]
port 184 nsew signal output
rlabel metal2 s 37278 44463 37334 44623 6 FrameStrobe_O[11]
port 185 nsew signal output
rlabel metal2 s 37554 44463 37610 44623 6 FrameStrobe_O[12]
port 186 nsew signal output
rlabel metal2 s 37830 44463 37886 44623 6 FrameStrobe_O[13]
port 187 nsew signal output
rlabel metal2 s 38106 44463 38162 44623 6 FrameStrobe_O[14]
port 188 nsew signal output
rlabel metal2 s 38382 44463 38438 44623 6 FrameStrobe_O[15]
port 189 nsew signal output
rlabel metal2 s 38658 44463 38714 44623 6 FrameStrobe_O[16]
port 190 nsew signal output
rlabel metal2 s 38934 44463 38990 44623 6 FrameStrobe_O[17]
port 191 nsew signal output
rlabel metal2 s 39210 44463 39266 44623 6 FrameStrobe_O[18]
port 192 nsew signal output
rlabel metal2 s 39486 44463 39542 44623 6 FrameStrobe_O[19]
port 193 nsew signal output
rlabel metal2 s 34518 44463 34574 44623 6 FrameStrobe_O[1]
port 194 nsew signal output
rlabel metal2 s 34794 44463 34850 44623 6 FrameStrobe_O[2]
port 195 nsew signal output
rlabel metal2 s 35070 44463 35126 44623 6 FrameStrobe_O[3]
port 196 nsew signal output
rlabel metal2 s 35346 44463 35402 44623 6 FrameStrobe_O[4]
port 197 nsew signal output
rlabel metal2 s 35622 44463 35678 44623 6 FrameStrobe_O[5]
port 198 nsew signal output
rlabel metal2 s 35898 44463 35954 44623 6 FrameStrobe_O[6]
port 199 nsew signal output
rlabel metal2 s 36174 44463 36230 44623 6 FrameStrobe_O[7]
port 200 nsew signal output
rlabel metal2 s 36450 44463 36506 44623 6 FrameStrobe_O[8]
port 201 nsew signal output
rlabel metal2 s 36726 44463 36782 44623 6 FrameStrobe_O[9]
port 202 nsew signal output
rlabel metal2 s 4986 44463 5042 44623 6 N1BEG[0]
port 203 nsew signal output
rlabel metal2 s 5262 44463 5318 44623 6 N1BEG[1]
port 204 nsew signal output
rlabel metal2 s 5538 44463 5594 44623 6 N1BEG[2]
port 205 nsew signal output
rlabel metal2 s 5814 44463 5870 44623 6 N1BEG[3]
port 206 nsew signal output
rlabel metal2 s 4986 0 5042 160 6 N1END[0]
port 207 nsew signal input
rlabel metal2 s 5262 0 5318 160 6 N1END[1]
port 208 nsew signal input
rlabel metal2 s 5538 0 5594 160 6 N1END[2]
port 209 nsew signal input
rlabel metal2 s 5814 0 5870 160 6 N1END[3]
port 210 nsew signal input
rlabel metal2 s 6090 44463 6146 44623 6 N2BEG[0]
port 211 nsew signal output
rlabel metal2 s 6366 44463 6422 44623 6 N2BEG[1]
port 212 nsew signal output
rlabel metal2 s 6642 44463 6698 44623 6 N2BEG[2]
port 213 nsew signal output
rlabel metal2 s 6918 44463 6974 44623 6 N2BEG[3]
port 214 nsew signal output
rlabel metal2 s 7194 44463 7250 44623 6 N2BEG[4]
port 215 nsew signal output
rlabel metal2 s 7470 44463 7526 44623 6 N2BEG[5]
port 216 nsew signal output
rlabel metal2 s 7746 44463 7802 44623 6 N2BEG[6]
port 217 nsew signal output
rlabel metal2 s 8022 44463 8078 44623 6 N2BEG[7]
port 218 nsew signal output
rlabel metal2 s 8298 44463 8354 44623 6 N2BEGb[0]
port 219 nsew signal output
rlabel metal2 s 8574 44463 8630 44623 6 N2BEGb[1]
port 220 nsew signal output
rlabel metal2 s 8850 44463 8906 44623 6 N2BEGb[2]
port 221 nsew signal output
rlabel metal2 s 9126 44463 9182 44623 6 N2BEGb[3]
port 222 nsew signal output
rlabel metal2 s 9402 44463 9458 44623 6 N2BEGb[4]
port 223 nsew signal output
rlabel metal2 s 9678 44463 9734 44623 6 N2BEGb[5]
port 224 nsew signal output
rlabel metal2 s 9954 44463 10010 44623 6 N2BEGb[6]
port 225 nsew signal output
rlabel metal2 s 10230 44463 10286 44623 6 N2BEGb[7]
port 226 nsew signal output
rlabel metal2 s 8298 0 8354 160 6 N2END[0]
port 227 nsew signal input
rlabel metal2 s 8574 0 8630 160 6 N2END[1]
port 228 nsew signal input
rlabel metal2 s 8850 0 8906 160 6 N2END[2]
port 229 nsew signal input
rlabel metal2 s 9126 0 9182 160 6 N2END[3]
port 230 nsew signal input
rlabel metal2 s 9402 0 9458 160 6 N2END[4]
port 231 nsew signal input
rlabel metal2 s 9678 0 9734 160 6 N2END[5]
port 232 nsew signal input
rlabel metal2 s 9954 0 10010 160 6 N2END[6]
port 233 nsew signal input
rlabel metal2 s 10230 0 10286 160 6 N2END[7]
port 234 nsew signal input
rlabel metal2 s 6090 0 6146 160 6 N2MID[0]
port 235 nsew signal input
rlabel metal2 s 6366 0 6422 160 6 N2MID[1]
port 236 nsew signal input
rlabel metal2 s 6642 0 6698 160 6 N2MID[2]
port 237 nsew signal input
rlabel metal2 s 6918 0 6974 160 6 N2MID[3]
port 238 nsew signal input
rlabel metal2 s 7194 0 7250 160 6 N2MID[4]
port 239 nsew signal input
rlabel metal2 s 7470 0 7526 160 6 N2MID[5]
port 240 nsew signal input
rlabel metal2 s 7746 0 7802 160 6 N2MID[6]
port 241 nsew signal input
rlabel metal2 s 8022 0 8078 160 6 N2MID[7]
port 242 nsew signal input
rlabel metal2 s 10506 44463 10562 44623 6 N4BEG[0]
port 243 nsew signal output
rlabel metal2 s 13266 44463 13322 44623 6 N4BEG[10]
port 244 nsew signal output
rlabel metal2 s 13542 44463 13598 44623 6 N4BEG[11]
port 245 nsew signal output
rlabel metal2 s 13818 44463 13874 44623 6 N4BEG[12]
port 246 nsew signal output
rlabel metal2 s 14094 44463 14150 44623 6 N4BEG[13]
port 247 nsew signal output
rlabel metal2 s 14370 44463 14426 44623 6 N4BEG[14]
port 248 nsew signal output
rlabel metal2 s 14646 44463 14702 44623 6 N4BEG[15]
port 249 nsew signal output
rlabel metal2 s 10782 44463 10838 44623 6 N4BEG[1]
port 250 nsew signal output
rlabel metal2 s 11058 44463 11114 44623 6 N4BEG[2]
port 251 nsew signal output
rlabel metal2 s 11334 44463 11390 44623 6 N4BEG[3]
port 252 nsew signal output
rlabel metal2 s 11610 44463 11666 44623 6 N4BEG[4]
port 253 nsew signal output
rlabel metal2 s 11886 44463 11942 44623 6 N4BEG[5]
port 254 nsew signal output
rlabel metal2 s 12162 44463 12218 44623 6 N4BEG[6]
port 255 nsew signal output
rlabel metal2 s 12438 44463 12494 44623 6 N4BEG[7]
port 256 nsew signal output
rlabel metal2 s 12714 44463 12770 44623 6 N4BEG[8]
port 257 nsew signal output
rlabel metal2 s 12990 44463 13046 44623 6 N4BEG[9]
port 258 nsew signal output
rlabel metal2 s 10506 0 10562 160 6 N4END[0]
port 259 nsew signal input
rlabel metal2 s 13266 0 13322 160 6 N4END[10]
port 260 nsew signal input
rlabel metal2 s 13542 0 13598 160 6 N4END[11]
port 261 nsew signal input
rlabel metal2 s 13818 0 13874 160 6 N4END[12]
port 262 nsew signal input
rlabel metal2 s 14094 0 14150 160 6 N4END[13]
port 263 nsew signal input
rlabel metal2 s 14370 0 14426 160 6 N4END[14]
port 264 nsew signal input
rlabel metal2 s 14646 0 14702 160 6 N4END[15]
port 265 nsew signal input
rlabel metal2 s 10782 0 10838 160 6 N4END[1]
port 266 nsew signal input
rlabel metal2 s 11058 0 11114 160 6 N4END[2]
port 267 nsew signal input
rlabel metal2 s 11334 0 11390 160 6 N4END[3]
port 268 nsew signal input
rlabel metal2 s 11610 0 11666 160 6 N4END[4]
port 269 nsew signal input
rlabel metal2 s 11886 0 11942 160 6 N4END[5]
port 270 nsew signal input
rlabel metal2 s 12162 0 12218 160 6 N4END[6]
port 271 nsew signal input
rlabel metal2 s 12438 0 12494 160 6 N4END[7]
port 272 nsew signal input
rlabel metal2 s 12714 0 12770 160 6 N4END[8]
port 273 nsew signal input
rlabel metal2 s 12990 0 13046 160 6 N4END[9]
port 274 nsew signal input
rlabel metal2 s 14922 44463 14978 44623 6 NN4BEG[0]
port 275 nsew signal output
rlabel metal2 s 17682 44463 17738 44623 6 NN4BEG[10]
port 276 nsew signal output
rlabel metal2 s 17958 44463 18014 44623 6 NN4BEG[11]
port 277 nsew signal output
rlabel metal2 s 18234 44463 18290 44623 6 NN4BEG[12]
port 278 nsew signal output
rlabel metal2 s 18510 44463 18566 44623 6 NN4BEG[13]
port 279 nsew signal output
rlabel metal2 s 18786 44463 18842 44623 6 NN4BEG[14]
port 280 nsew signal output
rlabel metal2 s 19062 44463 19118 44623 6 NN4BEG[15]
port 281 nsew signal output
rlabel metal2 s 15198 44463 15254 44623 6 NN4BEG[1]
port 282 nsew signal output
rlabel metal2 s 15474 44463 15530 44623 6 NN4BEG[2]
port 283 nsew signal output
rlabel metal2 s 15750 44463 15806 44623 6 NN4BEG[3]
port 284 nsew signal output
rlabel metal2 s 16026 44463 16082 44623 6 NN4BEG[4]
port 285 nsew signal output
rlabel metal2 s 16302 44463 16358 44623 6 NN4BEG[5]
port 286 nsew signal output
rlabel metal2 s 16578 44463 16634 44623 6 NN4BEG[6]
port 287 nsew signal output
rlabel metal2 s 16854 44463 16910 44623 6 NN4BEG[7]
port 288 nsew signal output
rlabel metal2 s 17130 44463 17186 44623 6 NN4BEG[8]
port 289 nsew signal output
rlabel metal2 s 17406 44463 17462 44623 6 NN4BEG[9]
port 290 nsew signal output
rlabel metal2 s 14922 0 14978 160 6 NN4END[0]
port 291 nsew signal input
rlabel metal2 s 17682 0 17738 160 6 NN4END[10]
port 292 nsew signal input
rlabel metal2 s 17958 0 18014 160 6 NN4END[11]
port 293 nsew signal input
rlabel metal2 s 18234 0 18290 160 6 NN4END[12]
port 294 nsew signal input
rlabel metal2 s 18510 0 18566 160 6 NN4END[13]
port 295 nsew signal input
rlabel metal2 s 18786 0 18842 160 6 NN4END[14]
port 296 nsew signal input
rlabel metal2 s 19062 0 19118 160 6 NN4END[15]
port 297 nsew signal input
rlabel metal2 s 15198 0 15254 160 6 NN4END[1]
port 298 nsew signal input
rlabel metal2 s 15474 0 15530 160 6 NN4END[2]
port 299 nsew signal input
rlabel metal2 s 15750 0 15806 160 6 NN4END[3]
port 300 nsew signal input
rlabel metal2 s 16026 0 16082 160 6 NN4END[4]
port 301 nsew signal input
rlabel metal2 s 16302 0 16358 160 6 NN4END[5]
port 302 nsew signal input
rlabel metal2 s 16578 0 16634 160 6 NN4END[6]
port 303 nsew signal input
rlabel metal2 s 16854 0 16910 160 6 NN4END[7]
port 304 nsew signal input
rlabel metal2 s 17130 0 17186 160 6 NN4END[8]
port 305 nsew signal input
rlabel metal2 s 17406 0 17462 160 6 NN4END[9]
port 306 nsew signal input
rlabel metal2 s 19338 0 19394 160 6 S1BEG[0]
port 307 nsew signal output
rlabel metal2 s 19614 0 19670 160 6 S1BEG[1]
port 308 nsew signal output
rlabel metal2 s 19890 0 19946 160 6 S1BEG[2]
port 309 nsew signal output
rlabel metal2 s 20166 0 20222 160 6 S1BEG[3]
port 310 nsew signal output
rlabel metal2 s 19338 44463 19394 44623 6 S1END[0]
port 311 nsew signal input
rlabel metal2 s 19614 44463 19670 44623 6 S1END[1]
port 312 nsew signal input
rlabel metal2 s 19890 44463 19946 44623 6 S1END[2]
port 313 nsew signal input
rlabel metal2 s 20166 44463 20222 44623 6 S1END[3]
port 314 nsew signal input
rlabel metal2 s 22650 0 22706 160 6 S2BEG[0]
port 315 nsew signal output
rlabel metal2 s 22926 0 22982 160 6 S2BEG[1]
port 316 nsew signal output
rlabel metal2 s 23202 0 23258 160 6 S2BEG[2]
port 317 nsew signal output
rlabel metal2 s 23478 0 23534 160 6 S2BEG[3]
port 318 nsew signal output
rlabel metal2 s 23754 0 23810 160 6 S2BEG[4]
port 319 nsew signal output
rlabel metal2 s 24030 0 24086 160 6 S2BEG[5]
port 320 nsew signal output
rlabel metal2 s 24306 0 24362 160 6 S2BEG[6]
port 321 nsew signal output
rlabel metal2 s 24582 0 24638 160 6 S2BEG[7]
port 322 nsew signal output
rlabel metal2 s 20442 0 20498 160 6 S2BEGb[0]
port 323 nsew signal output
rlabel metal2 s 20718 0 20774 160 6 S2BEGb[1]
port 324 nsew signal output
rlabel metal2 s 20994 0 21050 160 6 S2BEGb[2]
port 325 nsew signal output
rlabel metal2 s 21270 0 21326 160 6 S2BEGb[3]
port 326 nsew signal output
rlabel metal2 s 21546 0 21602 160 6 S2BEGb[4]
port 327 nsew signal output
rlabel metal2 s 21822 0 21878 160 6 S2BEGb[5]
port 328 nsew signal output
rlabel metal2 s 22098 0 22154 160 6 S2BEGb[6]
port 329 nsew signal output
rlabel metal2 s 22374 0 22430 160 6 S2BEGb[7]
port 330 nsew signal output
rlabel metal2 s 20442 44463 20498 44623 6 S2END[0]
port 331 nsew signal input
rlabel metal2 s 20718 44463 20774 44623 6 S2END[1]
port 332 nsew signal input
rlabel metal2 s 20994 44463 21050 44623 6 S2END[2]
port 333 nsew signal input
rlabel metal2 s 21270 44463 21326 44623 6 S2END[3]
port 334 nsew signal input
rlabel metal2 s 21546 44463 21602 44623 6 S2END[4]
port 335 nsew signal input
rlabel metal2 s 21822 44463 21878 44623 6 S2END[5]
port 336 nsew signal input
rlabel metal2 s 22098 44463 22154 44623 6 S2END[6]
port 337 nsew signal input
rlabel metal2 s 22374 44463 22430 44623 6 S2END[7]
port 338 nsew signal input
rlabel metal2 s 22650 44463 22706 44623 6 S2MID[0]
port 339 nsew signal input
rlabel metal2 s 22926 44463 22982 44623 6 S2MID[1]
port 340 nsew signal input
rlabel metal2 s 23202 44463 23258 44623 6 S2MID[2]
port 341 nsew signal input
rlabel metal2 s 23478 44463 23534 44623 6 S2MID[3]
port 342 nsew signal input
rlabel metal2 s 23754 44463 23810 44623 6 S2MID[4]
port 343 nsew signal input
rlabel metal2 s 24030 44463 24086 44623 6 S2MID[5]
port 344 nsew signal input
rlabel metal2 s 24306 44463 24362 44623 6 S2MID[6]
port 345 nsew signal input
rlabel metal2 s 24582 44463 24638 44623 6 S2MID[7]
port 346 nsew signal input
rlabel metal2 s 24858 0 24914 160 6 S4BEG[0]
port 347 nsew signal output
rlabel metal2 s 27618 0 27674 160 6 S4BEG[10]
port 348 nsew signal output
rlabel metal2 s 27894 0 27950 160 6 S4BEG[11]
port 349 nsew signal output
rlabel metal2 s 28170 0 28226 160 6 S4BEG[12]
port 350 nsew signal output
rlabel metal2 s 28446 0 28502 160 6 S4BEG[13]
port 351 nsew signal output
rlabel metal2 s 28722 0 28778 160 6 S4BEG[14]
port 352 nsew signal output
rlabel metal2 s 28998 0 29054 160 6 S4BEG[15]
port 353 nsew signal output
rlabel metal2 s 25134 0 25190 160 6 S4BEG[1]
port 354 nsew signal output
rlabel metal2 s 25410 0 25466 160 6 S4BEG[2]
port 355 nsew signal output
rlabel metal2 s 25686 0 25742 160 6 S4BEG[3]
port 356 nsew signal output
rlabel metal2 s 25962 0 26018 160 6 S4BEG[4]
port 357 nsew signal output
rlabel metal2 s 26238 0 26294 160 6 S4BEG[5]
port 358 nsew signal output
rlabel metal2 s 26514 0 26570 160 6 S4BEG[6]
port 359 nsew signal output
rlabel metal2 s 26790 0 26846 160 6 S4BEG[7]
port 360 nsew signal output
rlabel metal2 s 27066 0 27122 160 6 S4BEG[8]
port 361 nsew signal output
rlabel metal2 s 27342 0 27398 160 6 S4BEG[9]
port 362 nsew signal output
rlabel metal2 s 24858 44463 24914 44623 6 S4END[0]
port 363 nsew signal input
rlabel metal2 s 27618 44463 27674 44623 6 S4END[10]
port 364 nsew signal input
rlabel metal2 s 27894 44463 27950 44623 6 S4END[11]
port 365 nsew signal input
rlabel metal2 s 28170 44463 28226 44623 6 S4END[12]
port 366 nsew signal input
rlabel metal2 s 28446 44463 28502 44623 6 S4END[13]
port 367 nsew signal input
rlabel metal2 s 28722 44463 28778 44623 6 S4END[14]
port 368 nsew signal input
rlabel metal2 s 28998 44463 29054 44623 6 S4END[15]
port 369 nsew signal input
rlabel metal2 s 25134 44463 25190 44623 6 S4END[1]
port 370 nsew signal input
rlabel metal2 s 25410 44463 25466 44623 6 S4END[2]
port 371 nsew signal input
rlabel metal2 s 25686 44463 25742 44623 6 S4END[3]
port 372 nsew signal input
rlabel metal2 s 25962 44463 26018 44623 6 S4END[4]
port 373 nsew signal input
rlabel metal2 s 26238 44463 26294 44623 6 S4END[5]
port 374 nsew signal input
rlabel metal2 s 26514 44463 26570 44623 6 S4END[6]
port 375 nsew signal input
rlabel metal2 s 26790 44463 26846 44623 6 S4END[7]
port 376 nsew signal input
rlabel metal2 s 27066 44463 27122 44623 6 S4END[8]
port 377 nsew signal input
rlabel metal2 s 27342 44463 27398 44623 6 S4END[9]
port 378 nsew signal input
rlabel metal2 s 29274 0 29330 160 6 SS4BEG[0]
port 379 nsew signal output
rlabel metal2 s 32034 0 32090 160 6 SS4BEG[10]
port 380 nsew signal output
rlabel metal2 s 32310 0 32366 160 6 SS4BEG[11]
port 381 nsew signal output
rlabel metal2 s 32586 0 32642 160 6 SS4BEG[12]
port 382 nsew signal output
rlabel metal2 s 32862 0 32918 160 6 SS4BEG[13]
port 383 nsew signal output
rlabel metal2 s 33138 0 33194 160 6 SS4BEG[14]
port 384 nsew signal output
rlabel metal2 s 33414 0 33470 160 6 SS4BEG[15]
port 385 nsew signal output
rlabel metal2 s 29550 0 29606 160 6 SS4BEG[1]
port 386 nsew signal output
rlabel metal2 s 29826 0 29882 160 6 SS4BEG[2]
port 387 nsew signal output
rlabel metal2 s 30102 0 30158 160 6 SS4BEG[3]
port 388 nsew signal output
rlabel metal2 s 30378 0 30434 160 6 SS4BEG[4]
port 389 nsew signal output
rlabel metal2 s 30654 0 30710 160 6 SS4BEG[5]
port 390 nsew signal output
rlabel metal2 s 30930 0 30986 160 6 SS4BEG[6]
port 391 nsew signal output
rlabel metal2 s 31206 0 31262 160 6 SS4BEG[7]
port 392 nsew signal output
rlabel metal2 s 31482 0 31538 160 6 SS4BEG[8]
port 393 nsew signal output
rlabel metal2 s 31758 0 31814 160 6 SS4BEG[9]
port 394 nsew signal output
rlabel metal2 s 29274 44463 29330 44623 6 SS4END[0]
port 395 nsew signal input
rlabel metal2 s 32034 44463 32090 44623 6 SS4END[10]
port 396 nsew signal input
rlabel metal2 s 32310 44463 32366 44623 6 SS4END[11]
port 397 nsew signal input
rlabel metal2 s 32586 44463 32642 44623 6 SS4END[12]
port 398 nsew signal input
rlabel metal2 s 32862 44463 32918 44623 6 SS4END[13]
port 399 nsew signal input
rlabel metal2 s 33138 44463 33194 44623 6 SS4END[14]
port 400 nsew signal input
rlabel metal2 s 33414 44463 33470 44623 6 SS4END[15]
port 401 nsew signal input
rlabel metal2 s 29550 44463 29606 44623 6 SS4END[1]
port 402 nsew signal input
rlabel metal2 s 29826 44463 29882 44623 6 SS4END[2]
port 403 nsew signal input
rlabel metal2 s 30102 44463 30158 44623 6 SS4END[3]
port 404 nsew signal input
rlabel metal2 s 30378 44463 30434 44623 6 SS4END[4]
port 405 nsew signal input
rlabel metal2 s 30654 44463 30710 44623 6 SS4END[5]
port 406 nsew signal input
rlabel metal2 s 30930 44463 30986 44623 6 SS4END[6]
port 407 nsew signal input
rlabel metal2 s 31206 44463 31262 44623 6 SS4END[7]
port 408 nsew signal input
rlabel metal2 s 31482 44463 31538 44623 6 SS4END[8]
port 409 nsew signal input
rlabel metal2 s 31758 44463 31814 44623 6 SS4END[9]
port 410 nsew signal input
rlabel metal2 s 33690 0 33746 160 6 UserCLK
port 411 nsew signal input
rlabel metal2 s 33690 44463 33746 44623 6 UserCLKo
port 412 nsew signal output
rlabel metal4 s 19568 1040 19888 43568 6 VGND
port 413 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 43568 6 VPWR
port 414 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 43568 6 VPWR
port 414 nsew power bidirectional
rlabel metal3 s 0 4904 160 5024 6 W1BEG[0]
port 415 nsew signal output
rlabel metal3 s 0 5176 160 5296 6 W1BEG[1]
port 416 nsew signal output
rlabel metal3 s 0 5448 160 5568 6 W1BEG[2]
port 417 nsew signal output
rlabel metal3 s 0 5720 160 5840 6 W1BEG[3]
port 418 nsew signal output
rlabel metal3 s 44495 4904 44655 5024 6 W1END[0]
port 419 nsew signal input
rlabel metal3 s 44495 5176 44655 5296 6 W1END[1]
port 420 nsew signal input
rlabel metal3 s 44495 5448 44655 5568 6 W1END[2]
port 421 nsew signal input
rlabel metal3 s 44495 5720 44655 5840 6 W1END[3]
port 422 nsew signal input
rlabel metal3 s 0 5992 160 6112 6 W2BEG[0]
port 423 nsew signal output
rlabel metal3 s 0 6264 160 6384 6 W2BEG[1]
port 424 nsew signal output
rlabel metal3 s 0 6536 160 6656 6 W2BEG[2]
port 425 nsew signal output
rlabel metal3 s 0 6808 160 6928 6 W2BEG[3]
port 426 nsew signal output
rlabel metal3 s 0 7080 160 7200 6 W2BEG[4]
port 427 nsew signal output
rlabel metal3 s 0 7352 160 7472 6 W2BEG[5]
port 428 nsew signal output
rlabel metal3 s 0 7624 160 7744 6 W2BEG[6]
port 429 nsew signal output
rlabel metal3 s 0 7896 160 8016 6 W2BEG[7]
port 430 nsew signal output
rlabel metal3 s 0 8168 160 8288 6 W2BEGb[0]
port 431 nsew signal output
rlabel metal3 s 0 8440 160 8560 6 W2BEGb[1]
port 432 nsew signal output
rlabel metal3 s 0 8712 160 8832 6 W2BEGb[2]
port 433 nsew signal output
rlabel metal3 s 0 8984 160 9104 6 W2BEGb[3]
port 434 nsew signal output
rlabel metal3 s 0 9256 160 9376 6 W2BEGb[4]
port 435 nsew signal output
rlabel metal3 s 0 9528 160 9648 6 W2BEGb[5]
port 436 nsew signal output
rlabel metal3 s 0 9800 160 9920 6 W2BEGb[6]
port 437 nsew signal output
rlabel metal3 s 0 10072 160 10192 6 W2BEGb[7]
port 438 nsew signal output
rlabel metal3 s 44495 8168 44655 8288 6 W2END[0]
port 439 nsew signal input
rlabel metal3 s 44495 8440 44655 8560 6 W2END[1]
port 440 nsew signal input
rlabel metal3 s 44495 8712 44655 8832 6 W2END[2]
port 441 nsew signal input
rlabel metal3 s 44495 8984 44655 9104 6 W2END[3]
port 442 nsew signal input
rlabel metal3 s 44495 9256 44655 9376 6 W2END[4]
port 443 nsew signal input
rlabel metal3 s 44495 9528 44655 9648 6 W2END[5]
port 444 nsew signal input
rlabel metal3 s 44495 9800 44655 9920 6 W2END[6]
port 445 nsew signal input
rlabel metal3 s 44495 10072 44655 10192 6 W2END[7]
port 446 nsew signal input
rlabel metal3 s 44495 5992 44655 6112 6 W2MID[0]
port 447 nsew signal input
rlabel metal3 s 44495 6264 44655 6384 6 W2MID[1]
port 448 nsew signal input
rlabel metal3 s 44495 6536 44655 6656 6 W2MID[2]
port 449 nsew signal input
rlabel metal3 s 44495 6808 44655 6928 6 W2MID[3]
port 450 nsew signal input
rlabel metal3 s 44495 7080 44655 7200 6 W2MID[4]
port 451 nsew signal input
rlabel metal3 s 44495 7352 44655 7472 6 W2MID[5]
port 452 nsew signal input
rlabel metal3 s 44495 7624 44655 7744 6 W2MID[6]
port 453 nsew signal input
rlabel metal3 s 44495 7896 44655 8016 6 W2MID[7]
port 454 nsew signal input
rlabel metal3 s 0 14696 160 14816 6 W6BEG[0]
port 455 nsew signal output
rlabel metal3 s 0 17416 160 17536 6 W6BEG[10]
port 456 nsew signal output
rlabel metal3 s 0 17688 160 17808 6 W6BEG[11]
port 457 nsew signal output
rlabel metal3 s 0 14968 160 15088 6 W6BEG[1]
port 458 nsew signal output
rlabel metal3 s 0 15240 160 15360 6 W6BEG[2]
port 459 nsew signal output
rlabel metal3 s 0 15512 160 15632 6 W6BEG[3]
port 460 nsew signal output
rlabel metal3 s 0 15784 160 15904 6 W6BEG[4]
port 461 nsew signal output
rlabel metal3 s 0 16056 160 16176 6 W6BEG[5]
port 462 nsew signal output
rlabel metal3 s 0 16328 160 16448 6 W6BEG[6]
port 463 nsew signal output
rlabel metal3 s 0 16600 160 16720 6 W6BEG[7]
port 464 nsew signal output
rlabel metal3 s 0 16872 160 16992 6 W6BEG[8]
port 465 nsew signal output
rlabel metal3 s 0 17144 160 17264 6 W6BEG[9]
port 466 nsew signal output
rlabel metal3 s 44495 14696 44655 14816 6 W6END[0]
port 467 nsew signal input
rlabel metal3 s 44495 17416 44655 17536 6 W6END[10]
port 468 nsew signal input
rlabel metal3 s 44495 17688 44655 17808 6 W6END[11]
port 469 nsew signal input
rlabel metal3 s 44495 14968 44655 15088 6 W6END[1]
port 470 nsew signal input
rlabel metal3 s 44495 15240 44655 15360 6 W6END[2]
port 471 nsew signal input
rlabel metal3 s 44495 15512 44655 15632 6 W6END[3]
port 472 nsew signal input
rlabel metal3 s 44495 15784 44655 15904 6 W6END[4]
port 473 nsew signal input
rlabel metal3 s 44495 16056 44655 16176 6 W6END[5]
port 474 nsew signal input
rlabel metal3 s 44495 16328 44655 16448 6 W6END[6]
port 475 nsew signal input
rlabel metal3 s 44495 16600 44655 16720 6 W6END[7]
port 476 nsew signal input
rlabel metal3 s 44495 16872 44655 16992 6 W6END[8]
port 477 nsew signal input
rlabel metal3 s 44495 17144 44655 17264 6 W6END[9]
port 478 nsew signal input
rlabel metal3 s 0 10344 160 10464 6 WW4BEG[0]
port 479 nsew signal output
rlabel metal3 s 0 13064 160 13184 6 WW4BEG[10]
port 480 nsew signal output
rlabel metal3 s 0 13336 160 13456 6 WW4BEG[11]
port 481 nsew signal output
rlabel metal3 s 0 13608 160 13728 6 WW4BEG[12]
port 482 nsew signal output
rlabel metal3 s 0 13880 160 14000 6 WW4BEG[13]
port 483 nsew signal output
rlabel metal3 s 0 14152 160 14272 6 WW4BEG[14]
port 484 nsew signal output
rlabel metal3 s 0 14424 160 14544 6 WW4BEG[15]
port 485 nsew signal output
rlabel metal3 s 0 10616 160 10736 6 WW4BEG[1]
port 486 nsew signal output
rlabel metal3 s 0 10888 160 11008 6 WW4BEG[2]
port 487 nsew signal output
rlabel metal3 s 0 11160 160 11280 6 WW4BEG[3]
port 488 nsew signal output
rlabel metal3 s 0 11432 160 11552 6 WW4BEG[4]
port 489 nsew signal output
rlabel metal3 s 0 11704 160 11824 6 WW4BEG[5]
port 490 nsew signal output
rlabel metal3 s 0 11976 160 12096 6 WW4BEG[6]
port 491 nsew signal output
rlabel metal3 s 0 12248 160 12368 6 WW4BEG[7]
port 492 nsew signal output
rlabel metal3 s 0 12520 160 12640 6 WW4BEG[8]
port 493 nsew signal output
rlabel metal3 s 0 12792 160 12912 6 WW4BEG[9]
port 494 nsew signal output
rlabel metal3 s 44495 10344 44655 10464 6 WW4END[0]
port 495 nsew signal input
rlabel metal3 s 44495 13064 44655 13184 6 WW4END[10]
port 496 nsew signal input
rlabel metal3 s 44495 13336 44655 13456 6 WW4END[11]
port 497 nsew signal input
rlabel metal3 s 44495 13608 44655 13728 6 WW4END[12]
port 498 nsew signal input
rlabel metal3 s 44495 13880 44655 14000 6 WW4END[13]
port 499 nsew signal input
rlabel metal3 s 44495 14152 44655 14272 6 WW4END[14]
port 500 nsew signal input
rlabel metal3 s 44495 14424 44655 14544 6 WW4END[15]
port 501 nsew signal input
rlabel metal3 s 44495 10616 44655 10736 6 WW4END[1]
port 502 nsew signal input
rlabel metal3 s 44495 10888 44655 11008 6 WW4END[2]
port 503 nsew signal input
rlabel metal3 s 44495 11160 44655 11280 6 WW4END[3]
port 504 nsew signal input
rlabel metal3 s 44495 11432 44655 11552 6 WW4END[4]
port 505 nsew signal input
rlabel metal3 s 44495 11704 44655 11824 6 WW4END[5]
port 506 nsew signal input
rlabel metal3 s 44495 11976 44655 12096 6 WW4END[6]
port 507 nsew signal input
rlabel metal3 s 44495 12248 44655 12368 6 WW4END[7]
port 508 nsew signal input
rlabel metal3 s 44495 12520 44655 12640 6 WW4END[8]
port 509 nsew signal input
rlabel metal3 s 44495 12792 44655 12912 6 WW4END[9]
port 510 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 44655 44623
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7918788
string GDS_FILE /home/asma/Desktop/FPGA_IGNITE_2024/openlane/LUT_redo/runs/24_11_24_22_23/results/signoff/LUT4AB.magic.gds
string GDS_START 224838
<< end >>

