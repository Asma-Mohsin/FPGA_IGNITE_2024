module eFPGA_top #(
    /* verilator lint_off UNUSEDSIGNAL */
    /* verilator lint_off UNUSEDPARAM*/

    parameter include_eFPGA = 1,
    parameter NumberOfRows = 6,
    parameter NumberOfCols = 10,
    parameter FrameBitsPerRow = 32,
    parameter MaxFramesPerCol = 20,
    parameter desync_flag = 20,
    parameter FrameSelectWidth = 5,
    parameter RowSelectWidth = 5
    /* verilator lint_on UNUSEDPARAM*/
) (
`ifdef USE_POWER_PINS
    input wire vccd1,
    input wire vssd1,
`endif
    //External IO port
    output [23:0] A_config_C,
    output [23:0] B_config_C,
    output [23:0] Config_accessC,
    output [11:0] I_top,
    input [11:0] O_top,
    output [11:0] T_top,
    input [159:0] UIO_BOT_UIN,
    output [159:0] UIO_BOT_UOUT,
    input [159:0] UIO_TOP_UIN,
    output [159:0] UIO_TOP_UOUT,
    //Config related ports
    input CLK,
    input resetn,
    input SelfWriteStrobe,
    input [31:0] SelfWriteData,
    input Rx,
    output ComActive,
    output ReceiveLED,
    input s_clk,
    input s_data
);
    //BlockRAM ports

    wire [96-1:0] RAM2FAB_D_I;
    wire [96-1:0] FAB2RAM_D_O;
    wire [48-1:0] FAB2RAM_A_O;
    wire [24-1:0] FAB2RAM_C_O;

    //Signal declarations
    wire [(NumberOfRows*FrameBitsPerRow)-1:0] FrameRegister;
    wire [(MaxFramesPerCol*NumberOfCols)-1:0] FrameSelect;
    wire [(FrameBitsPerRow*(NumberOfRows+2))-1:0] FrameData;
    wire [FrameBitsPerRow-1:0] FrameAddressRegister;
    wire LongFrameStrobe;
    wire [31:0] LocalWriteData;
    wire LocalWriteStrobe;
    wire [RowSelectWidth-1:0] RowSelect;
    wire resten;
`ifndef EMULATION

    eFPGA_Config #(
        .RowSelectWidth(RowSelectWidth),
        .NumberOfRows(NumberOfRows),
        .desync_flag(desync_flag),
        .FrameBitsPerRow(FrameBitsPerRow)
    ) eFPGA_Config_inst (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .CLK(CLK),
        .resetn(resetn),
        .Rx(Rx),
        .ComActive(ComActive),
        .ReceiveLED(ReceiveLED),
        .s_clk(s_clk),
        .s_data(s_data),
        .SelfWriteData(SelfWriteData),
        .SelfWriteStrobe(SelfWriteStrobe),
        .ConfigWriteData(LocalWriteData),
        .ConfigWriteStrobe(LocalWriteStrobe),
        .FrameAddressRegister(FrameAddressRegister),
        .LongFrameStrobe(LongFrameStrobe),
        .RowSelect(RowSelect)
    );


    Frame_Data_Reg #(
        .FrameBitsPerRow(FrameBitsPerRow),
        .RowSelectWidth(RowSelectWidth),
        .Row(1)
    ) inst_Frame_Data_Reg_0 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameData_I(LocalWriteData),
        .FrameData_O(FrameRegister[0*FrameBitsPerRow+FrameBitsPerRow-1:0*FrameBitsPerRow]),
        .RowSelect(RowSelect),
        .CLK(CLK)
    );

    Frame_Data_Reg #(
        .FrameBitsPerRow(FrameBitsPerRow),
        .RowSelectWidth(RowSelectWidth),
        .Row(2)
    ) inst_Frame_Data_Reg_1 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameData_I(LocalWriteData),
        .FrameData_O(FrameRegister[1*FrameBitsPerRow+FrameBitsPerRow-1:1*FrameBitsPerRow]),
        .RowSelect(RowSelect),
        .CLK(CLK)
    );

    Frame_Data_Reg #(
        .FrameBitsPerRow(FrameBitsPerRow),
        .RowSelectWidth(RowSelectWidth),
        .Row(3)
    ) inst_Frame_Data_Reg_2 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameData_I(LocalWriteData),
        .FrameData_O(FrameRegister[2*FrameBitsPerRow+FrameBitsPerRow-1:2*FrameBitsPerRow]),
        .RowSelect(RowSelect),
        .CLK(CLK)
    );

    Frame_Data_Reg #(
        .FrameBitsPerRow(FrameBitsPerRow),
        .RowSelectWidth(RowSelectWidth),
        .Row(4)
    ) inst_Frame_Data_Reg_3 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameData_I(LocalWriteData),
        .FrameData_O(FrameRegister[3*FrameBitsPerRow+FrameBitsPerRow-1:3*FrameBitsPerRow]),
        .RowSelect(RowSelect),
        .CLK(CLK)
    );

    Frame_Data_Reg #(
        .FrameBitsPerRow(FrameBitsPerRow),
        .RowSelectWidth(RowSelectWidth),
        .Row(5)
    ) inst_Frame_Data_Reg_4 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameData_I(LocalWriteData),
        .FrameData_O(FrameRegister[4*FrameBitsPerRow+FrameBitsPerRow-1:4*FrameBitsPerRow]),
        .RowSelect(RowSelect),
        .CLK(CLK)
    );

    Frame_Data_Reg #(
        .FrameBitsPerRow(FrameBitsPerRow),
        .RowSelectWidth(RowSelectWidth),
        .Row(6)
    ) inst_Frame_Data_Reg_5 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameData_I(LocalWriteData),
        .FrameData_O(FrameRegister[5*FrameBitsPerRow+FrameBitsPerRow-1:5*FrameBitsPerRow]),
        .RowSelect(RowSelect),
        .CLK(CLK)
    );


    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(0)
    ) inst_Frame_Select_0 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[0*MaxFramesPerCol+MaxFramesPerCol-1:0*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(1)
    ) inst_Frame_Select_1 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[1*MaxFramesPerCol+MaxFramesPerCol-1:1*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(2)
    ) inst_Frame_Select_2 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[2*MaxFramesPerCol+MaxFramesPerCol-1:2*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(3)
    ) inst_Frame_Select_3 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[3*MaxFramesPerCol+MaxFramesPerCol-1:3*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(4)
    ) inst_Frame_Select_4 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[4*MaxFramesPerCol+MaxFramesPerCol-1:4*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(5)
    ) inst_Frame_Select_5 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[5*MaxFramesPerCol+MaxFramesPerCol-1:5*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(6)
    ) inst_Frame_Select_6 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[6*MaxFramesPerCol+MaxFramesPerCol-1:6*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(7)
    ) inst_Frame_Select_7 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[7*MaxFramesPerCol+MaxFramesPerCol-1:7*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(8)
    ) inst_Frame_Select_8 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[8*MaxFramesPerCol+MaxFramesPerCol-1:8*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );

    Frame_Select #(
        .MaxFramesPerCol(MaxFramesPerCol),
        .FrameSelectWidth(FrameSelectWidth),
        .Col(9)
    ) inst_Frame_Select_9 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .FrameStrobe_I(FrameAddressRegister[MaxFramesPerCol-1:0]),
        .FrameStrobe_O(FrameSelect[9*MaxFramesPerCol+MaxFramesPerCol-1:9*MaxFramesPerCol]),
        .FrameSelect(FrameAddressRegister[FrameBitsPerRow-1:FrameBitsPerRow-FrameSelectWidth]),
        .FrameStrobe(LongFrameStrobe)
    );


`endif
    eFPGA eFPGA_inst (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .Tile_X0Y6_A_config_C_bit0(A_config_C[0]),
        .Tile_X0Y6_A_config_C_bit1(A_config_C[1]),
        .Tile_X0Y6_A_config_C_bit2(A_config_C[2]),
        .Tile_X0Y6_A_config_C_bit3(A_config_C[3]),
        .Tile_X0Y5_A_config_C_bit0(A_config_C[4]),
        .Tile_X0Y5_A_config_C_bit1(A_config_C[5]),
        .Tile_X0Y5_A_config_C_bit2(A_config_C[6]),
        .Tile_X0Y5_A_config_C_bit3(A_config_C[7]),
        .Tile_X0Y4_A_config_C_bit0(A_config_C[8]),
        .Tile_X0Y4_A_config_C_bit1(A_config_C[9]),
        .Tile_X0Y4_A_config_C_bit2(A_config_C[10]),
        .Tile_X0Y4_A_config_C_bit3(A_config_C[11]),
        .Tile_X0Y3_A_config_C_bit0(A_config_C[12]),
        .Tile_X0Y3_A_config_C_bit1(A_config_C[13]),
        .Tile_X0Y3_A_config_C_bit2(A_config_C[14]),
        .Tile_X0Y3_A_config_C_bit3(A_config_C[15]),
        .Tile_X0Y2_A_config_C_bit0(A_config_C[16]),
        .Tile_X0Y2_A_config_C_bit1(A_config_C[17]),
        .Tile_X0Y2_A_config_C_bit2(A_config_C[18]),
        .Tile_X0Y2_A_config_C_bit3(A_config_C[19]),
        .Tile_X0Y1_A_config_C_bit0(A_config_C[20]),
        .Tile_X0Y1_A_config_C_bit1(A_config_C[21]),
        .Tile_X0Y1_A_config_C_bit2(A_config_C[22]),
        .Tile_X0Y1_A_config_C_bit3(A_config_C[23]),
        .Tile_X0Y6_B_config_C_bit0(B_config_C[0]),
        .Tile_X0Y6_B_config_C_bit1(B_config_C[1]),
        .Tile_X0Y6_B_config_C_bit2(B_config_C[2]),
        .Tile_X0Y6_B_config_C_bit3(B_config_C[3]),
        .Tile_X0Y5_B_config_C_bit0(B_config_C[4]),
        .Tile_X0Y5_B_config_C_bit1(B_config_C[5]),
        .Tile_X0Y5_B_config_C_bit2(B_config_C[6]),
        .Tile_X0Y5_B_config_C_bit3(B_config_C[7]),
        .Tile_X0Y4_B_config_C_bit0(B_config_C[8]),
        .Tile_X0Y4_B_config_C_bit1(B_config_C[9]),
        .Tile_X0Y4_B_config_C_bit2(B_config_C[10]),
        .Tile_X0Y4_B_config_C_bit3(B_config_C[11]),
        .Tile_X0Y3_B_config_C_bit0(B_config_C[12]),
        .Tile_X0Y3_B_config_C_bit1(B_config_C[13]),
        .Tile_X0Y3_B_config_C_bit2(B_config_C[14]),
        .Tile_X0Y3_B_config_C_bit3(B_config_C[15]),
        .Tile_X0Y2_B_config_C_bit0(B_config_C[16]),
        .Tile_X0Y2_B_config_C_bit1(B_config_C[17]),
        .Tile_X0Y2_B_config_C_bit2(B_config_C[18]),
        .Tile_X0Y2_B_config_C_bit3(B_config_C[19]),
        .Tile_X0Y1_B_config_C_bit0(B_config_C[20]),
        .Tile_X0Y1_B_config_C_bit1(B_config_C[21]),
        .Tile_X0Y1_B_config_C_bit2(B_config_C[22]),
        .Tile_X0Y1_B_config_C_bit3(B_config_C[23]),
        .Tile_X9Y6_Config_accessC_bit0(Config_accessC[0]),
        .Tile_X9Y6_Config_accessC_bit1(Config_accessC[1]),
        .Tile_X9Y6_Config_accessC_bit2(Config_accessC[2]),
        .Tile_X9Y6_Config_accessC_bit3(Config_accessC[3]),
        .Tile_X9Y5_Config_accessC_bit0(Config_accessC[4]),
        .Tile_X9Y5_Config_accessC_bit1(Config_accessC[5]),
        .Tile_X9Y5_Config_accessC_bit2(Config_accessC[6]),
        .Tile_X9Y5_Config_accessC_bit3(Config_accessC[7]),
        .Tile_X9Y4_Config_accessC_bit0(Config_accessC[8]),
        .Tile_X9Y4_Config_accessC_bit1(Config_accessC[9]),
        .Tile_X9Y4_Config_accessC_bit2(Config_accessC[10]),
        .Tile_X9Y4_Config_accessC_bit3(Config_accessC[11]),
        .Tile_X9Y3_Config_accessC_bit0(Config_accessC[12]),
        .Tile_X9Y3_Config_accessC_bit1(Config_accessC[13]),
        .Tile_X9Y3_Config_accessC_bit2(Config_accessC[14]),
        .Tile_X9Y3_Config_accessC_bit3(Config_accessC[15]),
        .Tile_X9Y2_Config_accessC_bit0(Config_accessC[16]),
        .Tile_X9Y2_Config_accessC_bit1(Config_accessC[17]),
        .Tile_X9Y2_Config_accessC_bit2(Config_accessC[18]),
        .Tile_X9Y2_Config_accessC_bit3(Config_accessC[19]),
        .Tile_X9Y1_Config_accessC_bit0(Config_accessC[20]),
        .Tile_X9Y1_Config_accessC_bit1(Config_accessC[21]),
        .Tile_X9Y1_Config_accessC_bit2(Config_accessC[22]),
        .Tile_X9Y1_Config_accessC_bit3(Config_accessC[23]),
        .Tile_X9Y6_FAB2RAM_A0_O0(FAB2RAM_A_O[0]),
        .Tile_X9Y6_FAB2RAM_A0_O1(FAB2RAM_A_O[1]),
        .Tile_X9Y6_FAB2RAM_A0_O2(FAB2RAM_A_O[2]),
        .Tile_X9Y6_FAB2RAM_A0_O3(FAB2RAM_A_O[3]),
        .Tile_X9Y6_FAB2RAM_A1_O0(FAB2RAM_A_O[4]),
        .Tile_X9Y6_FAB2RAM_A1_O1(FAB2RAM_A_O[5]),
        .Tile_X9Y6_FAB2RAM_A1_O2(FAB2RAM_A_O[6]),
        .Tile_X9Y6_FAB2RAM_A1_O3(FAB2RAM_A_O[7]),
        .Tile_X9Y5_FAB2RAM_A0_O0(FAB2RAM_A_O[8]),
        .Tile_X9Y5_FAB2RAM_A0_O1(FAB2RAM_A_O[9]),
        .Tile_X9Y5_FAB2RAM_A0_O2(FAB2RAM_A_O[10]),
        .Tile_X9Y5_FAB2RAM_A0_O3(FAB2RAM_A_O[11]),
        .Tile_X9Y5_FAB2RAM_A1_O0(FAB2RAM_A_O[12]),
        .Tile_X9Y5_FAB2RAM_A1_O1(FAB2RAM_A_O[13]),
        .Tile_X9Y5_FAB2RAM_A1_O2(FAB2RAM_A_O[14]),
        .Tile_X9Y5_FAB2RAM_A1_O3(FAB2RAM_A_O[15]),
        .Tile_X9Y4_FAB2RAM_A0_O0(FAB2RAM_A_O[16]),
        .Tile_X9Y4_FAB2RAM_A0_O1(FAB2RAM_A_O[17]),
        .Tile_X9Y4_FAB2RAM_A0_O2(FAB2RAM_A_O[18]),
        .Tile_X9Y4_FAB2RAM_A0_O3(FAB2RAM_A_O[19]),
        .Tile_X9Y4_FAB2RAM_A1_O0(FAB2RAM_A_O[20]),
        .Tile_X9Y4_FAB2RAM_A1_O1(FAB2RAM_A_O[21]),
        .Tile_X9Y4_FAB2RAM_A1_O2(FAB2RAM_A_O[22]),
        .Tile_X9Y4_FAB2RAM_A1_O3(FAB2RAM_A_O[23]),
        .Tile_X9Y3_FAB2RAM_A0_O0(FAB2RAM_A_O[24]),
        .Tile_X9Y3_FAB2RAM_A0_O1(FAB2RAM_A_O[25]),
        .Tile_X9Y3_FAB2RAM_A0_O2(FAB2RAM_A_O[26]),
        .Tile_X9Y3_FAB2RAM_A0_O3(FAB2RAM_A_O[27]),
        .Tile_X9Y3_FAB2RAM_A1_O0(FAB2RAM_A_O[28]),
        .Tile_X9Y3_FAB2RAM_A1_O1(FAB2RAM_A_O[29]),
        .Tile_X9Y3_FAB2RAM_A1_O2(FAB2RAM_A_O[30]),
        .Tile_X9Y3_FAB2RAM_A1_O3(FAB2RAM_A_O[31]),
        .Tile_X9Y2_FAB2RAM_A0_O0(FAB2RAM_A_O[32]),
        .Tile_X9Y2_FAB2RAM_A0_O1(FAB2RAM_A_O[33]),
        .Tile_X9Y2_FAB2RAM_A0_O2(FAB2RAM_A_O[34]),
        .Tile_X9Y2_FAB2RAM_A0_O3(FAB2RAM_A_O[35]),
        .Tile_X9Y2_FAB2RAM_A1_O0(FAB2RAM_A_O[36]),
        .Tile_X9Y2_FAB2RAM_A1_O1(FAB2RAM_A_O[37]),
        .Tile_X9Y2_FAB2RAM_A1_O2(FAB2RAM_A_O[38]),
        .Tile_X9Y2_FAB2RAM_A1_O3(FAB2RAM_A_O[39]),
        .Tile_X9Y1_FAB2RAM_A0_O0(FAB2RAM_A_O[40]),
        .Tile_X9Y1_FAB2RAM_A0_O1(FAB2RAM_A_O[41]),
        .Tile_X9Y1_FAB2RAM_A0_O2(FAB2RAM_A_O[42]),
        .Tile_X9Y1_FAB2RAM_A0_O3(FAB2RAM_A_O[43]),
        .Tile_X9Y1_FAB2RAM_A1_O0(FAB2RAM_A_O[44]),
        .Tile_X9Y1_FAB2RAM_A1_O1(FAB2RAM_A_O[45]),
        .Tile_X9Y1_FAB2RAM_A1_O2(FAB2RAM_A_O[46]),
        .Tile_X9Y1_FAB2RAM_A1_O3(FAB2RAM_A_O[47]),
        .Tile_X9Y6_FAB2RAM_C_O0(FAB2RAM_C_O[0]),
        .Tile_X9Y6_FAB2RAM_C_O1(FAB2RAM_C_O[1]),
        .Tile_X9Y6_FAB2RAM_C_O2(FAB2RAM_C_O[2]),
        .Tile_X9Y6_FAB2RAM_C_O3(FAB2RAM_C_O[3]),
        .Tile_X9Y5_FAB2RAM_C_O0(FAB2RAM_C_O[4]),
        .Tile_X9Y5_FAB2RAM_C_O1(FAB2RAM_C_O[5]),
        .Tile_X9Y5_FAB2RAM_C_O2(FAB2RAM_C_O[6]),
        .Tile_X9Y5_FAB2RAM_C_O3(FAB2RAM_C_O[7]),
        .Tile_X9Y4_FAB2RAM_C_O0(FAB2RAM_C_O[8]),
        .Tile_X9Y4_FAB2RAM_C_O1(FAB2RAM_C_O[9]),
        .Tile_X9Y4_FAB2RAM_C_O2(FAB2RAM_C_O[10]),
        .Tile_X9Y4_FAB2RAM_C_O3(FAB2RAM_C_O[11]),
        .Tile_X9Y3_FAB2RAM_C_O0(FAB2RAM_C_O[12]),
        .Tile_X9Y3_FAB2RAM_C_O1(FAB2RAM_C_O[13]),
        .Tile_X9Y3_FAB2RAM_C_O2(FAB2RAM_C_O[14]),
        .Tile_X9Y3_FAB2RAM_C_O3(FAB2RAM_C_O[15]),
        .Tile_X9Y2_FAB2RAM_C_O0(FAB2RAM_C_O[16]),
        .Tile_X9Y2_FAB2RAM_C_O1(FAB2RAM_C_O[17]),
        .Tile_X9Y2_FAB2RAM_C_O2(FAB2RAM_C_O[18]),
        .Tile_X9Y2_FAB2RAM_C_O3(FAB2RAM_C_O[19]),
        .Tile_X9Y1_FAB2RAM_C_O0(FAB2RAM_C_O[20]),
        .Tile_X9Y1_FAB2RAM_C_O1(FAB2RAM_C_O[21]),
        .Tile_X9Y1_FAB2RAM_C_O2(FAB2RAM_C_O[22]),
        .Tile_X9Y1_FAB2RAM_C_O3(FAB2RAM_C_O[23]),
        .Tile_X9Y6_FAB2RAM_D0_O0(FAB2RAM_D_O[0]),
        .Tile_X9Y6_FAB2RAM_D0_O1(FAB2RAM_D_O[1]),
        .Tile_X9Y6_FAB2RAM_D0_O2(FAB2RAM_D_O[2]),
        .Tile_X9Y6_FAB2RAM_D0_O3(FAB2RAM_D_O[3]),
        .Tile_X9Y6_FAB2RAM_D1_O0(FAB2RAM_D_O[4]),
        .Tile_X9Y6_FAB2RAM_D1_O1(FAB2RAM_D_O[5]),
        .Tile_X9Y6_FAB2RAM_D1_O2(FAB2RAM_D_O[6]),
        .Tile_X9Y6_FAB2RAM_D1_O3(FAB2RAM_D_O[7]),
        .Tile_X9Y6_FAB2RAM_D2_O0(FAB2RAM_D_O[8]),
        .Tile_X9Y6_FAB2RAM_D2_O1(FAB2RAM_D_O[9]),
        .Tile_X9Y6_FAB2RAM_D2_O2(FAB2RAM_D_O[10]),
        .Tile_X9Y6_FAB2RAM_D2_O3(FAB2RAM_D_O[11]),
        .Tile_X9Y6_FAB2RAM_D3_O0(FAB2RAM_D_O[12]),
        .Tile_X9Y6_FAB2RAM_D3_O1(FAB2RAM_D_O[13]),
        .Tile_X9Y6_FAB2RAM_D3_O2(FAB2RAM_D_O[14]),
        .Tile_X9Y6_FAB2RAM_D3_O3(FAB2RAM_D_O[15]),
        .Tile_X9Y5_FAB2RAM_D0_O0(FAB2RAM_D_O[16]),
        .Tile_X9Y5_FAB2RAM_D0_O1(FAB2RAM_D_O[17]),
        .Tile_X9Y5_FAB2RAM_D0_O2(FAB2RAM_D_O[18]),
        .Tile_X9Y5_FAB2RAM_D0_O3(FAB2RAM_D_O[19]),
        .Tile_X9Y5_FAB2RAM_D1_O0(FAB2RAM_D_O[20]),
        .Tile_X9Y5_FAB2RAM_D1_O1(FAB2RAM_D_O[21]),
        .Tile_X9Y5_FAB2RAM_D1_O2(FAB2RAM_D_O[22]),
        .Tile_X9Y5_FAB2RAM_D1_O3(FAB2RAM_D_O[23]),
        .Tile_X9Y5_FAB2RAM_D2_O0(FAB2RAM_D_O[24]),
        .Tile_X9Y5_FAB2RAM_D2_O1(FAB2RAM_D_O[25]),
        .Tile_X9Y5_FAB2RAM_D2_O2(FAB2RAM_D_O[26]),
        .Tile_X9Y5_FAB2RAM_D2_O3(FAB2RAM_D_O[27]),
        .Tile_X9Y5_FAB2RAM_D3_O0(FAB2RAM_D_O[28]),
        .Tile_X9Y5_FAB2RAM_D3_O1(FAB2RAM_D_O[29]),
        .Tile_X9Y5_FAB2RAM_D3_O2(FAB2RAM_D_O[30]),
        .Tile_X9Y5_FAB2RAM_D3_O3(FAB2RAM_D_O[31]),
        .Tile_X9Y4_FAB2RAM_D0_O0(FAB2RAM_D_O[32]),
        .Tile_X9Y4_FAB2RAM_D0_O1(FAB2RAM_D_O[33]),
        .Tile_X9Y4_FAB2RAM_D0_O2(FAB2RAM_D_O[34]),
        .Tile_X9Y4_FAB2RAM_D0_O3(FAB2RAM_D_O[35]),
        .Tile_X9Y4_FAB2RAM_D1_O0(FAB2RAM_D_O[36]),
        .Tile_X9Y4_FAB2RAM_D1_O1(FAB2RAM_D_O[37]),
        .Tile_X9Y4_FAB2RAM_D1_O2(FAB2RAM_D_O[38]),
        .Tile_X9Y4_FAB2RAM_D1_O3(FAB2RAM_D_O[39]),
        .Tile_X9Y4_FAB2RAM_D2_O0(FAB2RAM_D_O[40]),
        .Tile_X9Y4_FAB2RAM_D2_O1(FAB2RAM_D_O[41]),
        .Tile_X9Y4_FAB2RAM_D2_O2(FAB2RAM_D_O[42]),
        .Tile_X9Y4_FAB2RAM_D2_O3(FAB2RAM_D_O[43]),
        .Tile_X9Y4_FAB2RAM_D3_O0(FAB2RAM_D_O[44]),
        .Tile_X9Y4_FAB2RAM_D3_O1(FAB2RAM_D_O[45]),
        .Tile_X9Y4_FAB2RAM_D3_O2(FAB2RAM_D_O[46]),
        .Tile_X9Y4_FAB2RAM_D3_O3(FAB2RAM_D_O[47]),
        .Tile_X9Y3_FAB2RAM_D0_O0(FAB2RAM_D_O[48]),
        .Tile_X9Y3_FAB2RAM_D0_O1(FAB2RAM_D_O[49]),
        .Tile_X9Y3_FAB2RAM_D0_O2(FAB2RAM_D_O[50]),
        .Tile_X9Y3_FAB2RAM_D0_O3(FAB2RAM_D_O[51]),
        .Tile_X9Y3_FAB2RAM_D1_O0(FAB2RAM_D_O[52]),
        .Tile_X9Y3_FAB2RAM_D1_O1(FAB2RAM_D_O[53]),
        .Tile_X9Y3_FAB2RAM_D1_O2(FAB2RAM_D_O[54]),
        .Tile_X9Y3_FAB2RAM_D1_O3(FAB2RAM_D_O[55]),
        .Tile_X9Y3_FAB2RAM_D2_O0(FAB2RAM_D_O[56]),
        .Tile_X9Y3_FAB2RAM_D2_O1(FAB2RAM_D_O[57]),
        .Tile_X9Y3_FAB2RAM_D2_O2(FAB2RAM_D_O[58]),
        .Tile_X9Y3_FAB2RAM_D2_O3(FAB2RAM_D_O[59]),
        .Tile_X9Y3_FAB2RAM_D3_O0(FAB2RAM_D_O[60]),
        .Tile_X9Y3_FAB2RAM_D3_O1(FAB2RAM_D_O[61]),
        .Tile_X9Y3_FAB2RAM_D3_O2(FAB2RAM_D_O[62]),
        .Tile_X9Y3_FAB2RAM_D3_O3(FAB2RAM_D_O[63]),
        .Tile_X9Y2_FAB2RAM_D0_O0(FAB2RAM_D_O[64]),
        .Tile_X9Y2_FAB2RAM_D0_O1(FAB2RAM_D_O[65]),
        .Tile_X9Y2_FAB2RAM_D0_O2(FAB2RAM_D_O[66]),
        .Tile_X9Y2_FAB2RAM_D0_O3(FAB2RAM_D_O[67]),
        .Tile_X9Y2_FAB2RAM_D1_O0(FAB2RAM_D_O[68]),
        .Tile_X9Y2_FAB2RAM_D1_O1(FAB2RAM_D_O[69]),
        .Tile_X9Y2_FAB2RAM_D1_O2(FAB2RAM_D_O[70]),
        .Tile_X9Y2_FAB2RAM_D1_O3(FAB2RAM_D_O[71]),
        .Tile_X9Y2_FAB2RAM_D2_O0(FAB2RAM_D_O[72]),
        .Tile_X9Y2_FAB2RAM_D2_O1(FAB2RAM_D_O[73]),
        .Tile_X9Y2_FAB2RAM_D2_O2(FAB2RAM_D_O[74]),
        .Tile_X9Y2_FAB2RAM_D2_O3(FAB2RAM_D_O[75]),
        .Tile_X9Y2_FAB2RAM_D3_O0(FAB2RAM_D_O[76]),
        .Tile_X9Y2_FAB2RAM_D3_O1(FAB2RAM_D_O[77]),
        .Tile_X9Y2_FAB2RAM_D3_O2(FAB2RAM_D_O[78]),
        .Tile_X9Y2_FAB2RAM_D3_O3(FAB2RAM_D_O[79]),
        .Tile_X9Y1_FAB2RAM_D0_O0(FAB2RAM_D_O[80]),
        .Tile_X9Y1_FAB2RAM_D0_O1(FAB2RAM_D_O[81]),
        .Tile_X9Y1_FAB2RAM_D0_O2(FAB2RAM_D_O[82]),
        .Tile_X9Y1_FAB2RAM_D0_O3(FAB2RAM_D_O[83]),
        .Tile_X9Y1_FAB2RAM_D1_O0(FAB2RAM_D_O[84]),
        .Tile_X9Y1_FAB2RAM_D1_O1(FAB2RAM_D_O[85]),
        .Tile_X9Y1_FAB2RAM_D1_O2(FAB2RAM_D_O[86]),
        .Tile_X9Y1_FAB2RAM_D1_O3(FAB2RAM_D_O[87]),
        .Tile_X9Y1_FAB2RAM_D2_O0(FAB2RAM_D_O[88]),
        .Tile_X9Y1_FAB2RAM_D2_O1(FAB2RAM_D_O[89]),
        .Tile_X9Y1_FAB2RAM_D2_O2(FAB2RAM_D_O[90]),
        .Tile_X9Y1_FAB2RAM_D2_O3(FAB2RAM_D_O[91]),
        .Tile_X9Y1_FAB2RAM_D3_O0(FAB2RAM_D_O[92]),
        .Tile_X9Y1_FAB2RAM_D3_O1(FAB2RAM_D_O[93]),
        .Tile_X9Y1_FAB2RAM_D3_O2(FAB2RAM_D_O[94]),
        .Tile_X9Y1_FAB2RAM_D3_O3(FAB2RAM_D_O[95]),
        .Tile_X0Y6_B_I_top(I_top[0]),
        .Tile_X0Y6_A_I_top(I_top[1]),
        .Tile_X0Y5_B_I_top(I_top[2]),
        .Tile_X0Y5_A_I_top(I_top[3]),
        .Tile_X0Y4_B_I_top(I_top[4]),
        .Tile_X0Y4_A_I_top(I_top[5]),
        .Tile_X0Y3_B_I_top(I_top[6]),
        .Tile_X0Y3_A_I_top(I_top[7]),
        .Tile_X0Y2_B_I_top(I_top[8]),
        .Tile_X0Y2_A_I_top(I_top[9]),
        .Tile_X0Y1_B_I_top(I_top[10]),
        .Tile_X0Y1_A_I_top(I_top[11]),
        .Tile_X0Y6_B_O_top(O_top[0]),
        .Tile_X0Y6_A_O_top(O_top[1]),
        .Tile_X0Y5_B_O_top(O_top[2]),
        .Tile_X0Y5_A_O_top(O_top[3]),
        .Tile_X0Y4_B_O_top(O_top[4]),
        .Tile_X0Y4_A_O_top(O_top[5]),
        .Tile_X0Y3_B_O_top(O_top[6]),
        .Tile_X0Y3_A_O_top(O_top[7]),
        .Tile_X0Y2_B_O_top(O_top[8]),
        .Tile_X0Y2_A_O_top(O_top[9]),
        .Tile_X0Y1_B_O_top(O_top[10]),
        .Tile_X0Y1_A_O_top(O_top[11]),
        .Tile_X9Y6_RAM2FAB_D0_I0(RAM2FAB_D_I[0]),
        .Tile_X9Y6_RAM2FAB_D0_I1(RAM2FAB_D_I[1]),
        .Tile_X9Y6_RAM2FAB_D0_I2(RAM2FAB_D_I[2]),
        .Tile_X9Y6_RAM2FAB_D0_I3(RAM2FAB_D_I[3]),
        .Tile_X9Y6_RAM2FAB_D1_I0(RAM2FAB_D_I[4]),
        .Tile_X9Y6_RAM2FAB_D1_I1(RAM2FAB_D_I[5]),
        .Tile_X9Y6_RAM2FAB_D1_I2(RAM2FAB_D_I[6]),
        .Tile_X9Y6_RAM2FAB_D1_I3(RAM2FAB_D_I[7]),
        .Tile_X9Y6_RAM2FAB_D2_I0(RAM2FAB_D_I[8]),
        .Tile_X9Y6_RAM2FAB_D2_I1(RAM2FAB_D_I[9]),
        .Tile_X9Y6_RAM2FAB_D2_I2(RAM2FAB_D_I[10]),
        .Tile_X9Y6_RAM2FAB_D2_I3(RAM2FAB_D_I[11]),
        .Tile_X9Y6_RAM2FAB_D3_I0(RAM2FAB_D_I[12]),
        .Tile_X9Y6_RAM2FAB_D3_I1(RAM2FAB_D_I[13]),
        .Tile_X9Y6_RAM2FAB_D3_I2(RAM2FAB_D_I[14]),
        .Tile_X9Y6_RAM2FAB_D3_I3(RAM2FAB_D_I[15]),
        .Tile_X9Y5_RAM2FAB_D0_I0(RAM2FAB_D_I[16]),
        .Tile_X9Y5_RAM2FAB_D0_I1(RAM2FAB_D_I[17]),
        .Tile_X9Y5_RAM2FAB_D0_I2(RAM2FAB_D_I[18]),
        .Tile_X9Y5_RAM2FAB_D0_I3(RAM2FAB_D_I[19]),
        .Tile_X9Y5_RAM2FAB_D1_I0(RAM2FAB_D_I[20]),
        .Tile_X9Y5_RAM2FAB_D1_I1(RAM2FAB_D_I[21]),
        .Tile_X9Y5_RAM2FAB_D1_I2(RAM2FAB_D_I[22]),
        .Tile_X9Y5_RAM2FAB_D1_I3(RAM2FAB_D_I[23]),
        .Tile_X9Y5_RAM2FAB_D2_I0(RAM2FAB_D_I[24]),
        .Tile_X9Y5_RAM2FAB_D2_I1(RAM2FAB_D_I[25]),
        .Tile_X9Y5_RAM2FAB_D2_I2(RAM2FAB_D_I[26]),
        .Tile_X9Y5_RAM2FAB_D2_I3(RAM2FAB_D_I[27]),
        .Tile_X9Y5_RAM2FAB_D3_I0(RAM2FAB_D_I[28]),
        .Tile_X9Y5_RAM2FAB_D3_I1(RAM2FAB_D_I[29]),
        .Tile_X9Y5_RAM2FAB_D3_I2(RAM2FAB_D_I[30]),
        .Tile_X9Y5_RAM2FAB_D3_I3(RAM2FAB_D_I[31]),
        .Tile_X9Y4_RAM2FAB_D0_I0(RAM2FAB_D_I[32]),
        .Tile_X9Y4_RAM2FAB_D0_I1(RAM2FAB_D_I[33]),
        .Tile_X9Y4_RAM2FAB_D0_I2(RAM2FAB_D_I[34]),
        .Tile_X9Y4_RAM2FAB_D0_I3(RAM2FAB_D_I[35]),
        .Tile_X9Y4_RAM2FAB_D1_I0(RAM2FAB_D_I[36]),
        .Tile_X9Y4_RAM2FAB_D1_I1(RAM2FAB_D_I[37]),
        .Tile_X9Y4_RAM2FAB_D1_I2(RAM2FAB_D_I[38]),
        .Tile_X9Y4_RAM2FAB_D1_I3(RAM2FAB_D_I[39]),
        .Tile_X9Y4_RAM2FAB_D2_I0(RAM2FAB_D_I[40]),
        .Tile_X9Y4_RAM2FAB_D2_I1(RAM2FAB_D_I[41]),
        .Tile_X9Y4_RAM2FAB_D2_I2(RAM2FAB_D_I[42]),
        .Tile_X9Y4_RAM2FAB_D2_I3(RAM2FAB_D_I[43]),
        .Tile_X9Y4_RAM2FAB_D3_I0(RAM2FAB_D_I[44]),
        .Tile_X9Y4_RAM2FAB_D3_I1(RAM2FAB_D_I[45]),
        .Tile_X9Y4_RAM2FAB_D3_I2(RAM2FAB_D_I[46]),
        .Tile_X9Y4_RAM2FAB_D3_I3(RAM2FAB_D_I[47]),
        .Tile_X9Y3_RAM2FAB_D0_I0(RAM2FAB_D_I[48]),
        .Tile_X9Y3_RAM2FAB_D0_I1(RAM2FAB_D_I[49]),
        .Tile_X9Y3_RAM2FAB_D0_I2(RAM2FAB_D_I[50]),
        .Tile_X9Y3_RAM2FAB_D0_I3(RAM2FAB_D_I[51]),
        .Tile_X9Y3_RAM2FAB_D1_I0(RAM2FAB_D_I[52]),
        .Tile_X9Y3_RAM2FAB_D1_I1(RAM2FAB_D_I[53]),
        .Tile_X9Y3_RAM2FAB_D1_I2(RAM2FAB_D_I[54]),
        .Tile_X9Y3_RAM2FAB_D1_I3(RAM2FAB_D_I[55]),
        .Tile_X9Y3_RAM2FAB_D2_I0(RAM2FAB_D_I[56]),
        .Tile_X9Y3_RAM2FAB_D2_I1(RAM2FAB_D_I[57]),
        .Tile_X9Y3_RAM2FAB_D2_I2(RAM2FAB_D_I[58]),
        .Tile_X9Y3_RAM2FAB_D2_I3(RAM2FAB_D_I[59]),
        .Tile_X9Y3_RAM2FAB_D3_I0(RAM2FAB_D_I[60]),
        .Tile_X9Y3_RAM2FAB_D3_I1(RAM2FAB_D_I[61]),
        .Tile_X9Y3_RAM2FAB_D3_I2(RAM2FAB_D_I[62]),
        .Tile_X9Y3_RAM2FAB_D3_I3(RAM2FAB_D_I[63]),
        .Tile_X9Y2_RAM2FAB_D0_I0(RAM2FAB_D_I[64]),
        .Tile_X9Y2_RAM2FAB_D0_I1(RAM2FAB_D_I[65]),
        .Tile_X9Y2_RAM2FAB_D0_I2(RAM2FAB_D_I[66]),
        .Tile_X9Y2_RAM2FAB_D0_I3(RAM2FAB_D_I[67]),
        .Tile_X9Y2_RAM2FAB_D1_I0(RAM2FAB_D_I[68]),
        .Tile_X9Y2_RAM2FAB_D1_I1(RAM2FAB_D_I[69]),
        .Tile_X9Y2_RAM2FAB_D1_I2(RAM2FAB_D_I[70]),
        .Tile_X9Y2_RAM2FAB_D1_I3(RAM2FAB_D_I[71]),
        .Tile_X9Y2_RAM2FAB_D2_I0(RAM2FAB_D_I[72]),
        .Tile_X9Y2_RAM2FAB_D2_I1(RAM2FAB_D_I[73]),
        .Tile_X9Y2_RAM2FAB_D2_I2(RAM2FAB_D_I[74]),
        .Tile_X9Y2_RAM2FAB_D2_I3(RAM2FAB_D_I[75]),
        .Tile_X9Y2_RAM2FAB_D3_I0(RAM2FAB_D_I[76]),
        .Tile_X9Y2_RAM2FAB_D3_I1(RAM2FAB_D_I[77]),
        .Tile_X9Y2_RAM2FAB_D3_I2(RAM2FAB_D_I[78]),
        .Tile_X9Y2_RAM2FAB_D3_I3(RAM2FAB_D_I[79]),
        .Tile_X9Y1_RAM2FAB_D0_I0(RAM2FAB_D_I[80]),
        .Tile_X9Y1_RAM2FAB_D0_I1(RAM2FAB_D_I[81]),
        .Tile_X9Y1_RAM2FAB_D0_I2(RAM2FAB_D_I[82]),
        .Tile_X9Y1_RAM2FAB_D0_I3(RAM2FAB_D_I[83]),
        .Tile_X9Y1_RAM2FAB_D1_I0(RAM2FAB_D_I[84]),
        .Tile_X9Y1_RAM2FAB_D1_I1(RAM2FAB_D_I[85]),
        .Tile_X9Y1_RAM2FAB_D1_I2(RAM2FAB_D_I[86]),
        .Tile_X9Y1_RAM2FAB_D1_I3(RAM2FAB_D_I[87]),
        .Tile_X9Y1_RAM2FAB_D2_I0(RAM2FAB_D_I[88]),
        .Tile_X9Y1_RAM2FAB_D2_I1(RAM2FAB_D_I[89]),
        .Tile_X9Y1_RAM2FAB_D2_I2(RAM2FAB_D_I[90]),
        .Tile_X9Y1_RAM2FAB_D2_I3(RAM2FAB_D_I[91]),
        .Tile_X9Y1_RAM2FAB_D3_I0(RAM2FAB_D_I[92]),
        .Tile_X9Y1_RAM2FAB_D3_I1(RAM2FAB_D_I[93]),
        .Tile_X9Y1_RAM2FAB_D3_I2(RAM2FAB_D_I[94]),
        .Tile_X9Y1_RAM2FAB_D3_I3(RAM2FAB_D_I[95]),
        .Tile_X0Y6_B_T_top(T_top[0]),
        .Tile_X0Y6_A_T_top(T_top[1]),
        .Tile_X0Y5_B_T_top(T_top[2]),
        .Tile_X0Y5_A_T_top(T_top[3]),
        .Tile_X0Y4_B_T_top(T_top[4]),
        .Tile_X0Y4_A_T_top(T_top[5]),
        .Tile_X0Y3_B_T_top(T_top[6]),
        .Tile_X0Y3_A_T_top(T_top[7]),
        .Tile_X0Y2_B_T_top(T_top[8]),
        .Tile_X0Y2_A_T_top(T_top[9]),
        .Tile_X0Y1_B_T_top(T_top[10]),
        .Tile_X0Y1_A_T_top(T_top[11]),
        .Tile_X1Y7_UIO_BOT_UIN0(UIO_BOT_UIN[0]),
        .Tile_X1Y7_UIO_BOT_UIN1(UIO_BOT_UIN[1]),
        .Tile_X1Y7_UIO_BOT_UIN2(UIO_BOT_UIN[2]),
        .Tile_X1Y7_UIO_BOT_UIN3(UIO_BOT_UIN[3]),
        .Tile_X1Y7_UIO_BOT_UIN4(UIO_BOT_UIN[4]),
        .Tile_X1Y7_UIO_BOT_UIN5(UIO_BOT_UIN[5]),
        .Tile_X1Y7_UIO_BOT_UIN6(UIO_BOT_UIN[6]),
        .Tile_X1Y7_UIO_BOT_UIN7(UIO_BOT_UIN[7]),
        .Tile_X1Y7_UIO_BOT_UIN8(UIO_BOT_UIN[8]),
        .Tile_X1Y7_UIO_BOT_UIN9(UIO_BOT_UIN[9]),
        .Tile_X1Y7_UIO_BOT_UIN10(UIO_BOT_UIN[10]),
        .Tile_X1Y7_UIO_BOT_UIN11(UIO_BOT_UIN[11]),
        .Tile_X1Y7_UIO_BOT_UIN12(UIO_BOT_UIN[12]),
        .Tile_X1Y7_UIO_BOT_UIN13(UIO_BOT_UIN[13]),
        .Tile_X1Y7_UIO_BOT_UIN14(UIO_BOT_UIN[14]),
        .Tile_X1Y7_UIO_BOT_UIN15(UIO_BOT_UIN[15]),
        .Tile_X1Y7_UIO_BOT_UIN16(UIO_BOT_UIN[16]),
        .Tile_X1Y7_UIO_BOT_UIN17(UIO_BOT_UIN[17]),
        .Tile_X1Y7_UIO_BOT_UIN18(UIO_BOT_UIN[18]),
        .Tile_X1Y7_UIO_BOT_UIN19(UIO_BOT_UIN[19]),
        .Tile_X2Y7_UIO_BOT_UIN0(UIO_BOT_UIN[20]),
        .Tile_X2Y7_UIO_BOT_UIN1(UIO_BOT_UIN[21]),
        .Tile_X2Y7_UIO_BOT_UIN2(UIO_BOT_UIN[22]),
        .Tile_X2Y7_UIO_BOT_UIN3(UIO_BOT_UIN[23]),
        .Tile_X2Y7_UIO_BOT_UIN4(UIO_BOT_UIN[24]),
        .Tile_X2Y7_UIO_BOT_UIN5(UIO_BOT_UIN[25]),
        .Tile_X2Y7_UIO_BOT_UIN6(UIO_BOT_UIN[26]),
        .Tile_X2Y7_UIO_BOT_UIN7(UIO_BOT_UIN[27]),
        .Tile_X2Y7_UIO_BOT_UIN8(UIO_BOT_UIN[28]),
        .Tile_X2Y7_UIO_BOT_UIN9(UIO_BOT_UIN[29]),
        .Tile_X2Y7_UIO_BOT_UIN10(UIO_BOT_UIN[30]),
        .Tile_X2Y7_UIO_BOT_UIN11(UIO_BOT_UIN[31]),
        .Tile_X2Y7_UIO_BOT_UIN12(UIO_BOT_UIN[32]),
        .Tile_X2Y7_UIO_BOT_UIN13(UIO_BOT_UIN[33]),
        .Tile_X2Y7_UIO_BOT_UIN14(UIO_BOT_UIN[34]),
        .Tile_X2Y7_UIO_BOT_UIN15(UIO_BOT_UIN[35]),
        .Tile_X2Y7_UIO_BOT_UIN16(UIO_BOT_UIN[36]),
        .Tile_X2Y7_UIO_BOT_UIN17(UIO_BOT_UIN[37]),
        .Tile_X2Y7_UIO_BOT_UIN18(UIO_BOT_UIN[38]),
        .Tile_X2Y7_UIO_BOT_UIN19(UIO_BOT_UIN[39]),
        .Tile_X3Y7_UIO_BOT_UIN0(UIO_BOT_UIN[40]),
        .Tile_X3Y7_UIO_BOT_UIN1(UIO_BOT_UIN[41]),
        .Tile_X3Y7_UIO_BOT_UIN2(UIO_BOT_UIN[42]),
        .Tile_X3Y7_UIO_BOT_UIN3(UIO_BOT_UIN[43]),
        .Tile_X3Y7_UIO_BOT_UIN4(UIO_BOT_UIN[44]),
        .Tile_X3Y7_UIO_BOT_UIN5(UIO_BOT_UIN[45]),
        .Tile_X3Y7_UIO_BOT_UIN6(UIO_BOT_UIN[46]),
        .Tile_X3Y7_UIO_BOT_UIN7(UIO_BOT_UIN[47]),
        .Tile_X3Y7_UIO_BOT_UIN8(UIO_BOT_UIN[48]),
        .Tile_X3Y7_UIO_BOT_UIN9(UIO_BOT_UIN[49]),
        .Tile_X3Y7_UIO_BOT_UIN10(UIO_BOT_UIN[50]),
        .Tile_X3Y7_UIO_BOT_UIN11(UIO_BOT_UIN[51]),
        .Tile_X3Y7_UIO_BOT_UIN12(UIO_BOT_UIN[52]),
        .Tile_X3Y7_UIO_BOT_UIN13(UIO_BOT_UIN[53]),
        .Tile_X3Y7_UIO_BOT_UIN14(UIO_BOT_UIN[54]),
        .Tile_X3Y7_UIO_BOT_UIN15(UIO_BOT_UIN[55]),
        .Tile_X3Y7_UIO_BOT_UIN16(UIO_BOT_UIN[56]),
        .Tile_X3Y7_UIO_BOT_UIN17(UIO_BOT_UIN[57]),
        .Tile_X3Y7_UIO_BOT_UIN18(UIO_BOT_UIN[58]),
        .Tile_X3Y7_UIO_BOT_UIN19(UIO_BOT_UIN[59]),
        .Tile_X4Y7_UIO_BOT_UIN0(UIO_BOT_UIN[60]),
        .Tile_X4Y7_UIO_BOT_UIN1(UIO_BOT_UIN[61]),
        .Tile_X4Y7_UIO_BOT_UIN2(UIO_BOT_UIN[62]),
        .Tile_X4Y7_UIO_BOT_UIN3(UIO_BOT_UIN[63]),
        .Tile_X4Y7_UIO_BOT_UIN4(UIO_BOT_UIN[64]),
        .Tile_X4Y7_UIO_BOT_UIN5(UIO_BOT_UIN[65]),
        .Tile_X4Y7_UIO_BOT_UIN6(UIO_BOT_UIN[66]),
        .Tile_X4Y7_UIO_BOT_UIN7(UIO_BOT_UIN[67]),
        .Tile_X4Y7_UIO_BOT_UIN8(UIO_BOT_UIN[68]),
        .Tile_X4Y7_UIO_BOT_UIN9(UIO_BOT_UIN[69]),
        .Tile_X4Y7_UIO_BOT_UIN10(UIO_BOT_UIN[70]),
        .Tile_X4Y7_UIO_BOT_UIN11(UIO_BOT_UIN[71]),
        .Tile_X4Y7_UIO_BOT_UIN12(UIO_BOT_UIN[72]),
        .Tile_X4Y7_UIO_BOT_UIN13(UIO_BOT_UIN[73]),
        .Tile_X4Y7_UIO_BOT_UIN14(UIO_BOT_UIN[74]),
        .Tile_X4Y7_UIO_BOT_UIN15(UIO_BOT_UIN[75]),
        .Tile_X4Y7_UIO_BOT_UIN16(UIO_BOT_UIN[76]),
        .Tile_X4Y7_UIO_BOT_UIN17(UIO_BOT_UIN[77]),
        .Tile_X4Y7_UIO_BOT_UIN18(UIO_BOT_UIN[78]),
        .Tile_X4Y7_UIO_BOT_UIN19(UIO_BOT_UIN[79]),
        .Tile_X5Y7_UIO_BOT_UIN0(UIO_BOT_UIN[80]),
        .Tile_X5Y7_UIO_BOT_UIN1(UIO_BOT_UIN[81]),
        .Tile_X5Y7_UIO_BOT_UIN2(UIO_BOT_UIN[82]),
        .Tile_X5Y7_UIO_BOT_UIN3(UIO_BOT_UIN[83]),
        .Tile_X5Y7_UIO_BOT_UIN4(UIO_BOT_UIN[84]),
        .Tile_X5Y7_UIO_BOT_UIN5(UIO_BOT_UIN[85]),
        .Tile_X5Y7_UIO_BOT_UIN6(UIO_BOT_UIN[86]),
        .Tile_X5Y7_UIO_BOT_UIN7(UIO_BOT_UIN[87]),
        .Tile_X5Y7_UIO_BOT_UIN8(UIO_BOT_UIN[88]),
        .Tile_X5Y7_UIO_BOT_UIN9(UIO_BOT_UIN[89]),
        .Tile_X5Y7_UIO_BOT_UIN10(UIO_BOT_UIN[90]),
        .Tile_X5Y7_UIO_BOT_UIN11(UIO_BOT_UIN[91]),
        .Tile_X5Y7_UIO_BOT_UIN12(UIO_BOT_UIN[92]),
        .Tile_X5Y7_UIO_BOT_UIN13(UIO_BOT_UIN[93]),
        .Tile_X5Y7_UIO_BOT_UIN14(UIO_BOT_UIN[94]),
        .Tile_X5Y7_UIO_BOT_UIN15(UIO_BOT_UIN[95]),
        .Tile_X5Y7_UIO_BOT_UIN16(UIO_BOT_UIN[96]),
        .Tile_X5Y7_UIO_BOT_UIN17(UIO_BOT_UIN[97]),
        .Tile_X5Y7_UIO_BOT_UIN18(UIO_BOT_UIN[98]),
        .Tile_X5Y7_UIO_BOT_UIN19(UIO_BOT_UIN[99]),
        .Tile_X6Y7_UIO_BOT_UIN0(UIO_BOT_UIN[100]),
        .Tile_X6Y7_UIO_BOT_UIN1(UIO_BOT_UIN[101]),
        .Tile_X6Y7_UIO_BOT_UIN2(UIO_BOT_UIN[102]),
        .Tile_X6Y7_UIO_BOT_UIN3(UIO_BOT_UIN[103]),
        .Tile_X6Y7_UIO_BOT_UIN4(UIO_BOT_UIN[104]),
        .Tile_X6Y7_UIO_BOT_UIN5(UIO_BOT_UIN[105]),
        .Tile_X6Y7_UIO_BOT_UIN6(UIO_BOT_UIN[106]),
        .Tile_X6Y7_UIO_BOT_UIN7(UIO_BOT_UIN[107]),
        .Tile_X6Y7_UIO_BOT_UIN8(UIO_BOT_UIN[108]),
        .Tile_X6Y7_UIO_BOT_UIN9(UIO_BOT_UIN[109]),
        .Tile_X6Y7_UIO_BOT_UIN10(UIO_BOT_UIN[110]),
        .Tile_X6Y7_UIO_BOT_UIN11(UIO_BOT_UIN[111]),
        .Tile_X6Y7_UIO_BOT_UIN12(UIO_BOT_UIN[112]),
        .Tile_X6Y7_UIO_BOT_UIN13(UIO_BOT_UIN[113]),
        .Tile_X6Y7_UIO_BOT_UIN14(UIO_BOT_UIN[114]),
        .Tile_X6Y7_UIO_BOT_UIN15(UIO_BOT_UIN[115]),
        .Tile_X6Y7_UIO_BOT_UIN16(UIO_BOT_UIN[116]),
        .Tile_X6Y7_UIO_BOT_UIN17(UIO_BOT_UIN[117]),
        .Tile_X6Y7_UIO_BOT_UIN18(UIO_BOT_UIN[118]),
        .Tile_X6Y7_UIO_BOT_UIN19(UIO_BOT_UIN[119]),
        .Tile_X7Y7_UIO_BOT_UIN0(UIO_BOT_UIN[120]),
        .Tile_X7Y7_UIO_BOT_UIN1(UIO_BOT_UIN[121]),
        .Tile_X7Y7_UIO_BOT_UIN2(UIO_BOT_UIN[122]),
        .Tile_X7Y7_UIO_BOT_UIN3(UIO_BOT_UIN[123]),
        .Tile_X7Y7_UIO_BOT_UIN4(UIO_BOT_UIN[124]),
        .Tile_X7Y7_UIO_BOT_UIN5(UIO_BOT_UIN[125]),
        .Tile_X7Y7_UIO_BOT_UIN6(UIO_BOT_UIN[126]),
        .Tile_X7Y7_UIO_BOT_UIN7(UIO_BOT_UIN[127]),
        .Tile_X7Y7_UIO_BOT_UIN8(UIO_BOT_UIN[128]),
        .Tile_X7Y7_UIO_BOT_UIN9(UIO_BOT_UIN[129]),
        .Tile_X7Y7_UIO_BOT_UIN10(UIO_BOT_UIN[130]),
        .Tile_X7Y7_UIO_BOT_UIN11(UIO_BOT_UIN[131]),
        .Tile_X7Y7_UIO_BOT_UIN12(UIO_BOT_UIN[132]),
        .Tile_X7Y7_UIO_BOT_UIN13(UIO_BOT_UIN[133]),
        .Tile_X7Y7_UIO_BOT_UIN14(UIO_BOT_UIN[134]),
        .Tile_X7Y7_UIO_BOT_UIN15(UIO_BOT_UIN[135]),
        .Tile_X7Y7_UIO_BOT_UIN16(UIO_BOT_UIN[136]),
        .Tile_X7Y7_UIO_BOT_UIN17(UIO_BOT_UIN[137]),
        .Tile_X7Y7_UIO_BOT_UIN18(UIO_BOT_UIN[138]),
        .Tile_X7Y7_UIO_BOT_UIN19(UIO_BOT_UIN[139]),
        .Tile_X8Y7_UIO_BOT_UIN0(UIO_BOT_UIN[140]),
        .Tile_X8Y7_UIO_BOT_UIN1(UIO_BOT_UIN[141]),
        .Tile_X8Y7_UIO_BOT_UIN2(UIO_BOT_UIN[142]),
        .Tile_X8Y7_UIO_BOT_UIN3(UIO_BOT_UIN[143]),
        .Tile_X8Y7_UIO_BOT_UIN4(UIO_BOT_UIN[144]),
        .Tile_X8Y7_UIO_BOT_UIN5(UIO_BOT_UIN[145]),
        .Tile_X8Y7_UIO_BOT_UIN6(UIO_BOT_UIN[146]),
        .Tile_X8Y7_UIO_BOT_UIN7(UIO_BOT_UIN[147]),
        .Tile_X8Y7_UIO_BOT_UIN8(UIO_BOT_UIN[148]),
        .Tile_X8Y7_UIO_BOT_UIN9(UIO_BOT_UIN[149]),
        .Tile_X8Y7_UIO_BOT_UIN10(UIO_BOT_UIN[150]),
        .Tile_X8Y7_UIO_BOT_UIN11(UIO_BOT_UIN[151]),
        .Tile_X8Y7_UIO_BOT_UIN12(UIO_BOT_UIN[152]),
        .Tile_X8Y7_UIO_BOT_UIN13(UIO_BOT_UIN[153]),
        .Tile_X8Y7_UIO_BOT_UIN14(UIO_BOT_UIN[154]),
        .Tile_X8Y7_UIO_BOT_UIN15(UIO_BOT_UIN[155]),
        .Tile_X8Y7_UIO_BOT_UIN16(UIO_BOT_UIN[156]),
        .Tile_X8Y7_UIO_BOT_UIN17(UIO_BOT_UIN[157]),
        .Tile_X8Y7_UIO_BOT_UIN18(UIO_BOT_UIN[158]),
        .Tile_X8Y7_UIO_BOT_UIN19(UIO_BOT_UIN[159]),
        .Tile_X1Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[0]),
        .Tile_X1Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[1]),
        .Tile_X1Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[2]),
        .Tile_X1Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[3]),
        .Tile_X1Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[4]),
        .Tile_X1Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[5]),
        .Tile_X1Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[6]),
        .Tile_X1Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[7]),
        .Tile_X1Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[8]),
        .Tile_X1Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[9]),
        .Tile_X1Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[10]),
        .Tile_X1Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[11]),
        .Tile_X1Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[12]),
        .Tile_X1Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[13]),
        .Tile_X1Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[14]),
        .Tile_X1Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[15]),
        .Tile_X1Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[16]),
        .Tile_X1Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[17]),
        .Tile_X1Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[18]),
        .Tile_X1Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[19]),
        .Tile_X2Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[20]),
        .Tile_X2Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[21]),
        .Tile_X2Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[22]),
        .Tile_X2Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[23]),
        .Tile_X2Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[24]),
        .Tile_X2Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[25]),
        .Tile_X2Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[26]),
        .Tile_X2Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[27]),
        .Tile_X2Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[28]),
        .Tile_X2Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[29]),
        .Tile_X2Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[30]),
        .Tile_X2Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[31]),
        .Tile_X2Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[32]),
        .Tile_X2Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[33]),
        .Tile_X2Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[34]),
        .Tile_X2Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[35]),
        .Tile_X2Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[36]),
        .Tile_X2Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[37]),
        .Tile_X2Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[38]),
        .Tile_X2Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[39]),
        .Tile_X3Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[40]),
        .Tile_X3Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[41]),
        .Tile_X3Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[42]),
        .Tile_X3Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[43]),
        .Tile_X3Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[44]),
        .Tile_X3Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[45]),
        .Tile_X3Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[46]),
        .Tile_X3Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[47]),
        .Tile_X3Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[48]),
        .Tile_X3Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[49]),
        .Tile_X3Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[50]),
        .Tile_X3Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[51]),
        .Tile_X3Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[52]),
        .Tile_X3Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[53]),
        .Tile_X3Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[54]),
        .Tile_X3Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[55]),
        .Tile_X3Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[56]),
        .Tile_X3Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[57]),
        .Tile_X3Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[58]),
        .Tile_X3Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[59]),
        .Tile_X4Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[60]),
        .Tile_X4Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[61]),
        .Tile_X4Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[62]),
        .Tile_X4Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[63]),
        .Tile_X4Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[64]),
        .Tile_X4Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[65]),
        .Tile_X4Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[66]),
        .Tile_X4Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[67]),
        .Tile_X4Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[68]),
        .Tile_X4Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[69]),
        .Tile_X4Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[70]),
        .Tile_X4Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[71]),
        .Tile_X4Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[72]),
        .Tile_X4Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[73]),
        .Tile_X4Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[74]),
        .Tile_X4Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[75]),
        .Tile_X4Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[76]),
        .Tile_X4Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[77]),
        .Tile_X4Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[78]),
        .Tile_X4Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[79]),
        .Tile_X5Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[80]),
        .Tile_X5Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[81]),
        .Tile_X5Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[82]),
        .Tile_X5Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[83]),
        .Tile_X5Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[84]),
        .Tile_X5Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[85]),
        .Tile_X5Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[86]),
        .Tile_X5Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[87]),
        .Tile_X5Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[88]),
        .Tile_X5Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[89]),
        .Tile_X5Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[90]),
        .Tile_X5Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[91]),
        .Tile_X5Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[92]),
        .Tile_X5Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[93]),
        .Tile_X5Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[94]),
        .Tile_X5Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[95]),
        .Tile_X5Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[96]),
        .Tile_X5Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[97]),
        .Tile_X5Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[98]),
        .Tile_X5Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[99]),
        .Tile_X6Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[100]),
        .Tile_X6Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[101]),
        .Tile_X6Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[102]),
        .Tile_X6Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[103]),
        .Tile_X6Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[104]),
        .Tile_X6Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[105]),
        .Tile_X6Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[106]),
        .Tile_X6Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[107]),
        .Tile_X6Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[108]),
        .Tile_X6Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[109]),
        .Tile_X6Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[110]),
        .Tile_X6Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[111]),
        .Tile_X6Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[112]),
        .Tile_X6Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[113]),
        .Tile_X6Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[114]),
        .Tile_X6Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[115]),
        .Tile_X6Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[116]),
        .Tile_X6Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[117]),
        .Tile_X6Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[118]),
        .Tile_X6Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[119]),
        .Tile_X7Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[120]),
        .Tile_X7Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[121]),
        .Tile_X7Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[122]),
        .Tile_X7Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[123]),
        .Tile_X7Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[124]),
        .Tile_X7Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[125]),
        .Tile_X7Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[126]),
        .Tile_X7Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[127]),
        .Tile_X7Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[128]),
        .Tile_X7Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[129]),
        .Tile_X7Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[130]),
        .Tile_X7Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[131]),
        .Tile_X7Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[132]),
        .Tile_X7Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[133]),
        .Tile_X7Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[134]),
        .Tile_X7Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[135]),
        .Tile_X7Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[136]),
        .Tile_X7Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[137]),
        .Tile_X7Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[138]),
        .Tile_X7Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[139]),
        .Tile_X8Y7_UIO_BOT_UOUT0(UIO_BOT_UOUT[140]),
        .Tile_X8Y7_UIO_BOT_UOUT1(UIO_BOT_UOUT[141]),
        .Tile_X8Y7_UIO_BOT_UOUT2(UIO_BOT_UOUT[142]),
        .Tile_X8Y7_UIO_BOT_UOUT3(UIO_BOT_UOUT[143]),
        .Tile_X8Y7_UIO_BOT_UOUT4(UIO_BOT_UOUT[144]),
        .Tile_X8Y7_UIO_BOT_UOUT5(UIO_BOT_UOUT[145]),
        .Tile_X8Y7_UIO_BOT_UOUT6(UIO_BOT_UOUT[146]),
        .Tile_X8Y7_UIO_BOT_UOUT7(UIO_BOT_UOUT[147]),
        .Tile_X8Y7_UIO_BOT_UOUT8(UIO_BOT_UOUT[148]),
        .Tile_X8Y7_UIO_BOT_UOUT9(UIO_BOT_UOUT[149]),
        .Tile_X8Y7_UIO_BOT_UOUT10(UIO_BOT_UOUT[150]),
        .Tile_X8Y7_UIO_BOT_UOUT11(UIO_BOT_UOUT[151]),
        .Tile_X8Y7_UIO_BOT_UOUT12(UIO_BOT_UOUT[152]),
        .Tile_X8Y7_UIO_BOT_UOUT13(UIO_BOT_UOUT[153]),
        .Tile_X8Y7_UIO_BOT_UOUT14(UIO_BOT_UOUT[154]),
        .Tile_X8Y7_UIO_BOT_UOUT15(UIO_BOT_UOUT[155]),
        .Tile_X8Y7_UIO_BOT_UOUT16(UIO_BOT_UOUT[156]),
        .Tile_X8Y7_UIO_BOT_UOUT17(UIO_BOT_UOUT[157]),
        .Tile_X8Y7_UIO_BOT_UOUT18(UIO_BOT_UOUT[158]),
        .Tile_X8Y7_UIO_BOT_UOUT19(UIO_BOT_UOUT[159]),
        .Tile_X1Y0_UIO_TOP_UIN0(UIO_TOP_UIN[0]),
        .Tile_X1Y0_UIO_TOP_UIN1(UIO_TOP_UIN[1]),
        .Tile_X1Y0_UIO_TOP_UIN2(UIO_TOP_UIN[2]),
        .Tile_X1Y0_UIO_TOP_UIN3(UIO_TOP_UIN[3]),
        .Tile_X1Y0_UIO_TOP_UIN4(UIO_TOP_UIN[4]),
        .Tile_X1Y0_UIO_TOP_UIN5(UIO_TOP_UIN[5]),
        .Tile_X1Y0_UIO_TOP_UIN6(UIO_TOP_UIN[6]),
        .Tile_X1Y0_UIO_TOP_UIN7(UIO_TOP_UIN[7]),
        .Tile_X1Y0_UIO_TOP_UIN8(UIO_TOP_UIN[8]),
        .Tile_X1Y0_UIO_TOP_UIN9(UIO_TOP_UIN[9]),
        .Tile_X1Y0_UIO_TOP_UIN10(UIO_TOP_UIN[10]),
        .Tile_X1Y0_UIO_TOP_UIN11(UIO_TOP_UIN[11]),
        .Tile_X1Y0_UIO_TOP_UIN12(UIO_TOP_UIN[12]),
        .Tile_X1Y0_UIO_TOP_UIN13(UIO_TOP_UIN[13]),
        .Tile_X1Y0_UIO_TOP_UIN14(UIO_TOP_UIN[14]),
        .Tile_X1Y0_UIO_TOP_UIN15(UIO_TOP_UIN[15]),
        .Tile_X1Y0_UIO_TOP_UIN16(UIO_TOP_UIN[16]),
        .Tile_X1Y0_UIO_TOP_UIN17(UIO_TOP_UIN[17]),
        .Tile_X1Y0_UIO_TOP_UIN18(UIO_TOP_UIN[18]),
        .Tile_X1Y0_UIO_TOP_UIN19(UIO_TOP_UIN[19]),
        .Tile_X2Y0_UIO_TOP_UIN0(UIO_TOP_UIN[20]),
        .Tile_X2Y0_UIO_TOP_UIN1(UIO_TOP_UIN[21]),
        .Tile_X2Y0_UIO_TOP_UIN2(UIO_TOP_UIN[22]),
        .Tile_X2Y0_UIO_TOP_UIN3(UIO_TOP_UIN[23]),
        .Tile_X2Y0_UIO_TOP_UIN4(UIO_TOP_UIN[24]),
        .Tile_X2Y0_UIO_TOP_UIN5(UIO_TOP_UIN[25]),
        .Tile_X2Y0_UIO_TOP_UIN6(UIO_TOP_UIN[26]),
        .Tile_X2Y0_UIO_TOP_UIN7(UIO_TOP_UIN[27]),
        .Tile_X2Y0_UIO_TOP_UIN8(UIO_TOP_UIN[28]),
        .Tile_X2Y0_UIO_TOP_UIN9(UIO_TOP_UIN[29]),
        .Tile_X2Y0_UIO_TOP_UIN10(UIO_TOP_UIN[30]),
        .Tile_X2Y0_UIO_TOP_UIN11(UIO_TOP_UIN[31]),
        .Tile_X2Y0_UIO_TOP_UIN12(UIO_TOP_UIN[32]),
        .Tile_X2Y0_UIO_TOP_UIN13(UIO_TOP_UIN[33]),
        .Tile_X2Y0_UIO_TOP_UIN14(UIO_TOP_UIN[34]),
        .Tile_X2Y0_UIO_TOP_UIN15(UIO_TOP_UIN[35]),
        .Tile_X2Y0_UIO_TOP_UIN16(UIO_TOP_UIN[36]),
        .Tile_X2Y0_UIO_TOP_UIN17(UIO_TOP_UIN[37]),
        .Tile_X2Y0_UIO_TOP_UIN18(UIO_TOP_UIN[38]),
        .Tile_X2Y0_UIO_TOP_UIN19(UIO_TOP_UIN[39]),
        .Tile_X3Y0_UIO_TOP_UIN0(UIO_TOP_UIN[40]),
        .Tile_X3Y0_UIO_TOP_UIN1(UIO_TOP_UIN[41]),
        .Tile_X3Y0_UIO_TOP_UIN2(UIO_TOP_UIN[42]),
        .Tile_X3Y0_UIO_TOP_UIN3(UIO_TOP_UIN[43]),
        .Tile_X3Y0_UIO_TOP_UIN4(UIO_TOP_UIN[44]),
        .Tile_X3Y0_UIO_TOP_UIN5(UIO_TOP_UIN[45]),
        .Tile_X3Y0_UIO_TOP_UIN6(UIO_TOP_UIN[46]),
        .Tile_X3Y0_UIO_TOP_UIN7(UIO_TOP_UIN[47]),
        .Tile_X3Y0_UIO_TOP_UIN8(UIO_TOP_UIN[48]),
        .Tile_X3Y0_UIO_TOP_UIN9(UIO_TOP_UIN[49]),
        .Tile_X3Y0_UIO_TOP_UIN10(UIO_TOP_UIN[50]),
        .Tile_X3Y0_UIO_TOP_UIN11(UIO_TOP_UIN[51]),
        .Tile_X3Y0_UIO_TOP_UIN12(UIO_TOP_UIN[52]),
        .Tile_X3Y0_UIO_TOP_UIN13(UIO_TOP_UIN[53]),
        .Tile_X3Y0_UIO_TOP_UIN14(UIO_TOP_UIN[54]),
        .Tile_X3Y0_UIO_TOP_UIN15(UIO_TOP_UIN[55]),
        .Tile_X3Y0_UIO_TOP_UIN16(UIO_TOP_UIN[56]),
        .Tile_X3Y0_UIO_TOP_UIN17(UIO_TOP_UIN[57]),
        .Tile_X3Y0_UIO_TOP_UIN18(UIO_TOP_UIN[58]),
        .Tile_X3Y0_UIO_TOP_UIN19(UIO_TOP_UIN[59]),
        .Tile_X4Y0_UIO_TOP_UIN0(UIO_TOP_UIN[60]),
        .Tile_X4Y0_UIO_TOP_UIN1(UIO_TOP_UIN[61]),
        .Tile_X4Y0_UIO_TOP_UIN2(UIO_TOP_UIN[62]),
        .Tile_X4Y0_UIO_TOP_UIN3(UIO_TOP_UIN[63]),
        .Tile_X4Y0_UIO_TOP_UIN4(UIO_TOP_UIN[64]),
        .Tile_X4Y0_UIO_TOP_UIN5(UIO_TOP_UIN[65]),
        .Tile_X4Y0_UIO_TOP_UIN6(UIO_TOP_UIN[66]),
        .Tile_X4Y0_UIO_TOP_UIN7(UIO_TOP_UIN[67]),
        .Tile_X4Y0_UIO_TOP_UIN8(UIO_TOP_UIN[68]),
        .Tile_X4Y0_UIO_TOP_UIN9(UIO_TOP_UIN[69]),
        .Tile_X4Y0_UIO_TOP_UIN10(UIO_TOP_UIN[70]),
        .Tile_X4Y0_UIO_TOP_UIN11(UIO_TOP_UIN[71]),
        .Tile_X4Y0_UIO_TOP_UIN12(UIO_TOP_UIN[72]),
        .Tile_X4Y0_UIO_TOP_UIN13(UIO_TOP_UIN[73]),
        .Tile_X4Y0_UIO_TOP_UIN14(UIO_TOP_UIN[74]),
        .Tile_X4Y0_UIO_TOP_UIN15(UIO_TOP_UIN[75]),
        .Tile_X4Y0_UIO_TOP_UIN16(UIO_TOP_UIN[76]),
        .Tile_X4Y0_UIO_TOP_UIN17(UIO_TOP_UIN[77]),
        .Tile_X4Y0_UIO_TOP_UIN18(UIO_TOP_UIN[78]),
        .Tile_X4Y0_UIO_TOP_UIN19(UIO_TOP_UIN[79]),
        .Tile_X5Y0_UIO_TOP_UIN0(UIO_TOP_UIN[80]),
        .Tile_X5Y0_UIO_TOP_UIN1(UIO_TOP_UIN[81]),
        .Tile_X5Y0_UIO_TOP_UIN2(UIO_TOP_UIN[82]),
        .Tile_X5Y0_UIO_TOP_UIN3(UIO_TOP_UIN[83]),
        .Tile_X5Y0_UIO_TOP_UIN4(UIO_TOP_UIN[84]),
        .Tile_X5Y0_UIO_TOP_UIN5(UIO_TOP_UIN[85]),
        .Tile_X5Y0_UIO_TOP_UIN6(UIO_TOP_UIN[86]),
        .Tile_X5Y0_UIO_TOP_UIN7(UIO_TOP_UIN[87]),
        .Tile_X5Y0_UIO_TOP_UIN8(UIO_TOP_UIN[88]),
        .Tile_X5Y0_UIO_TOP_UIN9(UIO_TOP_UIN[89]),
        .Tile_X5Y0_UIO_TOP_UIN10(UIO_TOP_UIN[90]),
        .Tile_X5Y0_UIO_TOP_UIN11(UIO_TOP_UIN[91]),
        .Tile_X5Y0_UIO_TOP_UIN12(UIO_TOP_UIN[92]),
        .Tile_X5Y0_UIO_TOP_UIN13(UIO_TOP_UIN[93]),
        .Tile_X5Y0_UIO_TOP_UIN14(UIO_TOP_UIN[94]),
        .Tile_X5Y0_UIO_TOP_UIN15(UIO_TOP_UIN[95]),
        .Tile_X5Y0_UIO_TOP_UIN16(UIO_TOP_UIN[96]),
        .Tile_X5Y0_UIO_TOP_UIN17(UIO_TOP_UIN[97]),
        .Tile_X5Y0_UIO_TOP_UIN18(UIO_TOP_UIN[98]),
        .Tile_X5Y0_UIO_TOP_UIN19(UIO_TOP_UIN[99]),
        .Tile_X6Y0_UIO_TOP_UIN0(UIO_TOP_UIN[100]),
        .Tile_X6Y0_UIO_TOP_UIN1(UIO_TOP_UIN[101]),
        .Tile_X6Y0_UIO_TOP_UIN2(UIO_TOP_UIN[102]),
        .Tile_X6Y0_UIO_TOP_UIN3(UIO_TOP_UIN[103]),
        .Tile_X6Y0_UIO_TOP_UIN4(UIO_TOP_UIN[104]),
        .Tile_X6Y0_UIO_TOP_UIN5(UIO_TOP_UIN[105]),
        .Tile_X6Y0_UIO_TOP_UIN6(UIO_TOP_UIN[106]),
        .Tile_X6Y0_UIO_TOP_UIN7(UIO_TOP_UIN[107]),
        .Tile_X6Y0_UIO_TOP_UIN8(UIO_TOP_UIN[108]),
        .Tile_X6Y0_UIO_TOP_UIN9(UIO_TOP_UIN[109]),
        .Tile_X6Y0_UIO_TOP_UIN10(UIO_TOP_UIN[110]),
        .Tile_X6Y0_UIO_TOP_UIN11(UIO_TOP_UIN[111]),
        .Tile_X6Y0_UIO_TOP_UIN12(UIO_TOP_UIN[112]),
        .Tile_X6Y0_UIO_TOP_UIN13(UIO_TOP_UIN[113]),
        .Tile_X6Y0_UIO_TOP_UIN14(UIO_TOP_UIN[114]),
        .Tile_X6Y0_UIO_TOP_UIN15(UIO_TOP_UIN[115]),
        .Tile_X6Y0_UIO_TOP_UIN16(UIO_TOP_UIN[116]),
        .Tile_X6Y0_UIO_TOP_UIN17(UIO_TOP_UIN[117]),
        .Tile_X6Y0_UIO_TOP_UIN18(UIO_TOP_UIN[118]),
        .Tile_X6Y0_UIO_TOP_UIN19(UIO_TOP_UIN[119]),
        .Tile_X7Y0_UIO_TOP_UIN0(UIO_TOP_UIN[120]),
        .Tile_X7Y0_UIO_TOP_UIN1(UIO_TOP_UIN[121]),
        .Tile_X7Y0_UIO_TOP_UIN2(UIO_TOP_UIN[122]),
        .Tile_X7Y0_UIO_TOP_UIN3(UIO_TOP_UIN[123]),
        .Tile_X7Y0_UIO_TOP_UIN4(UIO_TOP_UIN[124]),
        .Tile_X7Y0_UIO_TOP_UIN5(UIO_TOP_UIN[125]),
        .Tile_X7Y0_UIO_TOP_UIN6(UIO_TOP_UIN[126]),
        .Tile_X7Y0_UIO_TOP_UIN7(UIO_TOP_UIN[127]),
        .Tile_X7Y0_UIO_TOP_UIN8(UIO_TOP_UIN[128]),
        .Tile_X7Y0_UIO_TOP_UIN9(UIO_TOP_UIN[129]),
        .Tile_X7Y0_UIO_TOP_UIN10(UIO_TOP_UIN[130]),
        .Tile_X7Y0_UIO_TOP_UIN11(UIO_TOP_UIN[131]),
        .Tile_X7Y0_UIO_TOP_UIN12(UIO_TOP_UIN[132]),
        .Tile_X7Y0_UIO_TOP_UIN13(UIO_TOP_UIN[133]),
        .Tile_X7Y0_UIO_TOP_UIN14(UIO_TOP_UIN[134]),
        .Tile_X7Y0_UIO_TOP_UIN15(UIO_TOP_UIN[135]),
        .Tile_X7Y0_UIO_TOP_UIN16(UIO_TOP_UIN[136]),
        .Tile_X7Y0_UIO_TOP_UIN17(UIO_TOP_UIN[137]),
        .Tile_X7Y0_UIO_TOP_UIN18(UIO_TOP_UIN[138]),
        .Tile_X7Y0_UIO_TOP_UIN19(UIO_TOP_UIN[139]),
        .Tile_X8Y0_UIO_TOP_UIN0(UIO_TOP_UIN[140]),
        .Tile_X8Y0_UIO_TOP_UIN1(UIO_TOP_UIN[141]),
        .Tile_X8Y0_UIO_TOP_UIN2(UIO_TOP_UIN[142]),
        .Tile_X8Y0_UIO_TOP_UIN3(UIO_TOP_UIN[143]),
        .Tile_X8Y0_UIO_TOP_UIN4(UIO_TOP_UIN[144]),
        .Tile_X8Y0_UIO_TOP_UIN5(UIO_TOP_UIN[145]),
        .Tile_X8Y0_UIO_TOP_UIN6(UIO_TOP_UIN[146]),
        .Tile_X8Y0_UIO_TOP_UIN7(UIO_TOP_UIN[147]),
        .Tile_X8Y0_UIO_TOP_UIN8(UIO_TOP_UIN[148]),
        .Tile_X8Y0_UIO_TOP_UIN9(UIO_TOP_UIN[149]),
        .Tile_X8Y0_UIO_TOP_UIN10(UIO_TOP_UIN[150]),
        .Tile_X8Y0_UIO_TOP_UIN11(UIO_TOP_UIN[151]),
        .Tile_X8Y0_UIO_TOP_UIN12(UIO_TOP_UIN[152]),
        .Tile_X8Y0_UIO_TOP_UIN13(UIO_TOP_UIN[153]),
        .Tile_X8Y0_UIO_TOP_UIN14(UIO_TOP_UIN[154]),
        .Tile_X8Y0_UIO_TOP_UIN15(UIO_TOP_UIN[155]),
        .Tile_X8Y0_UIO_TOP_UIN16(UIO_TOP_UIN[156]),
        .Tile_X8Y0_UIO_TOP_UIN17(UIO_TOP_UIN[157]),
        .Tile_X8Y0_UIO_TOP_UIN18(UIO_TOP_UIN[158]),
        .Tile_X8Y0_UIO_TOP_UIN19(UIO_TOP_UIN[159]),
        .Tile_X1Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[0]),
        .Tile_X1Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[1]),
        .Tile_X1Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[2]),
        .Tile_X1Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[3]),
        .Tile_X1Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[4]),
        .Tile_X1Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[5]),
        .Tile_X1Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[6]),
        .Tile_X1Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[7]),
        .Tile_X1Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[8]),
        .Tile_X1Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[9]),
        .Tile_X1Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[10]),
        .Tile_X1Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[11]),
        .Tile_X1Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[12]),
        .Tile_X1Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[13]),
        .Tile_X1Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[14]),
        .Tile_X1Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[15]),
        .Tile_X1Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[16]),
        .Tile_X1Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[17]),
        .Tile_X1Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[18]),
        .Tile_X1Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[19]),
        .Tile_X2Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[20]),
        .Tile_X2Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[21]),
        .Tile_X2Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[22]),
        .Tile_X2Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[23]),
        .Tile_X2Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[24]),
        .Tile_X2Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[25]),
        .Tile_X2Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[26]),
        .Tile_X2Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[27]),
        .Tile_X2Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[28]),
        .Tile_X2Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[29]),
        .Tile_X2Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[30]),
        .Tile_X2Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[31]),
        .Tile_X2Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[32]),
        .Tile_X2Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[33]),
        .Tile_X2Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[34]),
        .Tile_X2Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[35]),
        .Tile_X2Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[36]),
        .Tile_X2Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[37]),
        .Tile_X2Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[38]),
        .Tile_X2Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[39]),
        .Tile_X3Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[40]),
        .Tile_X3Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[41]),
        .Tile_X3Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[42]),
        .Tile_X3Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[43]),
        .Tile_X3Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[44]),
        .Tile_X3Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[45]),
        .Tile_X3Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[46]),
        .Tile_X3Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[47]),
        .Tile_X3Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[48]),
        .Tile_X3Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[49]),
        .Tile_X3Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[50]),
        .Tile_X3Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[51]),
        .Tile_X3Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[52]),
        .Tile_X3Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[53]),
        .Tile_X3Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[54]),
        .Tile_X3Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[55]),
        .Tile_X3Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[56]),
        .Tile_X3Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[57]),
        .Tile_X3Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[58]),
        .Tile_X3Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[59]),
        .Tile_X4Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[60]),
        .Tile_X4Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[61]),
        .Tile_X4Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[62]),
        .Tile_X4Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[63]),
        .Tile_X4Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[64]),
        .Tile_X4Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[65]),
        .Tile_X4Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[66]),
        .Tile_X4Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[67]),
        .Tile_X4Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[68]),
        .Tile_X4Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[69]),
        .Tile_X4Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[70]),
        .Tile_X4Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[71]),
        .Tile_X4Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[72]),
        .Tile_X4Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[73]),
        .Tile_X4Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[74]),
        .Tile_X4Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[75]),
        .Tile_X4Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[76]),
        .Tile_X4Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[77]),
        .Tile_X4Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[78]),
        .Tile_X4Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[79]),
        .Tile_X5Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[80]),
        .Tile_X5Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[81]),
        .Tile_X5Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[82]),
        .Tile_X5Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[83]),
        .Tile_X5Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[84]),
        .Tile_X5Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[85]),
        .Tile_X5Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[86]),
        .Tile_X5Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[87]),
        .Tile_X5Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[88]),
        .Tile_X5Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[89]),
        .Tile_X5Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[90]),
        .Tile_X5Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[91]),
        .Tile_X5Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[92]),
        .Tile_X5Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[93]),
        .Tile_X5Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[94]),
        .Tile_X5Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[95]),
        .Tile_X5Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[96]),
        .Tile_X5Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[97]),
        .Tile_X5Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[98]),
        .Tile_X5Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[99]),
        .Tile_X6Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[100]),
        .Tile_X6Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[101]),
        .Tile_X6Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[102]),
        .Tile_X6Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[103]),
        .Tile_X6Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[104]),
        .Tile_X6Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[105]),
        .Tile_X6Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[106]),
        .Tile_X6Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[107]),
        .Tile_X6Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[108]),
        .Tile_X6Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[109]),
        .Tile_X6Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[110]),
        .Tile_X6Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[111]),
        .Tile_X6Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[112]),
        .Tile_X6Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[113]),
        .Tile_X6Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[114]),
        .Tile_X6Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[115]),
        .Tile_X6Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[116]),
        .Tile_X6Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[117]),
        .Tile_X6Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[118]),
        .Tile_X6Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[119]),
        .Tile_X7Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[120]),
        .Tile_X7Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[121]),
        .Tile_X7Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[122]),
        .Tile_X7Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[123]),
        .Tile_X7Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[124]),
        .Tile_X7Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[125]),
        .Tile_X7Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[126]),
        .Tile_X7Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[127]),
        .Tile_X7Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[128]),
        .Tile_X7Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[129]),
        .Tile_X7Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[130]),
        .Tile_X7Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[131]),
        .Tile_X7Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[132]),
        .Tile_X7Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[133]),
        .Tile_X7Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[134]),
        .Tile_X7Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[135]),
        .Tile_X7Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[136]),
        .Tile_X7Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[137]),
        .Tile_X7Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[138]),
        .Tile_X7Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[139]),
        .Tile_X8Y0_UIO_TOP_UOUT0(UIO_TOP_UOUT[140]),
        .Tile_X8Y0_UIO_TOP_UOUT1(UIO_TOP_UOUT[141]),
        .Tile_X8Y0_UIO_TOP_UOUT2(UIO_TOP_UOUT[142]),
        .Tile_X8Y0_UIO_TOP_UOUT3(UIO_TOP_UOUT[143]),
        .Tile_X8Y0_UIO_TOP_UOUT4(UIO_TOP_UOUT[144]),
        .Tile_X8Y0_UIO_TOP_UOUT5(UIO_TOP_UOUT[145]),
        .Tile_X8Y0_UIO_TOP_UOUT6(UIO_TOP_UOUT[146]),
        .Tile_X8Y0_UIO_TOP_UOUT7(UIO_TOP_UOUT[147]),
        .Tile_X8Y0_UIO_TOP_UOUT8(UIO_TOP_UOUT[148]),
        .Tile_X8Y0_UIO_TOP_UOUT9(UIO_TOP_UOUT[149]),
        .Tile_X8Y0_UIO_TOP_UOUT10(UIO_TOP_UOUT[150]),
        .Tile_X8Y0_UIO_TOP_UOUT11(UIO_TOP_UOUT[151]),
        .Tile_X8Y0_UIO_TOP_UOUT12(UIO_TOP_UOUT[152]),
        .Tile_X8Y0_UIO_TOP_UOUT13(UIO_TOP_UOUT[153]),
        .Tile_X8Y0_UIO_TOP_UOUT14(UIO_TOP_UOUT[154]),
        .Tile_X8Y0_UIO_TOP_UOUT15(UIO_TOP_UOUT[155]),
        .Tile_X8Y0_UIO_TOP_UOUT16(UIO_TOP_UOUT[156]),
        .Tile_X8Y0_UIO_TOP_UOUT17(UIO_TOP_UOUT[157]),
        .Tile_X8Y0_UIO_TOP_UOUT18(UIO_TOP_UOUT[158]),
        .Tile_X8Y0_UIO_TOP_UOUT19(UIO_TOP_UOUT[159]),
        .UserCLK(CLK),
        .FrameData(FrameData),
        .FrameStrobe(FrameSelect)
    );


    BlockRAM_1KB Inst_BlockRAM_0 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .clk(CLK),
        .rd_addr(FAB2RAM_A_O[7:0]),
        .rd_data(RAM2FAB_D_I[31:0]),
        .wr_addr(FAB2RAM_A_O[15:8]),
        .wr_data(FAB2RAM_D_O[31:0]),
        .C0(FAB2RAM_C_O[0]),
        .C1(FAB2RAM_C_O[1]),
        .C2(FAB2RAM_C_O[2]),
        .C3(FAB2RAM_C_O[3]),
        .C4(FAB2RAM_C_O[4]),
        .C5(FAB2RAM_C_O[5])
    );

    BlockRAM_1KB Inst_BlockRAM_1 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .clk(CLK),
        .rd_addr(FAB2RAM_A_O[23:16]),
        .rd_data(RAM2FAB_D_I[63:32]),
        .wr_addr(FAB2RAM_A_O[31:24]),
        .wr_data(FAB2RAM_D_O[63:32]),
        .C0(FAB2RAM_C_O[8]),
        .C1(FAB2RAM_C_O[9]),
        .C2(FAB2RAM_C_O[10]),
        .C3(FAB2RAM_C_O[11]),
        .C4(FAB2RAM_C_O[12]),
        .C5(FAB2RAM_C_O[13])
    );

    BlockRAM_1KB Inst_BlockRAM_2 (
`ifdef USE_POWER_PINS
        .vccd1(vccd1),
        .vssd1(vssd1),
`endif
        .clk(CLK),
        .rd_addr(FAB2RAM_A_O[39:32]),
        .rd_data(RAM2FAB_D_I[95:64]),
        .wr_addr(FAB2RAM_A_O[47:40]),
        .wr_data(FAB2RAM_D_O[95:64]),
        .C0(FAB2RAM_C_O[16]),
        .C1(FAB2RAM_C_O[17]),
        .C2(FAB2RAM_C_O[18]),
        .C3(FAB2RAM_C_O[19]),
        .C4(FAB2RAM_C_O[20]),
        .C5(FAB2RAM_C_O[21])
    );

    assign FrameData = {32'h12345678, FrameRegister, 32'h12345678};
endmodule
/* verilator lint_on UNUSEDSIGNAL */

