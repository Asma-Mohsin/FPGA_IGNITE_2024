magic
tech sky130A
magscale 1 2
timestamp 1732405368
<< obsli1 >>
rect 1104 2159 44896 5457
<< obsm1 >>
rect 842 1164 45051 6588
<< metal2 >>
rect 5722 7840 5778 8000
rect 5998 7840 6054 8000
rect 6274 7840 6330 8000
rect 6550 7840 6606 8000
rect 6826 7840 6882 8000
rect 7102 7840 7158 8000
rect 7378 7840 7434 8000
rect 7654 7840 7710 8000
rect 7930 7840 7986 8000
rect 8206 7840 8262 8000
rect 8482 7840 8538 8000
rect 8758 7840 8814 8000
rect 9034 7840 9090 8000
rect 9310 7840 9366 8000
rect 9586 7840 9642 8000
rect 9862 7840 9918 8000
rect 10138 7840 10194 8000
rect 10414 7840 10470 8000
rect 10690 7840 10746 8000
rect 10966 7840 11022 8000
rect 11242 7840 11298 8000
rect 11518 7840 11574 8000
rect 11794 7840 11850 8000
rect 12070 7840 12126 8000
rect 12346 7840 12402 8000
rect 12622 7840 12678 8000
rect 12898 7840 12954 8000
rect 13174 7840 13230 8000
rect 13450 7840 13506 8000
rect 13726 7840 13782 8000
rect 14002 7840 14058 8000
rect 14278 7840 14334 8000
rect 14554 7840 14610 8000
rect 14830 7840 14886 8000
rect 15106 7840 15162 8000
rect 15382 7840 15438 8000
rect 15658 7840 15714 8000
rect 15934 7840 15990 8000
rect 16210 7840 16266 8000
rect 16486 7840 16542 8000
rect 16762 7840 16818 8000
rect 17038 7840 17094 8000
rect 17314 7840 17370 8000
rect 17590 7840 17646 8000
rect 17866 7840 17922 8000
rect 18142 7840 18198 8000
rect 18418 7840 18474 8000
rect 18694 7840 18750 8000
rect 18970 7840 19026 8000
rect 19246 7840 19302 8000
rect 19522 7840 19578 8000
rect 19798 7840 19854 8000
rect 20074 7840 20130 8000
rect 20350 7840 20406 8000
rect 20626 7840 20682 8000
rect 20902 7840 20958 8000
rect 21178 7840 21234 8000
rect 21454 7840 21510 8000
rect 21730 7840 21786 8000
rect 22006 7840 22062 8000
rect 22282 7840 22338 8000
rect 22558 7840 22614 8000
rect 22834 7840 22890 8000
rect 23110 7840 23166 8000
rect 23386 7840 23442 8000
rect 23662 7840 23718 8000
rect 23938 7840 23994 8000
rect 24214 7840 24270 8000
rect 24490 7840 24546 8000
rect 24766 7840 24822 8000
rect 25042 7840 25098 8000
rect 25318 7840 25374 8000
rect 25594 7840 25650 8000
rect 25870 7840 25926 8000
rect 26146 7840 26202 8000
rect 26422 7840 26478 8000
rect 26698 7840 26754 8000
rect 26974 7840 27030 8000
rect 27250 7840 27306 8000
rect 27526 7840 27582 8000
rect 27802 7840 27858 8000
rect 28078 7840 28134 8000
rect 28354 7840 28410 8000
rect 28630 7840 28686 8000
rect 28906 7840 28962 8000
rect 29182 7840 29238 8000
rect 29458 7840 29514 8000
rect 29734 7840 29790 8000
rect 30010 7840 30066 8000
rect 30286 7840 30342 8000
rect 30562 7840 30618 8000
rect 30838 7840 30894 8000
rect 31114 7840 31170 8000
rect 31390 7840 31446 8000
rect 31666 7840 31722 8000
rect 31942 7840 31998 8000
rect 32218 7840 32274 8000
rect 32494 7840 32550 8000
rect 32770 7840 32826 8000
rect 33046 7840 33102 8000
rect 33322 7840 33378 8000
rect 33598 7840 33654 8000
rect 33874 7840 33930 8000
rect 34150 7840 34206 8000
rect 34426 7840 34482 8000
rect 34702 7840 34758 8000
rect 34978 7840 35034 8000
rect 35254 7840 35310 8000
rect 35530 7840 35586 8000
rect 35806 7840 35862 8000
rect 36082 7840 36138 8000
rect 36358 7840 36414 8000
rect 36634 7840 36690 8000
rect 36910 7840 36966 8000
rect 37186 7840 37242 8000
rect 37462 7840 37518 8000
rect 37738 7840 37794 8000
rect 38014 7840 38070 8000
rect 38290 7840 38346 8000
rect 38566 7840 38622 8000
rect 38842 7840 38898 8000
rect 39118 7840 39174 8000
rect 39394 7840 39450 8000
rect 39670 7840 39726 8000
rect 39946 7840 40002 8000
rect 40222 7840 40278 8000
rect 846 0 902 160
rect 1582 0 1638 160
rect 2318 0 2374 160
rect 3054 0 3110 160
rect 3790 0 3846 160
rect 4526 0 4582 160
rect 5262 0 5318 160
rect 5998 0 6054 160
rect 6734 0 6790 160
rect 7470 0 7526 160
rect 8206 0 8262 160
rect 8942 0 8998 160
rect 9678 0 9734 160
rect 10414 0 10470 160
rect 11150 0 11206 160
rect 11886 0 11942 160
rect 12622 0 12678 160
rect 13358 0 13414 160
rect 14094 0 14150 160
rect 14830 0 14886 160
rect 15566 0 15622 160
rect 16302 0 16358 160
rect 17038 0 17094 160
rect 17774 0 17830 160
rect 18510 0 18566 160
rect 19246 0 19302 160
rect 19982 0 20038 160
rect 20718 0 20774 160
rect 21454 0 21510 160
rect 22190 0 22246 160
rect 22926 0 22982 160
rect 23662 0 23718 160
rect 24398 0 24454 160
rect 25134 0 25190 160
rect 25870 0 25926 160
rect 26606 0 26662 160
rect 27342 0 27398 160
rect 28078 0 28134 160
rect 28814 0 28870 160
rect 29550 0 29606 160
rect 30286 0 30342 160
rect 31022 0 31078 160
rect 31758 0 31814 160
rect 32494 0 32550 160
rect 33230 0 33286 160
rect 33966 0 34022 160
rect 34702 0 34758 160
rect 35438 0 35494 160
rect 36174 0 36230 160
rect 36910 0 36966 160
rect 37646 0 37702 160
rect 38382 0 38438 160
rect 39118 0 39174 160
rect 39854 0 39910 160
rect 40590 0 40646 160
rect 41326 0 41382 160
rect 42062 0 42118 160
rect 42798 0 42854 160
rect 43534 0 43590 160
rect 44270 0 44326 160
rect 45006 0 45062 160
<< obsm2 >>
rect 848 7784 5666 7970
rect 5834 7784 5942 7970
rect 6110 7784 6218 7970
rect 6386 7784 6494 7970
rect 6662 7784 6770 7970
rect 6938 7784 7046 7970
rect 7214 7784 7322 7970
rect 7490 7784 7598 7970
rect 7766 7784 7874 7970
rect 8042 7784 8150 7970
rect 8318 7784 8426 7970
rect 8594 7784 8702 7970
rect 8870 7784 8978 7970
rect 9146 7784 9254 7970
rect 9422 7784 9530 7970
rect 9698 7784 9806 7970
rect 9974 7784 10082 7970
rect 10250 7784 10358 7970
rect 10526 7784 10634 7970
rect 10802 7784 10910 7970
rect 11078 7784 11186 7970
rect 11354 7784 11462 7970
rect 11630 7784 11738 7970
rect 11906 7784 12014 7970
rect 12182 7784 12290 7970
rect 12458 7784 12566 7970
rect 12734 7784 12842 7970
rect 13010 7784 13118 7970
rect 13286 7784 13394 7970
rect 13562 7784 13670 7970
rect 13838 7784 13946 7970
rect 14114 7784 14222 7970
rect 14390 7784 14498 7970
rect 14666 7784 14774 7970
rect 14942 7784 15050 7970
rect 15218 7784 15326 7970
rect 15494 7784 15602 7970
rect 15770 7784 15878 7970
rect 16046 7784 16154 7970
rect 16322 7784 16430 7970
rect 16598 7784 16706 7970
rect 16874 7784 16982 7970
rect 17150 7784 17258 7970
rect 17426 7784 17534 7970
rect 17702 7784 17810 7970
rect 17978 7784 18086 7970
rect 18254 7784 18362 7970
rect 18530 7784 18638 7970
rect 18806 7784 18914 7970
rect 19082 7784 19190 7970
rect 19358 7784 19466 7970
rect 19634 7784 19742 7970
rect 19910 7784 20018 7970
rect 20186 7784 20294 7970
rect 20462 7784 20570 7970
rect 20738 7784 20846 7970
rect 21014 7784 21122 7970
rect 21290 7784 21398 7970
rect 21566 7784 21674 7970
rect 21842 7784 21950 7970
rect 22118 7784 22226 7970
rect 22394 7784 22502 7970
rect 22670 7784 22778 7970
rect 22946 7784 23054 7970
rect 23222 7784 23330 7970
rect 23498 7784 23606 7970
rect 23774 7784 23882 7970
rect 24050 7784 24158 7970
rect 24326 7784 24434 7970
rect 24602 7784 24710 7970
rect 24878 7784 24986 7970
rect 25154 7784 25262 7970
rect 25430 7784 25538 7970
rect 25706 7784 25814 7970
rect 25982 7784 26090 7970
rect 26258 7784 26366 7970
rect 26534 7784 26642 7970
rect 26810 7784 26918 7970
rect 27086 7784 27194 7970
rect 27362 7784 27470 7970
rect 27638 7784 27746 7970
rect 27914 7784 28022 7970
rect 28190 7784 28298 7970
rect 28466 7784 28574 7970
rect 28742 7784 28850 7970
rect 29018 7784 29126 7970
rect 29294 7784 29402 7970
rect 29570 7784 29678 7970
rect 29846 7784 29954 7970
rect 30122 7784 30230 7970
rect 30398 7784 30506 7970
rect 30674 7784 30782 7970
rect 30950 7784 31058 7970
rect 31226 7784 31334 7970
rect 31502 7784 31610 7970
rect 31778 7784 31886 7970
rect 32054 7784 32162 7970
rect 32330 7784 32438 7970
rect 32606 7784 32714 7970
rect 32882 7784 32990 7970
rect 33158 7784 33266 7970
rect 33434 7784 33542 7970
rect 33710 7784 33818 7970
rect 33986 7784 34094 7970
rect 34262 7784 34370 7970
rect 34538 7784 34646 7970
rect 34814 7784 34922 7970
rect 35090 7784 35198 7970
rect 35366 7784 35474 7970
rect 35642 7784 35750 7970
rect 35918 7784 36026 7970
rect 36194 7784 36302 7970
rect 36470 7784 36578 7970
rect 36746 7784 36854 7970
rect 37022 7784 37130 7970
rect 37298 7784 37406 7970
rect 37574 7784 37682 7970
rect 37850 7784 37958 7970
rect 38126 7784 38234 7970
rect 38402 7784 38510 7970
rect 38678 7784 38786 7970
rect 38954 7784 39062 7970
rect 39230 7784 39338 7970
rect 39506 7784 39614 7970
rect 39782 7784 39890 7970
rect 40058 7784 40166 7970
rect 40334 7784 45045 7970
rect 848 216 45045 7784
rect 958 54 1526 216
rect 1694 54 2262 216
rect 2430 54 2998 216
rect 3166 54 3734 216
rect 3902 54 4470 216
rect 4638 54 5206 216
rect 5374 54 5942 216
rect 6110 54 6678 216
rect 6846 54 7414 216
rect 7582 54 8150 216
rect 8318 54 8886 216
rect 9054 54 9622 216
rect 9790 54 10358 216
rect 10526 54 11094 216
rect 11262 54 11830 216
rect 11998 54 12566 216
rect 12734 54 13302 216
rect 13470 54 14038 216
rect 14206 54 14774 216
rect 14942 54 15510 216
rect 15678 54 16246 216
rect 16414 54 16982 216
rect 17150 54 17718 216
rect 17886 54 18454 216
rect 18622 54 19190 216
rect 19358 54 19926 216
rect 20094 54 20662 216
rect 20830 54 21398 216
rect 21566 54 22134 216
rect 22302 54 22870 216
rect 23038 54 23606 216
rect 23774 54 24342 216
rect 24510 54 25078 216
rect 25246 54 25814 216
rect 25982 54 26550 216
rect 26718 54 27286 216
rect 27454 54 28022 216
rect 28190 54 28758 216
rect 28926 54 29494 216
rect 29662 54 30230 216
rect 30398 54 30966 216
rect 31134 54 31702 216
rect 31870 54 32438 216
rect 32606 54 33174 216
rect 33342 54 33910 216
rect 34078 54 34646 216
rect 34814 54 35382 216
rect 35550 54 36118 216
rect 36286 54 36854 216
rect 37022 54 37590 216
rect 37758 54 38326 216
rect 38494 54 39062 216
rect 39230 54 39798 216
rect 39966 54 40534 216
rect 40702 54 41270 216
rect 41438 54 42006 216
rect 42174 54 42742 216
rect 42910 54 43478 216
rect 43646 54 44214 216
rect 44382 54 44950 216
<< obsm3 >>
rect 4705 1667 45049 5813
<< metal4 >>
rect 6417 2128 6737 5488
rect 11890 2128 12210 5488
rect 17364 2128 17684 5488
rect 22837 2128 23157 5488
rect 28311 2128 28631 5488
rect 33784 2128 34104 5488
rect 39258 2128 39578 5488
rect 44731 2128 45051 5488
<< obsm4 >>
rect 37227 3843 37293 4317
<< labels >>
rlabel metal2 s 34702 7840 34758 8000 6 Co
port 1 nsew signal output
rlabel metal2 s 1582 0 1638 160 6 FrameStrobe[0]
port 2 nsew signal input
rlabel metal2 s 8942 0 8998 160 6 FrameStrobe[10]
port 3 nsew signal input
rlabel metal2 s 9678 0 9734 160 6 FrameStrobe[11]
port 4 nsew signal input
rlabel metal2 s 10414 0 10470 160 6 FrameStrobe[12]
port 5 nsew signal input
rlabel metal2 s 11150 0 11206 160 6 FrameStrobe[13]
port 6 nsew signal input
rlabel metal2 s 11886 0 11942 160 6 FrameStrobe[14]
port 7 nsew signal input
rlabel metal2 s 12622 0 12678 160 6 FrameStrobe[15]
port 8 nsew signal input
rlabel metal2 s 13358 0 13414 160 6 FrameStrobe[16]
port 9 nsew signal input
rlabel metal2 s 14094 0 14150 160 6 FrameStrobe[17]
port 10 nsew signal input
rlabel metal2 s 14830 0 14886 160 6 FrameStrobe[18]
port 11 nsew signal input
rlabel metal2 s 15566 0 15622 160 6 FrameStrobe[19]
port 12 nsew signal input
rlabel metal2 s 2318 0 2374 160 6 FrameStrobe[1]
port 13 nsew signal input
rlabel metal2 s 3054 0 3110 160 6 FrameStrobe[2]
port 14 nsew signal input
rlabel metal2 s 3790 0 3846 160 6 FrameStrobe[3]
port 15 nsew signal input
rlabel metal2 s 4526 0 4582 160 6 FrameStrobe[4]
port 16 nsew signal input
rlabel metal2 s 5262 0 5318 160 6 FrameStrobe[5]
port 17 nsew signal input
rlabel metal2 s 5998 0 6054 160 6 FrameStrobe[6]
port 18 nsew signal input
rlabel metal2 s 6734 0 6790 160 6 FrameStrobe[7]
port 19 nsew signal input
rlabel metal2 s 7470 0 7526 160 6 FrameStrobe[8]
port 20 nsew signal input
rlabel metal2 s 8206 0 8262 160 6 FrameStrobe[9]
port 21 nsew signal input
rlabel metal2 s 34978 7840 35034 8000 6 FrameStrobe_O[0]
port 22 nsew signal output
rlabel metal2 s 37738 7840 37794 8000 6 FrameStrobe_O[10]
port 23 nsew signal output
rlabel metal2 s 38014 7840 38070 8000 6 FrameStrobe_O[11]
port 24 nsew signal output
rlabel metal2 s 38290 7840 38346 8000 6 FrameStrobe_O[12]
port 25 nsew signal output
rlabel metal2 s 38566 7840 38622 8000 6 FrameStrobe_O[13]
port 26 nsew signal output
rlabel metal2 s 38842 7840 38898 8000 6 FrameStrobe_O[14]
port 27 nsew signal output
rlabel metal2 s 39118 7840 39174 8000 6 FrameStrobe_O[15]
port 28 nsew signal output
rlabel metal2 s 39394 7840 39450 8000 6 FrameStrobe_O[16]
port 29 nsew signal output
rlabel metal2 s 39670 7840 39726 8000 6 FrameStrobe_O[17]
port 30 nsew signal output
rlabel metal2 s 39946 7840 40002 8000 6 FrameStrobe_O[18]
port 31 nsew signal output
rlabel metal2 s 40222 7840 40278 8000 6 FrameStrobe_O[19]
port 32 nsew signal output
rlabel metal2 s 35254 7840 35310 8000 6 FrameStrobe_O[1]
port 33 nsew signal output
rlabel metal2 s 35530 7840 35586 8000 6 FrameStrobe_O[2]
port 34 nsew signal output
rlabel metal2 s 35806 7840 35862 8000 6 FrameStrobe_O[3]
port 35 nsew signal output
rlabel metal2 s 36082 7840 36138 8000 6 FrameStrobe_O[4]
port 36 nsew signal output
rlabel metal2 s 36358 7840 36414 8000 6 FrameStrobe_O[5]
port 37 nsew signal output
rlabel metal2 s 36634 7840 36690 8000 6 FrameStrobe_O[6]
port 38 nsew signal output
rlabel metal2 s 36910 7840 36966 8000 6 FrameStrobe_O[7]
port 39 nsew signal output
rlabel metal2 s 37186 7840 37242 8000 6 FrameStrobe_O[8]
port 40 nsew signal output
rlabel metal2 s 37462 7840 37518 8000 6 FrameStrobe_O[9]
port 41 nsew signal output
rlabel metal2 s 5722 7840 5778 8000 6 N1BEG[0]
port 42 nsew signal output
rlabel metal2 s 5998 7840 6054 8000 6 N1BEG[1]
port 43 nsew signal output
rlabel metal2 s 6274 7840 6330 8000 6 N1BEG[2]
port 44 nsew signal output
rlabel metal2 s 6550 7840 6606 8000 6 N1BEG[3]
port 45 nsew signal output
rlabel metal2 s 6826 7840 6882 8000 6 N2BEG[0]
port 46 nsew signal output
rlabel metal2 s 7102 7840 7158 8000 6 N2BEG[1]
port 47 nsew signal output
rlabel metal2 s 7378 7840 7434 8000 6 N2BEG[2]
port 48 nsew signal output
rlabel metal2 s 7654 7840 7710 8000 6 N2BEG[3]
port 49 nsew signal output
rlabel metal2 s 7930 7840 7986 8000 6 N2BEG[4]
port 50 nsew signal output
rlabel metal2 s 8206 7840 8262 8000 6 N2BEG[5]
port 51 nsew signal output
rlabel metal2 s 8482 7840 8538 8000 6 N2BEG[6]
port 52 nsew signal output
rlabel metal2 s 8758 7840 8814 8000 6 N2BEG[7]
port 53 nsew signal output
rlabel metal2 s 9034 7840 9090 8000 6 N2BEGb[0]
port 54 nsew signal output
rlabel metal2 s 9310 7840 9366 8000 6 N2BEGb[1]
port 55 nsew signal output
rlabel metal2 s 9586 7840 9642 8000 6 N2BEGb[2]
port 56 nsew signal output
rlabel metal2 s 9862 7840 9918 8000 6 N2BEGb[3]
port 57 nsew signal output
rlabel metal2 s 10138 7840 10194 8000 6 N2BEGb[4]
port 58 nsew signal output
rlabel metal2 s 10414 7840 10470 8000 6 N2BEGb[5]
port 59 nsew signal output
rlabel metal2 s 10690 7840 10746 8000 6 N2BEGb[6]
port 60 nsew signal output
rlabel metal2 s 10966 7840 11022 8000 6 N2BEGb[7]
port 61 nsew signal output
rlabel metal2 s 11242 7840 11298 8000 6 N4BEG[0]
port 62 nsew signal output
rlabel metal2 s 14002 7840 14058 8000 6 N4BEG[10]
port 63 nsew signal output
rlabel metal2 s 14278 7840 14334 8000 6 N4BEG[11]
port 64 nsew signal output
rlabel metal2 s 14554 7840 14610 8000 6 N4BEG[12]
port 65 nsew signal output
rlabel metal2 s 14830 7840 14886 8000 6 N4BEG[13]
port 66 nsew signal output
rlabel metal2 s 15106 7840 15162 8000 6 N4BEG[14]
port 67 nsew signal output
rlabel metal2 s 15382 7840 15438 8000 6 N4BEG[15]
port 68 nsew signal output
rlabel metal2 s 11518 7840 11574 8000 6 N4BEG[1]
port 69 nsew signal output
rlabel metal2 s 11794 7840 11850 8000 6 N4BEG[2]
port 70 nsew signal output
rlabel metal2 s 12070 7840 12126 8000 6 N4BEG[3]
port 71 nsew signal output
rlabel metal2 s 12346 7840 12402 8000 6 N4BEG[4]
port 72 nsew signal output
rlabel metal2 s 12622 7840 12678 8000 6 N4BEG[5]
port 73 nsew signal output
rlabel metal2 s 12898 7840 12954 8000 6 N4BEG[6]
port 74 nsew signal output
rlabel metal2 s 13174 7840 13230 8000 6 N4BEG[7]
port 75 nsew signal output
rlabel metal2 s 13450 7840 13506 8000 6 N4BEG[8]
port 76 nsew signal output
rlabel metal2 s 13726 7840 13782 8000 6 N4BEG[9]
port 77 nsew signal output
rlabel metal2 s 15658 7840 15714 8000 6 NN4BEG[0]
port 78 nsew signal output
rlabel metal2 s 18418 7840 18474 8000 6 NN4BEG[10]
port 79 nsew signal output
rlabel metal2 s 18694 7840 18750 8000 6 NN4BEG[11]
port 80 nsew signal output
rlabel metal2 s 18970 7840 19026 8000 6 NN4BEG[12]
port 81 nsew signal output
rlabel metal2 s 19246 7840 19302 8000 6 NN4BEG[13]
port 82 nsew signal output
rlabel metal2 s 19522 7840 19578 8000 6 NN4BEG[14]
port 83 nsew signal output
rlabel metal2 s 19798 7840 19854 8000 6 NN4BEG[15]
port 84 nsew signal output
rlabel metal2 s 15934 7840 15990 8000 6 NN4BEG[1]
port 85 nsew signal output
rlabel metal2 s 16210 7840 16266 8000 6 NN4BEG[2]
port 86 nsew signal output
rlabel metal2 s 16486 7840 16542 8000 6 NN4BEG[3]
port 87 nsew signal output
rlabel metal2 s 16762 7840 16818 8000 6 NN4BEG[4]
port 88 nsew signal output
rlabel metal2 s 17038 7840 17094 8000 6 NN4BEG[5]
port 89 nsew signal output
rlabel metal2 s 17314 7840 17370 8000 6 NN4BEG[6]
port 90 nsew signal output
rlabel metal2 s 17590 7840 17646 8000 6 NN4BEG[7]
port 91 nsew signal output
rlabel metal2 s 17866 7840 17922 8000 6 NN4BEG[8]
port 92 nsew signal output
rlabel metal2 s 18142 7840 18198 8000 6 NN4BEG[9]
port 93 nsew signal output
rlabel metal2 s 20074 7840 20130 8000 6 S1END[0]
port 94 nsew signal input
rlabel metal2 s 20350 7840 20406 8000 6 S1END[1]
port 95 nsew signal input
rlabel metal2 s 20626 7840 20682 8000 6 S1END[2]
port 96 nsew signal input
rlabel metal2 s 20902 7840 20958 8000 6 S1END[3]
port 97 nsew signal input
rlabel metal2 s 21178 7840 21234 8000 6 S2END[0]
port 98 nsew signal input
rlabel metal2 s 21454 7840 21510 8000 6 S2END[1]
port 99 nsew signal input
rlabel metal2 s 21730 7840 21786 8000 6 S2END[2]
port 100 nsew signal input
rlabel metal2 s 22006 7840 22062 8000 6 S2END[3]
port 101 nsew signal input
rlabel metal2 s 22282 7840 22338 8000 6 S2END[4]
port 102 nsew signal input
rlabel metal2 s 22558 7840 22614 8000 6 S2END[5]
port 103 nsew signal input
rlabel metal2 s 22834 7840 22890 8000 6 S2END[6]
port 104 nsew signal input
rlabel metal2 s 23110 7840 23166 8000 6 S2END[7]
port 105 nsew signal input
rlabel metal2 s 23386 7840 23442 8000 6 S2MID[0]
port 106 nsew signal input
rlabel metal2 s 23662 7840 23718 8000 6 S2MID[1]
port 107 nsew signal input
rlabel metal2 s 23938 7840 23994 8000 6 S2MID[2]
port 108 nsew signal input
rlabel metal2 s 24214 7840 24270 8000 6 S2MID[3]
port 109 nsew signal input
rlabel metal2 s 24490 7840 24546 8000 6 S2MID[4]
port 110 nsew signal input
rlabel metal2 s 24766 7840 24822 8000 6 S2MID[5]
port 111 nsew signal input
rlabel metal2 s 25042 7840 25098 8000 6 S2MID[6]
port 112 nsew signal input
rlabel metal2 s 25318 7840 25374 8000 6 S2MID[7]
port 113 nsew signal input
rlabel metal2 s 25594 7840 25650 8000 6 S4END[0]
port 114 nsew signal input
rlabel metal2 s 28354 7840 28410 8000 6 S4END[10]
port 115 nsew signal input
rlabel metal2 s 28630 7840 28686 8000 6 S4END[11]
port 116 nsew signal input
rlabel metal2 s 28906 7840 28962 8000 6 S4END[12]
port 117 nsew signal input
rlabel metal2 s 29182 7840 29238 8000 6 S4END[13]
port 118 nsew signal input
rlabel metal2 s 29458 7840 29514 8000 6 S4END[14]
port 119 nsew signal input
rlabel metal2 s 29734 7840 29790 8000 6 S4END[15]
port 120 nsew signal input
rlabel metal2 s 25870 7840 25926 8000 6 S4END[1]
port 121 nsew signal input
rlabel metal2 s 26146 7840 26202 8000 6 S4END[2]
port 122 nsew signal input
rlabel metal2 s 26422 7840 26478 8000 6 S4END[3]
port 123 nsew signal input
rlabel metal2 s 26698 7840 26754 8000 6 S4END[4]
port 124 nsew signal input
rlabel metal2 s 26974 7840 27030 8000 6 S4END[5]
port 125 nsew signal input
rlabel metal2 s 27250 7840 27306 8000 6 S4END[6]
port 126 nsew signal input
rlabel metal2 s 27526 7840 27582 8000 6 S4END[7]
port 127 nsew signal input
rlabel metal2 s 27802 7840 27858 8000 6 S4END[8]
port 128 nsew signal input
rlabel metal2 s 28078 7840 28134 8000 6 S4END[9]
port 129 nsew signal input
rlabel metal2 s 30010 7840 30066 8000 6 SS4END[0]
port 130 nsew signal input
rlabel metal2 s 32770 7840 32826 8000 6 SS4END[10]
port 131 nsew signal input
rlabel metal2 s 33046 7840 33102 8000 6 SS4END[11]
port 132 nsew signal input
rlabel metal2 s 33322 7840 33378 8000 6 SS4END[12]
port 133 nsew signal input
rlabel metal2 s 33598 7840 33654 8000 6 SS4END[13]
port 134 nsew signal input
rlabel metal2 s 33874 7840 33930 8000 6 SS4END[14]
port 135 nsew signal input
rlabel metal2 s 34150 7840 34206 8000 6 SS4END[15]
port 136 nsew signal input
rlabel metal2 s 30286 7840 30342 8000 6 SS4END[1]
port 137 nsew signal input
rlabel metal2 s 30562 7840 30618 8000 6 SS4END[2]
port 138 nsew signal input
rlabel metal2 s 30838 7840 30894 8000 6 SS4END[3]
port 139 nsew signal input
rlabel metal2 s 31114 7840 31170 8000 6 SS4END[4]
port 140 nsew signal input
rlabel metal2 s 31390 7840 31446 8000 6 SS4END[5]
port 141 nsew signal input
rlabel metal2 s 31666 7840 31722 8000 6 SS4END[6]
port 142 nsew signal input
rlabel metal2 s 31942 7840 31998 8000 6 SS4END[7]
port 143 nsew signal input
rlabel metal2 s 32218 7840 32274 8000 6 SS4END[8]
port 144 nsew signal input
rlabel metal2 s 32494 7840 32550 8000 6 SS4END[9]
port 145 nsew signal input
rlabel metal2 s 16302 0 16358 160 6 UIO_BOT_UIN0
port 146 nsew signal input
rlabel metal2 s 17038 0 17094 160 6 UIO_BOT_UIN1
port 147 nsew signal input
rlabel metal2 s 17774 0 17830 160 6 UIO_BOT_UIN10
port 148 nsew signal input
rlabel metal2 s 18510 0 18566 160 6 UIO_BOT_UIN11
port 149 nsew signal input
rlabel metal2 s 19246 0 19302 160 6 UIO_BOT_UIN12
port 150 nsew signal input
rlabel metal2 s 19982 0 20038 160 6 UIO_BOT_UIN13
port 151 nsew signal input
rlabel metal2 s 20718 0 20774 160 6 UIO_BOT_UIN14
port 152 nsew signal input
rlabel metal2 s 21454 0 21510 160 6 UIO_BOT_UIN15
port 153 nsew signal input
rlabel metal2 s 22190 0 22246 160 6 UIO_BOT_UIN16
port 154 nsew signal input
rlabel metal2 s 22926 0 22982 160 6 UIO_BOT_UIN17
port 155 nsew signal input
rlabel metal2 s 23662 0 23718 160 6 UIO_BOT_UIN18
port 156 nsew signal input
rlabel metal2 s 24398 0 24454 160 6 UIO_BOT_UIN19
port 157 nsew signal input
rlabel metal2 s 25134 0 25190 160 6 UIO_BOT_UIN2
port 158 nsew signal input
rlabel metal2 s 25870 0 25926 160 6 UIO_BOT_UIN3
port 159 nsew signal input
rlabel metal2 s 26606 0 26662 160 6 UIO_BOT_UIN4
port 160 nsew signal input
rlabel metal2 s 27342 0 27398 160 6 UIO_BOT_UIN5
port 161 nsew signal input
rlabel metal2 s 28078 0 28134 160 6 UIO_BOT_UIN6
port 162 nsew signal input
rlabel metal2 s 28814 0 28870 160 6 UIO_BOT_UIN7
port 163 nsew signal input
rlabel metal2 s 29550 0 29606 160 6 UIO_BOT_UIN8
port 164 nsew signal input
rlabel metal2 s 30286 0 30342 160 6 UIO_BOT_UIN9
port 165 nsew signal input
rlabel metal2 s 31022 0 31078 160 6 UIO_BOT_UOUT0
port 166 nsew signal output
rlabel metal2 s 31758 0 31814 160 6 UIO_BOT_UOUT1
port 167 nsew signal output
rlabel metal2 s 32494 0 32550 160 6 UIO_BOT_UOUT10
port 168 nsew signal output
rlabel metal2 s 33230 0 33286 160 6 UIO_BOT_UOUT11
port 169 nsew signal output
rlabel metal2 s 33966 0 34022 160 6 UIO_BOT_UOUT12
port 170 nsew signal output
rlabel metal2 s 34702 0 34758 160 6 UIO_BOT_UOUT13
port 171 nsew signal output
rlabel metal2 s 35438 0 35494 160 6 UIO_BOT_UOUT14
port 172 nsew signal output
rlabel metal2 s 36174 0 36230 160 6 UIO_BOT_UOUT15
port 173 nsew signal output
rlabel metal2 s 36910 0 36966 160 6 UIO_BOT_UOUT16
port 174 nsew signal output
rlabel metal2 s 37646 0 37702 160 6 UIO_BOT_UOUT17
port 175 nsew signal output
rlabel metal2 s 38382 0 38438 160 6 UIO_BOT_UOUT18
port 176 nsew signal output
rlabel metal2 s 39118 0 39174 160 6 UIO_BOT_UOUT19
port 177 nsew signal output
rlabel metal2 s 39854 0 39910 160 6 UIO_BOT_UOUT2
port 178 nsew signal output
rlabel metal2 s 40590 0 40646 160 6 UIO_BOT_UOUT3
port 179 nsew signal output
rlabel metal2 s 41326 0 41382 160 6 UIO_BOT_UOUT4
port 180 nsew signal output
rlabel metal2 s 42062 0 42118 160 6 UIO_BOT_UOUT5
port 181 nsew signal output
rlabel metal2 s 42798 0 42854 160 6 UIO_BOT_UOUT6
port 182 nsew signal output
rlabel metal2 s 43534 0 43590 160 6 UIO_BOT_UOUT7
port 183 nsew signal output
rlabel metal2 s 44270 0 44326 160 6 UIO_BOT_UOUT8
port 184 nsew signal output
rlabel metal2 s 45006 0 45062 160 6 UIO_BOT_UOUT9
port 185 nsew signal output
rlabel metal2 s 846 0 902 160 6 UserCLK
port 186 nsew signal input
rlabel metal2 s 34426 7840 34482 8000 6 UserCLKo
port 187 nsew signal output
rlabel metal4 s 6417 2128 6737 5488 6 vccd1
port 188 nsew power bidirectional
rlabel metal4 s 17364 2128 17684 5488 6 vccd1
port 188 nsew power bidirectional
rlabel metal4 s 28311 2128 28631 5488 6 vccd1
port 188 nsew power bidirectional
rlabel metal4 s 39258 2128 39578 5488 6 vccd1
port 188 nsew power bidirectional
rlabel metal4 s 11890 2128 12210 5488 6 vssd1
port 189 nsew ground bidirectional
rlabel metal4 s 22837 2128 23157 5488 6 vssd1
port 189 nsew ground bidirectional
rlabel metal4 s 33784 2128 34104 5488 6 vssd1
port 189 nsew ground bidirectional
rlabel metal4 s 44731 2128 45051 5488 6 vssd1
port 189 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 46000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 544600
string GDS_FILE /home/user/Desktop/FPGA_IGNITE_2024/openlane/S_term_Tiles/runs/24_11_24_00_41/results/signoff/S_term_single.magic.gds
string GDS_START 49188
<< end >>

