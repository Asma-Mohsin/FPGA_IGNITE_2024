VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_IO
  CLASS BLOCK ;
  FOREIGN W_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 181.000 BY 231.000 ;
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.310 0.700 161.690 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.830 0.700 171.210 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.070 0.700 166.450 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.870 0.700 190.250 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.310 0.700 195.690 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.070 0.700 200.450 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.830 0.700 205.210 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.590 0.700 175.970 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.110 0.700 185.490 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.350 0.700 180.730 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.590 0.700 209.970 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.350 0.700 214.730 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.110 0.700 219.490 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.870 0.700 224.250 ;
    END
  END B_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 3.550 181.000 3.930 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 5.590 181.000 5.970 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 6.950 181.000 7.330 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 8.990 181.000 9.370 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 10.350 181.000 10.730 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 12.390 181.000 12.770 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 13.750 181.000 14.130 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 15.790 181.000 16.170 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 17.150 181.000 17.530 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 19.190 181.000 19.570 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 21.230 181.000 21.610 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 22.590 181.000 22.970 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 24.630 181.000 25.010 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 25.990 181.000 26.370 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 28.030 181.000 28.410 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 29.390 181.000 29.770 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 31.430 181.000 31.810 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 33.470 181.000 33.850 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 34.830 181.000 35.210 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 36.870 181.000 37.250 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 66.110 181.000 66.490 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 83.790 181.000 84.170 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 85.150 181.000 85.530 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 68.150 181.000 68.530 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 69.510 181.000 69.890 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 71.550 181.000 71.930 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 72.910 181.000 73.290 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 74.950 181.000 75.330 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 76.310 181.000 76.690 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 78.350 181.000 78.730 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 80.390 181.000 80.770 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 81.750 181.000 82.130 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 38.230 181.000 38.610 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 55.910 181.000 56.290 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 57.270 181.000 57.650 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 59.310 181.000 59.690 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 60.670 181.000 61.050 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 62.710 181.000 63.090 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 64.750 181.000 65.130 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 40.270 181.000 40.650 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 41.630 181.000 42.010 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 43.670 181.000 44.050 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 45.030 181.000 45.410 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 47.070 181.000 47.450 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 49.110 181.000 49.490 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 50.470 181.000 50.850 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 52.510 181.000 52.890 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 53.870 181.000 54.250 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.950 0.700 7.330 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.230 0.700 55.610 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.990 0.700 60.370 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.750 0.700 65.130 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.510 0.700 69.890 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.270 0.700 74.650 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.030 0.700 79.410 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.790 0.700 84.170 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.550 0.700 88.930 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.310 0.700 93.690 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.750 0.700 99.130 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.710 0.700 12.090 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.510 0.700 103.890 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.270 0.700 108.650 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.030 0.700 113.410 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.790 0.700 118.170 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.550 0.700 122.930 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.310 0.700 127.690 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.070 0.700 132.450 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.830 0.700 137.210 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.590 0.700 141.970 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.030 0.700 147.410 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.470 0.700 16.850 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.790 0.700 152.170 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.550 0.700 156.930 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.230 0.700 21.610 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.990 0.700 26.370 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.750 0.700 31.130 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.510 0.700 35.890 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.270 0.700 40.650 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.030 0.700 45.410 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.790 0.700 50.170 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 170.830 181.000 171.210 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 187.830 181.000 188.210 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 189.870 181.000 190.250 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 191.230 181.000 191.610 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 193.270 181.000 193.650 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 194.630 181.000 195.010 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 196.670 181.000 197.050 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 198.710 181.000 199.090 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 200.070 181.000 200.450 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 202.110 181.000 202.490 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 203.470 181.000 203.850 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 172.190 181.000 172.570 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 205.510 181.000 205.890 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 206.870 181.000 207.250 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 208.910 181.000 209.290 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 210.950 181.000 211.330 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 212.310 181.000 212.690 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 214.350 181.000 214.730 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 215.710 181.000 216.090 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 217.750 181.000 218.130 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 219.110 181.000 219.490 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 221.150 181.000 221.530 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 174.230 181.000 174.610 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 222.510 181.000 222.890 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 224.550 181.000 224.930 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 175.590 181.000 175.970 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 177.630 181.000 178.010 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 178.990 181.000 179.370 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 181.030 181.000 181.410 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 183.070 181.000 183.450 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 184.430 181.000 184.810 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 186.470 181.000 186.850 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 9.700 0.000 10.080 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.200 0.000 90.580 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 98.480 0.000 98.860 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.300 0.000 106.680 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 114.580 0.000 114.960 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 122.400 0.000 122.780 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 130.680 0.000 131.060 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 138.500 0.000 138.880 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 146.320 0.000 146.700 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 154.600 0.000 154.980 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 162.420 0.000 162.800 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 17.980 0.000 18.360 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 25.800 0.000 26.180 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 34.080 0.000 34.460 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.900 0.000 42.280 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 50.180 0.000 50.560 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.000 0.000 58.380 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 66.280 0.000 66.660 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.100 0.000 74.480 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 82.380 0.000 82.760 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.700 230.300 10.080 231.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.200 230.300 90.580 231.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.480 230.300 98.860 231.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.300 230.300 106.680 231.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.580 230.300 114.960 231.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.400 230.300 122.780 231.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.680 230.300 131.060 231.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.500 230.300 138.880 231.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 230.300 146.700 231.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.600 230.300 154.980 231.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.420 230.300 162.800 231.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.980 230.300 18.360 231.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.800 230.300 26.180 231.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 34.080 230.300 34.460 231.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.900 230.300 42.280 231.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.180 230.300 50.560 231.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 230.300 58.380 231.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.280 230.300 66.660 231.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.100 230.300 74.480 231.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.380 230.300 82.760 231.000 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 170.700 0.000 171.080 0.700 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 170.700 230.300 171.080 231.000 ;
    END
  END UserCLKo
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 87.190 181.000 87.570 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 88.550 181.000 88.930 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 90.590 181.000 90.970 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 92.630 181.000 93.010 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 108.270 181.000 108.650 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 109.630 181.000 110.010 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 111.670 181.000 112.050 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 113.030 181.000 113.410 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 115.070 181.000 115.450 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 116.430 181.000 116.810 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 118.470 181.000 118.850 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 119.830 181.000 120.210 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 93.990 181.000 94.370 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 96.030 181.000 96.410 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 97.390 181.000 97.770 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 99.430 181.000 99.810 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 100.790 181.000 101.170 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 102.830 181.000 103.210 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 104.190 181.000 104.570 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 106.230 181.000 106.610 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 149.750 181.000 150.130 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 167.430 181.000 167.810 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 168.790 181.000 169.170 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 151.790 181.000 152.170 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 153.150 181.000 153.530 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 155.190 181.000 155.570 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 156.550 181.000 156.930 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 158.590 181.000 158.970 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 159.950 181.000 160.330 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 161.990 181.000 162.370 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 163.350 181.000 163.730 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 165.390 181.000 165.770 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 121.870 181.000 122.250 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 139.550 181.000 139.930 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 140.910 181.000 141.290 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 180.300 142.950 181.000 143.330 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 144.310 181.000 144.690 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 146.350 181.000 146.730 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 147.710 181.000 148.090 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 123.910 181.000 124.290 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 125.270 181.000 125.650 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 127.310 181.000 127.690 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 128.670 181.000 129.050 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 130.710 181.000 131.090 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 132.070 181.000 132.450 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 134.110 181.000 134.490 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 135.470 181.000 135.850 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 137.510 181.000 137.890 ;
    END
  END WW4END[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -12.040 -11.660 -8.940 242.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 -11.660 192.820 -8.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 239.760 192.820 242.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 -11.660 192.820 242.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.580 -16.460 22.180 247.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 -16.460 175.780 247.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 21.290 197.620 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 174.470 197.620 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.840 -16.460 -13.740 247.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 -16.460 197.620 -13.360 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 244.560 197.620 247.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 194.520 -16.460 197.620 247.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.880 -16.460 25.480 247.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 24.590 197.620 26.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 177.770 197.620 179.370 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 4.870 5.355 175.910 225.950 ;
      LAYER li1 ;
        RECT 5.060 5.355 175.720 225.845 ;
      LAYER met1 ;
        RECT 1.910 4.800 179.330 226.000 ;
      LAYER met2 ;
        RECT 1.930 230.020 9.420 230.300 ;
        RECT 10.360 230.020 17.700 230.300 ;
        RECT 18.640 230.020 25.520 230.300 ;
        RECT 26.460 230.020 33.800 230.300 ;
        RECT 34.740 230.020 41.620 230.300 ;
        RECT 42.560 230.020 49.900 230.300 ;
        RECT 50.840 230.020 57.720 230.300 ;
        RECT 58.660 230.020 66.000 230.300 ;
        RECT 66.940 230.020 73.820 230.300 ;
        RECT 74.760 230.020 82.100 230.300 ;
        RECT 83.040 230.020 89.920 230.300 ;
        RECT 90.860 230.020 98.200 230.300 ;
        RECT 99.140 230.020 106.020 230.300 ;
        RECT 106.960 230.020 114.300 230.300 ;
        RECT 115.240 230.020 122.120 230.300 ;
        RECT 123.060 230.020 130.400 230.300 ;
        RECT 131.340 230.020 138.220 230.300 ;
        RECT 139.160 230.020 146.040 230.300 ;
        RECT 146.980 230.020 154.320 230.300 ;
        RECT 155.260 230.020 162.140 230.300 ;
        RECT 163.080 230.020 170.420 230.300 ;
        RECT 171.360 230.020 179.310 230.300 ;
        RECT 1.930 0.980 179.310 230.020 ;
        RECT 1.930 0.700 9.420 0.980 ;
        RECT 10.360 0.700 17.700 0.980 ;
        RECT 18.640 0.700 25.520 0.980 ;
        RECT 26.460 0.700 33.800 0.980 ;
        RECT 34.740 0.700 41.620 0.980 ;
        RECT 42.560 0.700 49.900 0.980 ;
        RECT 50.840 0.700 57.720 0.980 ;
        RECT 58.660 0.700 66.000 0.980 ;
        RECT 66.940 0.700 73.820 0.980 ;
        RECT 74.760 0.700 82.100 0.980 ;
        RECT 83.040 0.700 89.920 0.980 ;
        RECT 90.860 0.700 98.200 0.980 ;
        RECT 99.140 0.700 106.020 0.980 ;
        RECT 106.960 0.700 114.300 0.980 ;
        RECT 115.240 0.700 122.120 0.980 ;
        RECT 123.060 0.700 130.400 0.980 ;
        RECT 131.340 0.700 138.220 0.980 ;
        RECT 139.160 0.700 146.040 0.980 ;
        RECT 146.980 0.700 154.320 0.980 ;
        RECT 155.260 0.700 162.140 0.980 ;
        RECT 163.080 0.700 170.420 0.980 ;
        RECT 171.360 0.700 179.310 0.980 ;
      LAYER met3 ;
        RECT 0.700 225.330 180.300 225.925 ;
        RECT 0.700 224.650 179.900 225.330 ;
        RECT 1.100 224.150 179.900 224.650 ;
        RECT 1.100 223.470 180.300 224.150 ;
        RECT 0.700 223.290 180.300 223.470 ;
        RECT 0.700 222.110 179.900 223.290 ;
        RECT 0.700 221.930 180.300 222.110 ;
        RECT 0.700 220.750 179.900 221.930 ;
        RECT 0.700 219.890 180.300 220.750 ;
        RECT 1.100 218.710 179.900 219.890 ;
        RECT 0.700 218.530 180.300 218.710 ;
        RECT 0.700 217.350 179.900 218.530 ;
        RECT 0.700 216.490 180.300 217.350 ;
        RECT 0.700 215.310 179.900 216.490 ;
        RECT 0.700 215.130 180.300 215.310 ;
        RECT 1.100 213.950 179.900 215.130 ;
        RECT 0.700 213.090 180.300 213.950 ;
        RECT 0.700 211.910 179.900 213.090 ;
        RECT 0.700 211.730 180.300 211.910 ;
        RECT 0.700 210.550 179.900 211.730 ;
        RECT 0.700 210.370 180.300 210.550 ;
        RECT 1.100 209.690 180.300 210.370 ;
        RECT 1.100 209.190 179.900 209.690 ;
        RECT 0.700 208.510 179.900 209.190 ;
        RECT 0.700 207.650 180.300 208.510 ;
        RECT 0.700 206.470 179.900 207.650 ;
        RECT 0.700 206.290 180.300 206.470 ;
        RECT 0.700 205.610 179.900 206.290 ;
        RECT 1.100 205.110 179.900 205.610 ;
        RECT 1.100 204.430 180.300 205.110 ;
        RECT 0.700 204.250 180.300 204.430 ;
        RECT 0.700 203.070 179.900 204.250 ;
        RECT 0.700 202.890 180.300 203.070 ;
        RECT 0.700 201.710 179.900 202.890 ;
        RECT 0.700 200.850 180.300 201.710 ;
        RECT 1.100 199.670 179.900 200.850 ;
        RECT 0.700 199.490 180.300 199.670 ;
        RECT 0.700 198.310 179.900 199.490 ;
        RECT 0.700 197.450 180.300 198.310 ;
        RECT 0.700 196.270 179.900 197.450 ;
        RECT 0.700 196.090 180.300 196.270 ;
        RECT 1.100 195.410 180.300 196.090 ;
        RECT 1.100 194.910 179.900 195.410 ;
        RECT 0.700 194.230 179.900 194.910 ;
        RECT 0.700 194.050 180.300 194.230 ;
        RECT 0.700 192.870 179.900 194.050 ;
        RECT 0.700 192.010 180.300 192.870 ;
        RECT 0.700 190.830 179.900 192.010 ;
        RECT 0.700 190.650 180.300 190.830 ;
        RECT 1.100 189.470 179.900 190.650 ;
        RECT 0.700 188.610 180.300 189.470 ;
        RECT 0.700 187.430 179.900 188.610 ;
        RECT 0.700 187.250 180.300 187.430 ;
        RECT 0.700 186.070 179.900 187.250 ;
        RECT 0.700 185.890 180.300 186.070 ;
        RECT 1.100 185.210 180.300 185.890 ;
        RECT 1.100 184.710 179.900 185.210 ;
        RECT 0.700 184.030 179.900 184.710 ;
        RECT 0.700 183.850 180.300 184.030 ;
        RECT 0.700 182.670 179.900 183.850 ;
        RECT 0.700 181.810 180.300 182.670 ;
        RECT 0.700 181.130 179.900 181.810 ;
        RECT 1.100 180.630 179.900 181.130 ;
        RECT 1.100 179.950 180.300 180.630 ;
        RECT 0.700 179.770 180.300 179.950 ;
        RECT 0.700 178.590 179.900 179.770 ;
        RECT 0.700 178.410 180.300 178.590 ;
        RECT 0.700 177.230 179.900 178.410 ;
        RECT 0.700 176.370 180.300 177.230 ;
        RECT 1.100 175.190 179.900 176.370 ;
        RECT 0.700 175.010 180.300 175.190 ;
        RECT 0.700 173.830 179.900 175.010 ;
        RECT 0.700 172.970 180.300 173.830 ;
        RECT 0.700 171.790 179.900 172.970 ;
        RECT 0.700 171.610 180.300 171.790 ;
        RECT 1.100 170.430 179.900 171.610 ;
        RECT 0.700 169.570 180.300 170.430 ;
        RECT 0.700 168.390 179.900 169.570 ;
        RECT 0.700 168.210 180.300 168.390 ;
        RECT 0.700 167.030 179.900 168.210 ;
        RECT 0.700 166.850 180.300 167.030 ;
        RECT 1.100 166.170 180.300 166.850 ;
        RECT 1.100 165.670 179.900 166.170 ;
        RECT 0.700 164.990 179.900 165.670 ;
        RECT 0.700 164.130 180.300 164.990 ;
        RECT 0.700 162.950 179.900 164.130 ;
        RECT 0.700 162.770 180.300 162.950 ;
        RECT 0.700 162.090 179.900 162.770 ;
        RECT 1.100 161.590 179.900 162.090 ;
        RECT 1.100 160.910 180.300 161.590 ;
        RECT 0.700 160.730 180.300 160.910 ;
        RECT 0.700 159.550 179.900 160.730 ;
        RECT 0.700 159.370 180.300 159.550 ;
        RECT 0.700 158.190 179.900 159.370 ;
        RECT 0.700 157.330 180.300 158.190 ;
        RECT 1.100 156.150 179.900 157.330 ;
        RECT 0.700 155.970 180.300 156.150 ;
        RECT 0.700 154.790 179.900 155.970 ;
        RECT 0.700 153.930 180.300 154.790 ;
        RECT 0.700 152.750 179.900 153.930 ;
        RECT 0.700 152.570 180.300 152.750 ;
        RECT 1.100 151.390 179.900 152.570 ;
        RECT 0.700 150.530 180.300 151.390 ;
        RECT 0.700 149.350 179.900 150.530 ;
        RECT 0.700 148.490 180.300 149.350 ;
        RECT 0.700 147.810 179.900 148.490 ;
        RECT 1.100 147.310 179.900 147.810 ;
        RECT 1.100 147.130 180.300 147.310 ;
        RECT 1.100 146.630 179.900 147.130 ;
        RECT 0.700 145.950 179.900 146.630 ;
        RECT 0.700 145.090 180.300 145.950 ;
        RECT 0.700 143.910 179.900 145.090 ;
        RECT 0.700 143.730 180.300 143.910 ;
        RECT 0.700 142.550 179.900 143.730 ;
        RECT 0.700 142.370 180.300 142.550 ;
        RECT 1.100 141.690 180.300 142.370 ;
        RECT 1.100 141.190 179.900 141.690 ;
        RECT 0.700 140.510 179.900 141.190 ;
        RECT 0.700 140.330 180.300 140.510 ;
        RECT 0.700 139.150 179.900 140.330 ;
        RECT 0.700 138.290 180.300 139.150 ;
        RECT 0.700 137.610 179.900 138.290 ;
        RECT 1.100 137.110 179.900 137.610 ;
        RECT 1.100 136.430 180.300 137.110 ;
        RECT 0.700 136.250 180.300 136.430 ;
        RECT 0.700 135.070 179.900 136.250 ;
        RECT 0.700 134.890 180.300 135.070 ;
        RECT 0.700 133.710 179.900 134.890 ;
        RECT 0.700 132.850 180.300 133.710 ;
        RECT 1.100 131.670 179.900 132.850 ;
        RECT 0.700 131.490 180.300 131.670 ;
        RECT 0.700 130.310 179.900 131.490 ;
        RECT 0.700 129.450 180.300 130.310 ;
        RECT 0.700 128.270 179.900 129.450 ;
        RECT 0.700 128.090 180.300 128.270 ;
        RECT 1.100 126.910 179.900 128.090 ;
        RECT 0.700 126.050 180.300 126.910 ;
        RECT 0.700 124.870 179.900 126.050 ;
        RECT 0.700 124.690 180.300 124.870 ;
        RECT 0.700 123.510 179.900 124.690 ;
        RECT 0.700 123.330 180.300 123.510 ;
        RECT 1.100 122.650 180.300 123.330 ;
        RECT 1.100 122.150 179.900 122.650 ;
        RECT 0.700 121.470 179.900 122.150 ;
        RECT 0.700 120.610 180.300 121.470 ;
        RECT 0.700 119.430 179.900 120.610 ;
        RECT 0.700 119.250 180.300 119.430 ;
        RECT 0.700 118.570 179.900 119.250 ;
        RECT 1.100 118.070 179.900 118.570 ;
        RECT 1.100 117.390 180.300 118.070 ;
        RECT 0.700 117.210 180.300 117.390 ;
        RECT 0.700 116.030 179.900 117.210 ;
        RECT 0.700 115.850 180.300 116.030 ;
        RECT 0.700 114.670 179.900 115.850 ;
        RECT 0.700 113.810 180.300 114.670 ;
        RECT 1.100 112.630 179.900 113.810 ;
        RECT 0.700 112.450 180.300 112.630 ;
        RECT 0.700 111.270 179.900 112.450 ;
        RECT 0.700 110.410 180.300 111.270 ;
        RECT 0.700 109.230 179.900 110.410 ;
        RECT 0.700 109.050 180.300 109.230 ;
        RECT 1.100 107.870 179.900 109.050 ;
        RECT 0.700 107.010 180.300 107.870 ;
        RECT 0.700 105.830 179.900 107.010 ;
        RECT 0.700 104.970 180.300 105.830 ;
        RECT 0.700 104.290 179.900 104.970 ;
        RECT 1.100 103.790 179.900 104.290 ;
        RECT 1.100 103.610 180.300 103.790 ;
        RECT 1.100 103.110 179.900 103.610 ;
        RECT 0.700 102.430 179.900 103.110 ;
        RECT 0.700 101.570 180.300 102.430 ;
        RECT 0.700 100.390 179.900 101.570 ;
        RECT 0.700 100.210 180.300 100.390 ;
        RECT 0.700 99.530 179.900 100.210 ;
        RECT 1.100 99.030 179.900 99.530 ;
        RECT 1.100 98.350 180.300 99.030 ;
        RECT 0.700 98.170 180.300 98.350 ;
        RECT 0.700 96.990 179.900 98.170 ;
        RECT 0.700 96.810 180.300 96.990 ;
        RECT 0.700 95.630 179.900 96.810 ;
        RECT 0.700 94.770 180.300 95.630 ;
        RECT 0.700 94.090 179.900 94.770 ;
        RECT 1.100 93.590 179.900 94.090 ;
        RECT 1.100 93.410 180.300 93.590 ;
        RECT 1.100 92.910 179.900 93.410 ;
        RECT 0.700 92.230 179.900 92.910 ;
        RECT 0.700 91.370 180.300 92.230 ;
        RECT 0.700 90.190 179.900 91.370 ;
        RECT 0.700 89.330 180.300 90.190 ;
        RECT 1.100 88.150 179.900 89.330 ;
        RECT 0.700 87.970 180.300 88.150 ;
        RECT 0.700 86.790 179.900 87.970 ;
        RECT 0.700 85.930 180.300 86.790 ;
        RECT 0.700 84.750 179.900 85.930 ;
        RECT 0.700 84.570 180.300 84.750 ;
        RECT 1.100 83.390 179.900 84.570 ;
        RECT 0.700 82.530 180.300 83.390 ;
        RECT 0.700 81.350 179.900 82.530 ;
        RECT 0.700 81.170 180.300 81.350 ;
        RECT 0.700 79.990 179.900 81.170 ;
        RECT 0.700 79.810 180.300 79.990 ;
        RECT 1.100 79.130 180.300 79.810 ;
        RECT 1.100 78.630 179.900 79.130 ;
        RECT 0.700 77.950 179.900 78.630 ;
        RECT 0.700 77.090 180.300 77.950 ;
        RECT 0.700 75.910 179.900 77.090 ;
        RECT 0.700 75.730 180.300 75.910 ;
        RECT 0.700 75.050 179.900 75.730 ;
        RECT 1.100 74.550 179.900 75.050 ;
        RECT 1.100 73.870 180.300 74.550 ;
        RECT 0.700 73.690 180.300 73.870 ;
        RECT 0.700 72.510 179.900 73.690 ;
        RECT 0.700 72.330 180.300 72.510 ;
        RECT 0.700 71.150 179.900 72.330 ;
        RECT 0.700 70.290 180.300 71.150 ;
        RECT 1.100 69.110 179.900 70.290 ;
        RECT 0.700 68.930 180.300 69.110 ;
        RECT 0.700 67.750 179.900 68.930 ;
        RECT 0.700 66.890 180.300 67.750 ;
        RECT 0.700 65.710 179.900 66.890 ;
        RECT 0.700 65.530 180.300 65.710 ;
        RECT 1.100 64.350 179.900 65.530 ;
        RECT 0.700 63.490 180.300 64.350 ;
        RECT 0.700 62.310 179.900 63.490 ;
        RECT 0.700 61.450 180.300 62.310 ;
        RECT 0.700 60.770 179.900 61.450 ;
        RECT 1.100 60.270 179.900 60.770 ;
        RECT 1.100 60.090 180.300 60.270 ;
        RECT 1.100 59.590 179.900 60.090 ;
        RECT 0.700 58.910 179.900 59.590 ;
        RECT 0.700 58.050 180.300 58.910 ;
        RECT 0.700 56.870 179.900 58.050 ;
        RECT 0.700 56.690 180.300 56.870 ;
        RECT 0.700 56.010 179.900 56.690 ;
        RECT 1.100 55.510 179.900 56.010 ;
        RECT 1.100 54.830 180.300 55.510 ;
        RECT 0.700 54.650 180.300 54.830 ;
        RECT 0.700 53.470 179.900 54.650 ;
        RECT 0.700 53.290 180.300 53.470 ;
        RECT 0.700 52.110 179.900 53.290 ;
        RECT 0.700 51.250 180.300 52.110 ;
        RECT 0.700 50.570 179.900 51.250 ;
        RECT 1.100 50.070 179.900 50.570 ;
        RECT 1.100 49.890 180.300 50.070 ;
        RECT 1.100 49.390 179.900 49.890 ;
        RECT 0.700 48.710 179.900 49.390 ;
        RECT 0.700 47.850 180.300 48.710 ;
        RECT 0.700 46.670 179.900 47.850 ;
        RECT 0.700 45.810 180.300 46.670 ;
        RECT 1.100 44.630 179.900 45.810 ;
        RECT 0.700 44.450 180.300 44.630 ;
        RECT 0.700 43.270 179.900 44.450 ;
        RECT 0.700 42.410 180.300 43.270 ;
        RECT 0.700 41.230 179.900 42.410 ;
        RECT 0.700 41.050 180.300 41.230 ;
        RECT 1.100 39.870 179.900 41.050 ;
        RECT 0.700 39.010 180.300 39.870 ;
        RECT 0.700 37.830 179.900 39.010 ;
        RECT 0.700 37.650 180.300 37.830 ;
        RECT 0.700 36.470 179.900 37.650 ;
        RECT 0.700 36.290 180.300 36.470 ;
        RECT 1.100 35.610 180.300 36.290 ;
        RECT 1.100 35.110 179.900 35.610 ;
        RECT 0.700 34.430 179.900 35.110 ;
        RECT 0.700 34.250 180.300 34.430 ;
        RECT 0.700 33.070 179.900 34.250 ;
        RECT 0.700 32.210 180.300 33.070 ;
        RECT 0.700 31.530 179.900 32.210 ;
        RECT 1.100 31.030 179.900 31.530 ;
        RECT 1.100 30.350 180.300 31.030 ;
        RECT 0.700 30.170 180.300 30.350 ;
        RECT 0.700 28.990 179.900 30.170 ;
        RECT 0.700 28.810 180.300 28.990 ;
        RECT 0.700 27.630 179.900 28.810 ;
        RECT 0.700 26.770 180.300 27.630 ;
        RECT 1.100 25.590 179.900 26.770 ;
        RECT 0.700 25.410 180.300 25.590 ;
        RECT 0.700 24.230 179.900 25.410 ;
        RECT 0.700 23.370 180.300 24.230 ;
        RECT 0.700 22.190 179.900 23.370 ;
        RECT 0.700 22.010 180.300 22.190 ;
        RECT 1.100 20.830 179.900 22.010 ;
        RECT 0.700 19.970 180.300 20.830 ;
        RECT 0.700 18.790 179.900 19.970 ;
        RECT 0.700 17.930 180.300 18.790 ;
        RECT 0.700 17.250 179.900 17.930 ;
        RECT 1.100 16.750 179.900 17.250 ;
        RECT 1.100 16.570 180.300 16.750 ;
        RECT 1.100 16.070 179.900 16.570 ;
        RECT 0.700 15.390 179.900 16.070 ;
        RECT 0.700 14.530 180.300 15.390 ;
        RECT 0.700 13.350 179.900 14.530 ;
        RECT 0.700 13.170 180.300 13.350 ;
        RECT 0.700 12.490 179.900 13.170 ;
        RECT 1.100 11.990 179.900 12.490 ;
        RECT 1.100 11.310 180.300 11.990 ;
        RECT 0.700 11.130 180.300 11.310 ;
        RECT 0.700 9.950 179.900 11.130 ;
        RECT 0.700 9.770 180.300 9.950 ;
        RECT 0.700 8.590 179.900 9.770 ;
        RECT 0.700 7.730 180.300 8.590 ;
        RECT 1.100 6.550 179.900 7.730 ;
        RECT 0.700 6.370 180.300 6.550 ;
        RECT 0.700 5.190 179.900 6.370 ;
        RECT 0.700 4.330 180.300 5.190 ;
        RECT 0.700 3.575 179.900 4.330 ;
      LAYER met4 ;
        RECT 59.175 6.295 172.665 221.505 ;
  END
END W_IO
END LIBRARY

