VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 182.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.000 0.000 104.380 0.700 ;
    END
  END Ci
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.120 0.000 206.500 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 225.440 0.000 225.820 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 227.280 0.000 227.660 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 229.120 0.000 229.500 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 230.960 0.000 231.340 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 233.260 0.000 233.640 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 235.100 0.000 235.480 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 236.940 0.000 237.320 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 238.780 0.000 239.160 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 240.620 0.000 241.000 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 242.920 0.000 243.300 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 207.960 0.000 208.340 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.800 0.000 210.180 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 211.640 0.000 212.020 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 213.940 0.000 214.320 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 215.780 0.000 216.160 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 217.620 0.000 218.000 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 219.460 0.000 219.840 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 221.300 0.000 221.680 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 223.600 0.000 223.980 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 5.560 181.300 5.940 182.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.040 181.300 46.420 182.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.180 181.300 50.560 182.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 53.860 181.300 54.240 182.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 181.300 58.380 182.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 62.140 181.300 62.520 182.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.280 181.300 66.660 182.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 69.960 181.300 70.340 182.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.100 181.300 74.480 182.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.240 181.300 78.620 182.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.380 181.300 82.760 182.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.700 181.300 10.080 182.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 13.840 181.300 14.220 182.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.520 181.300 17.900 182.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 21.660 181.300 22.040 182.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.800 181.300 26.180 182.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.940 181.300 30.320 182.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 33.620 181.300 34.000 182.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.760 181.300 38.140 182.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.900 181.300 42.280 182.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 3.720 0.000 4.100 0.700 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 5.560 0.000 5.940 0.700 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 7.400 0.000 7.780 0.700 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 9.240 0.000 9.620 0.700 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 26.720 0.000 27.100 0.700 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 28.560 0.000 28.940 0.700 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 30.400 0.000 30.780 0.700 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.240 0.000 32.620 0.700 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 34.540 0.000 34.920 0.700 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 36.380 0.000 36.760 0.700 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 38.220 0.000 38.600 0.700 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 40.060 0.000 40.440 0.700 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 11.080 0.000 11.460 0.700 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 13.380 0.000 13.760 0.700 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 15.220 0.000 15.600 0.700 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 17.060 0.000 17.440 0.700 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 18.900 0.000 19.280 0.700 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 20.740 0.000 21.120 0.700 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 22.580 0.000 22.960 0.700 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 24.880 0.000 25.260 0.700 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.900 0.000 42.280 0.700 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 61.220 0.000 61.600 0.700 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.520 0.000 63.900 0.700 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.360 0.000 65.740 0.700 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.200 0.000 67.580 0.700 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.040 0.000 69.420 0.700 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.880 0.000 71.260 0.700 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 44.200 0.000 44.580 0.700 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 46.040 0.000 46.420 0.700 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 47.880 0.000 48.260 0.700 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 49.720 0.000 50.100 0.700 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.560 0.000 51.940 0.700 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 53.860 0.000 54.240 0.700 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 55.700 0.000 56.080 0.700 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 57.540 0.000 57.920 0.700 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 59.380 0.000 59.760 0.700 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 73.180 0.000 73.560 0.700 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 92.040 0.000 92.420 0.700 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 94.340 0.000 94.720 0.700 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 96.180 0.000 96.560 0.700 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 98.020 0.000 98.400 0.700 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.860 0.000 100.240 0.700 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 101.700 0.000 102.080 0.700 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 75.020 0.000 75.400 0.700 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 76.860 0.000 77.240 0.700 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 78.700 0.000 79.080 0.700 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 80.540 0.000 80.920 0.700 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.380 0.000 82.760 0.700 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 84.680 0.000 85.060 0.700 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 0.000 86.900 0.700 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 88.360 0.000 88.740 0.700 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.200 0.000 90.580 0.700 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.840 0.000 106.220 0.700 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.680 0.000 108.060 0.700 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.520 0.000 109.900 0.700 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 111.360 0.000 111.740 0.700 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.660 0.000 114.040 0.700 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 115.500 0.000 115.880 0.700 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 117.340 0.000 117.720 0.700 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.180 0.000 119.560 0.700 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.020 0.000 121.400 0.700 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 123.320 0.000 123.700 0.700 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.160 0.000 125.540 0.700 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.000 0.000 127.380 0.700 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.840 0.000 129.220 0.700 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.680 0.000 131.060 0.700 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.980 0.000 133.360 0.700 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.820 0.000 135.200 0.700 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 136.660 0.000 137.040 0.700 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.500 0.000 138.880 0.700 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.340 0.000 140.720 0.700 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.180 0.000 142.560 0.700 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.480 0.000 144.860 0.700 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 163.800 0.000 164.180 0.700 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 165.640 0.000 166.020 0.700 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 167.480 0.000 167.860 0.700 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 169.320 0.000 169.700 0.700 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 171.160 0.000 171.540 0.700 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.460 0.000 173.840 0.700 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 0.000 146.700 0.700 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 148.160 0.000 148.540 0.700 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.000 0.000 150.380 0.700 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.840 0.000 152.220 0.700 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.140 0.000 154.520 0.700 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 155.980 0.000 156.360 0.700 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 157.820 0.000 158.200 0.700 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 159.660 0.000 160.040 0.700 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 161.500 0.000 161.880 0.700 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 175.300 0.000 175.680 0.700 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 194.620 0.000 195.000 0.700 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 196.460 0.000 196.840 0.700 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 198.300 0.000 198.680 0.700 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 200.140 0.000 200.520 0.700 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 201.980 0.000 202.360 0.700 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 204.280 0.000 204.660 0.700 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.140 0.000 177.520 0.700 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 178.980 0.000 179.360 0.700 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 180.820 0.000 181.200 0.700 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 183.120 0.000 183.500 0.700 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 184.960 0.000 185.340 0.700 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 186.800 0.000 187.180 0.700 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.640 0.000 189.020 0.700 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 190.480 0.000 190.860 0.700 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 192.780 0.000 193.160 0.700 ;
    END
  END SS4BEG[9]
  PIN UIO_TOP_UIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.020 181.300 167.400 182.000 ;
    END
  END UIO_TOP_UIN0
  PIN UIO_TOP_UIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 171.160 181.300 171.540 182.000 ;
    END
  END UIO_TOP_UIN1
  PIN UIO_TOP_UIN10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 174.840 181.300 175.220 182.000 ;
    END
  END UIO_TOP_UIN10
  PIN UIO_TOP_UIN11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 178.980 181.300 179.360 182.000 ;
    END
  END UIO_TOP_UIN11
  PIN UIO_TOP_UIN12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.120 181.300 183.500 182.000 ;
    END
  END UIO_TOP_UIN12
  PIN UIO_TOP_UIN13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 187.260 181.300 187.640 182.000 ;
    END
  END UIO_TOP_UIN13
  PIN UIO_TOP_UIN14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 190.940 181.300 191.320 182.000 ;
    END
  END UIO_TOP_UIN14
  PIN UIO_TOP_UIN15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 195.080 181.300 195.460 182.000 ;
    END
  END UIO_TOP_UIN15
  PIN UIO_TOP_UIN16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 199.220 181.300 199.600 182.000 ;
    END
  END UIO_TOP_UIN16
  PIN UIO_TOP_UIN17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 203.360 181.300 203.740 182.000 ;
    END
  END UIO_TOP_UIN17
  PIN UIO_TOP_UIN18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 207.040 181.300 207.420 182.000 ;
    END
  END UIO_TOP_UIN18
  PIN UIO_TOP_UIN19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 211.180 181.300 211.560 182.000 ;
    END
  END UIO_TOP_UIN19
  PIN UIO_TOP_UIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 215.320 181.300 215.700 182.000 ;
    END
  END UIO_TOP_UIN2
  PIN UIO_TOP_UIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 219.460 181.300 219.840 182.000 ;
    END
  END UIO_TOP_UIN3
  PIN UIO_TOP_UIN4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 223.600 181.300 223.980 182.000 ;
    END
  END UIO_TOP_UIN4
  PIN UIO_TOP_UIN5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 227.280 181.300 227.660 182.000 ;
    END
  END UIO_TOP_UIN5
  PIN UIO_TOP_UIN6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 231.420 181.300 231.800 182.000 ;
    END
  END UIO_TOP_UIN6
  PIN UIO_TOP_UIN7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 235.560 181.300 235.940 182.000 ;
    END
  END UIO_TOP_UIN7
  PIN UIO_TOP_UIN8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 239.700 181.300 240.080 182.000 ;
    END
  END UIO_TOP_UIN8
  PIN UIO_TOP_UIN9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 243.380 181.300 243.760 182.000 ;
    END
  END UIO_TOP_UIN9
  PIN UIO_TOP_UOUT0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.060 181.300 86.440 182.000 ;
    END
  END UIO_TOP_UOUT0
  PIN UIO_TOP_UOUT1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.200 181.300 90.580 182.000 ;
    END
  END UIO_TOP_UOUT1
  PIN UIO_TOP_UOUT10
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 94.340 181.300 94.720 182.000 ;
    END
  END UIO_TOP_UOUT10
  PIN UIO_TOP_UOUT11
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.480 181.300 98.860 182.000 ;
    END
  END UIO_TOP_UOUT11
  PIN UIO_TOP_UOUT12
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 102.620 181.300 103.000 182.000 ;
    END
  END UIO_TOP_UOUT12
  PIN UIO_TOP_UOUT13
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.300 181.300 106.680 182.000 ;
    END
  END UIO_TOP_UOUT13
  PIN UIO_TOP_UOUT14
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.440 181.300 110.820 182.000 ;
    END
  END UIO_TOP_UOUT14
  PIN UIO_TOP_UOUT15
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.580 181.300 114.960 182.000 ;
    END
  END UIO_TOP_UOUT15
  PIN UIO_TOP_UOUT16
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.720 181.300 119.100 182.000 ;
    END
  END UIO_TOP_UOUT16
  PIN UIO_TOP_UOUT17
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.400 181.300 122.780 182.000 ;
    END
  END UIO_TOP_UOUT17
  PIN UIO_TOP_UOUT18
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 126.540 181.300 126.920 182.000 ;
    END
  END UIO_TOP_UOUT18
  PIN UIO_TOP_UOUT19
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.680 181.300 131.060 182.000 ;
    END
  END UIO_TOP_UOUT19
  PIN UIO_TOP_UOUT2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.820 181.300 135.200 182.000 ;
    END
  END UIO_TOP_UOUT2
  PIN UIO_TOP_UOUT3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 138.500 181.300 138.880 182.000 ;
    END
  END UIO_TOP_UOUT3
  PIN UIO_TOP_UOUT4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 142.640 181.300 143.020 182.000 ;
    END
  END UIO_TOP_UOUT4
  PIN UIO_TOP_UOUT5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.780 181.300 147.160 182.000 ;
    END
  END UIO_TOP_UOUT5
  PIN UIO_TOP_UOUT6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.920 181.300 151.300 182.000 ;
    END
  END UIO_TOP_UOUT6
  PIN UIO_TOP_UOUT7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.060 181.300 155.440 182.000 ;
    END
  END UIO_TOP_UOUT7
  PIN UIO_TOP_UOUT8
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 158.740 181.300 159.120 182.000 ;
    END
  END UIO_TOP_UOUT8
  PIN UIO_TOP_UOUT9
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.880 181.300 163.260 182.000 ;
    END
  END UIO_TOP_UOUT9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 181.300 129.170 182.000 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 125.670 181.300 125.950 182.000 ;
    END
  END UserCLKo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.580 5.200 22.180 177.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 5.200 175.780 177.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 21.290 244.960 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 174.470 244.960 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.880 5.200 25.480 177.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.480 5.200 179.080 177.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 24.590 244.960 26.190 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 244.720 176.885 ;
      LAYER met1 ;
        RECT 3.750 1.060 244.720 178.120 ;
      LAYER met2 ;
        RECT 3.780 181.020 5.280 181.300 ;
        RECT 6.220 181.020 9.420 181.300 ;
        RECT 10.360 181.020 13.560 181.300 ;
        RECT 14.500 181.020 17.240 181.300 ;
        RECT 18.180 181.020 21.380 181.300 ;
        RECT 22.320 181.020 25.520 181.300 ;
        RECT 26.460 181.020 29.660 181.300 ;
        RECT 30.600 181.020 33.340 181.300 ;
        RECT 34.280 181.020 37.480 181.300 ;
        RECT 38.420 181.020 41.620 181.300 ;
        RECT 42.560 181.020 45.760 181.300 ;
        RECT 46.700 181.020 49.900 181.300 ;
        RECT 50.840 181.020 53.580 181.300 ;
        RECT 54.520 181.020 57.720 181.300 ;
        RECT 58.660 181.020 61.860 181.300 ;
        RECT 62.800 181.020 66.000 181.300 ;
        RECT 66.940 181.020 69.680 181.300 ;
        RECT 70.620 181.020 73.820 181.300 ;
        RECT 74.760 181.020 77.960 181.300 ;
        RECT 78.900 181.020 82.100 181.300 ;
        RECT 83.040 181.020 85.780 181.300 ;
        RECT 86.720 181.020 89.920 181.300 ;
        RECT 90.860 181.020 94.060 181.300 ;
        RECT 95.000 181.020 98.200 181.300 ;
        RECT 99.140 181.020 102.340 181.300 ;
        RECT 103.280 181.020 106.020 181.300 ;
        RECT 106.960 181.020 110.160 181.300 ;
        RECT 111.100 181.020 114.300 181.300 ;
        RECT 115.240 181.020 118.440 181.300 ;
        RECT 119.380 181.020 122.120 181.300 ;
        RECT 123.060 181.020 125.390 181.300 ;
        RECT 126.230 181.020 126.260 181.300 ;
        RECT 127.200 181.020 128.610 181.300 ;
        RECT 129.450 181.020 130.400 181.300 ;
        RECT 131.340 181.020 134.540 181.300 ;
        RECT 135.480 181.020 138.220 181.300 ;
        RECT 139.160 181.020 142.360 181.300 ;
        RECT 143.300 181.020 146.500 181.300 ;
        RECT 147.440 181.020 150.640 181.300 ;
        RECT 151.580 181.020 154.780 181.300 ;
        RECT 155.720 181.020 158.460 181.300 ;
        RECT 159.400 181.020 162.600 181.300 ;
        RECT 163.540 181.020 166.740 181.300 ;
        RECT 167.680 181.020 170.880 181.300 ;
        RECT 171.820 181.020 174.560 181.300 ;
        RECT 175.500 181.020 178.700 181.300 ;
        RECT 179.640 181.020 182.840 181.300 ;
        RECT 183.780 181.020 186.980 181.300 ;
        RECT 187.920 181.020 190.660 181.300 ;
        RECT 191.600 181.020 194.800 181.300 ;
        RECT 195.740 181.020 198.940 181.300 ;
        RECT 199.880 181.020 203.080 181.300 ;
        RECT 204.020 181.020 206.760 181.300 ;
        RECT 207.700 181.020 210.900 181.300 ;
        RECT 211.840 181.020 215.040 181.300 ;
        RECT 215.980 181.020 219.180 181.300 ;
        RECT 220.120 181.020 223.320 181.300 ;
        RECT 224.260 181.020 227.000 181.300 ;
        RECT 227.940 181.020 231.140 181.300 ;
        RECT 232.080 181.020 235.280 181.300 ;
        RECT 236.220 181.020 239.420 181.300 ;
        RECT 240.360 181.020 243.100 181.300 ;
        RECT 3.780 0.980 243.640 181.020 ;
        RECT 4.380 0.270 5.280 0.980 ;
        RECT 6.220 0.270 7.120 0.980 ;
        RECT 8.060 0.270 8.960 0.980 ;
        RECT 9.900 0.270 10.800 0.980 ;
        RECT 11.740 0.270 13.100 0.980 ;
        RECT 14.040 0.270 14.940 0.980 ;
        RECT 15.880 0.270 16.780 0.980 ;
        RECT 17.720 0.270 18.620 0.980 ;
        RECT 19.560 0.270 20.460 0.980 ;
        RECT 21.400 0.270 22.300 0.980 ;
        RECT 23.240 0.270 24.600 0.980 ;
        RECT 25.540 0.270 26.440 0.980 ;
        RECT 27.380 0.270 28.280 0.980 ;
        RECT 29.220 0.270 30.120 0.980 ;
        RECT 31.060 0.270 31.960 0.980 ;
        RECT 32.900 0.270 34.260 0.980 ;
        RECT 35.200 0.270 36.100 0.980 ;
        RECT 37.040 0.270 37.940 0.980 ;
        RECT 38.880 0.270 39.780 0.980 ;
        RECT 40.720 0.270 41.620 0.980 ;
        RECT 42.560 0.270 43.920 0.980 ;
        RECT 44.860 0.270 45.760 0.980 ;
        RECT 46.700 0.270 47.600 0.980 ;
        RECT 48.540 0.270 49.440 0.980 ;
        RECT 50.380 0.270 51.280 0.980 ;
        RECT 52.220 0.270 53.580 0.980 ;
        RECT 54.520 0.270 55.420 0.980 ;
        RECT 56.360 0.270 57.260 0.980 ;
        RECT 58.200 0.270 59.100 0.980 ;
        RECT 60.040 0.270 60.940 0.980 ;
        RECT 61.880 0.270 63.240 0.980 ;
        RECT 64.180 0.270 65.080 0.980 ;
        RECT 66.020 0.270 66.920 0.980 ;
        RECT 67.860 0.270 68.760 0.980 ;
        RECT 69.700 0.270 70.600 0.980 ;
        RECT 71.540 0.270 72.900 0.980 ;
        RECT 73.840 0.270 74.740 0.980 ;
        RECT 75.680 0.270 76.580 0.980 ;
        RECT 77.520 0.270 78.420 0.980 ;
        RECT 79.360 0.270 80.260 0.980 ;
        RECT 81.200 0.270 82.100 0.980 ;
        RECT 83.040 0.270 84.400 0.980 ;
        RECT 85.340 0.270 86.240 0.980 ;
        RECT 87.180 0.270 88.080 0.980 ;
        RECT 89.020 0.270 89.920 0.980 ;
        RECT 90.860 0.270 91.760 0.980 ;
        RECT 92.700 0.270 94.060 0.980 ;
        RECT 95.000 0.270 95.900 0.980 ;
        RECT 96.840 0.270 97.740 0.980 ;
        RECT 98.680 0.270 99.580 0.980 ;
        RECT 100.520 0.270 101.420 0.980 ;
        RECT 102.360 0.270 103.720 0.980 ;
        RECT 104.660 0.270 105.560 0.980 ;
        RECT 106.500 0.270 107.400 0.980 ;
        RECT 108.340 0.270 109.240 0.980 ;
        RECT 110.180 0.270 111.080 0.980 ;
        RECT 112.020 0.270 113.380 0.980 ;
        RECT 114.320 0.270 115.220 0.980 ;
        RECT 116.160 0.270 117.060 0.980 ;
        RECT 118.000 0.270 118.900 0.980 ;
        RECT 119.840 0.270 120.740 0.980 ;
        RECT 121.680 0.270 123.040 0.980 ;
        RECT 123.980 0.270 124.880 0.980 ;
        RECT 125.820 0.270 126.720 0.980 ;
        RECT 127.660 0.270 128.560 0.980 ;
        RECT 129.500 0.270 130.400 0.980 ;
        RECT 131.340 0.270 132.700 0.980 ;
        RECT 133.640 0.270 134.540 0.980 ;
        RECT 135.480 0.270 136.380 0.980 ;
        RECT 137.320 0.270 138.220 0.980 ;
        RECT 139.160 0.270 140.060 0.980 ;
        RECT 141.000 0.270 141.900 0.980 ;
        RECT 142.840 0.270 144.200 0.980 ;
        RECT 145.140 0.270 146.040 0.980 ;
        RECT 146.980 0.270 147.880 0.980 ;
        RECT 148.820 0.270 149.720 0.980 ;
        RECT 150.660 0.270 151.560 0.980 ;
        RECT 152.500 0.270 153.860 0.980 ;
        RECT 154.800 0.270 155.700 0.980 ;
        RECT 156.640 0.270 157.540 0.980 ;
        RECT 158.480 0.270 159.380 0.980 ;
        RECT 160.320 0.270 161.220 0.980 ;
        RECT 162.160 0.270 163.520 0.980 ;
        RECT 164.460 0.270 165.360 0.980 ;
        RECT 166.300 0.270 167.200 0.980 ;
        RECT 168.140 0.270 169.040 0.980 ;
        RECT 169.980 0.270 170.880 0.980 ;
        RECT 171.820 0.270 173.180 0.980 ;
        RECT 174.120 0.270 175.020 0.980 ;
        RECT 175.960 0.270 176.860 0.980 ;
        RECT 177.800 0.270 178.700 0.980 ;
        RECT 179.640 0.270 180.540 0.980 ;
        RECT 181.480 0.270 182.840 0.980 ;
        RECT 183.780 0.270 184.680 0.980 ;
        RECT 185.620 0.270 186.520 0.980 ;
        RECT 187.460 0.270 188.360 0.980 ;
        RECT 189.300 0.270 190.200 0.980 ;
        RECT 191.140 0.270 192.500 0.980 ;
        RECT 193.440 0.270 194.340 0.980 ;
        RECT 195.280 0.270 196.180 0.980 ;
        RECT 197.120 0.270 198.020 0.980 ;
        RECT 198.960 0.270 199.860 0.980 ;
        RECT 200.800 0.270 201.700 0.980 ;
        RECT 202.640 0.270 204.000 0.980 ;
        RECT 204.940 0.270 205.840 0.980 ;
        RECT 206.780 0.270 207.680 0.980 ;
        RECT 208.620 0.270 209.520 0.980 ;
        RECT 210.460 0.270 211.360 0.980 ;
        RECT 212.300 0.270 213.660 0.980 ;
        RECT 214.600 0.270 215.500 0.980 ;
        RECT 216.440 0.270 217.340 0.980 ;
        RECT 218.280 0.270 219.180 0.980 ;
        RECT 220.120 0.270 221.020 0.980 ;
        RECT 221.960 0.270 223.320 0.980 ;
        RECT 224.260 0.270 225.160 0.980 ;
        RECT 226.100 0.270 227.000 0.980 ;
        RECT 227.940 0.270 228.840 0.980 ;
        RECT 229.780 0.270 230.680 0.980 ;
        RECT 231.620 0.270 232.980 0.980 ;
        RECT 233.920 0.270 234.820 0.980 ;
        RECT 235.760 0.270 236.660 0.980 ;
        RECT 237.600 0.270 238.500 0.980 ;
        RECT 239.440 0.270 240.340 0.980 ;
        RECT 241.280 0.270 242.640 0.980 ;
        RECT 243.580 0.270 243.640 0.980 ;
      LAYER met3 ;
        RECT 8.345 2.215 240.515 176.965 ;
      LAYER met4 ;
        RECT 107.935 4.800 173.780 103.865 ;
        RECT 176.180 4.800 177.080 103.865 ;
        RECT 179.480 4.800 192.905 103.865 ;
        RECT 107.935 2.215 192.905 4.800 ;
  END
END N_term_single
END LIBRARY

