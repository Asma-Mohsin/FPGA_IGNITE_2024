VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO N_term_single
  CLASS BLOCK ;
  FOREIGN N_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 231.000 BY 218.000 ;
  PIN Ci
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.260 0.000 95.640 0.700 ;
    END
  END Ci
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 188.180 0.000 188.560 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 206.120 0.000 206.500 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 207.960 0.000 208.340 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 209.340 0.000 209.720 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 211.180 0.000 211.560 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 213.020 0.000 213.400 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 214.860 0.000 215.240 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 216.700 0.000 217.080 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 218.080 0.000 218.460 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 219.920 0.000 220.300 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 221.760 0.000 222.140 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 190.020 0.000 190.400 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.860 0.000 192.240 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 193.700 0.000 194.080 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.540 0.000 195.920 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 197.380 0.000 197.760 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 198.760 0.000 199.140 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 200.600 0.000 200.980 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 202.440 0.000 202.820 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 204.280 0.000 204.660 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 5.560 217.300 5.940 218.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 42.820 217.300 43.200 218.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.500 217.300 46.880 218.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.180 217.300 50.560 218.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.860 217.300 54.240 218.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 57.540 217.300 57.920 218.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.220 217.300 61.600 218.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.900 217.300 65.280 218.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 68.580 217.300 68.960 218.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 72.720 217.300 73.100 218.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.400 217.300 76.780 218.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.240 217.300 9.620 218.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 12.920 217.300 13.300 218.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 16.600 217.300 16.980 218.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 20.280 217.300 20.660 218.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 23.960 217.300 24.340 218.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 27.640 217.300 28.020 218.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 31.780 217.300 32.160 218.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.460 217.300 35.840 218.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.140 217.300 39.520 218.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 3.720 0.000 4.100 0.700 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 5.560 0.000 5.940 0.700 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.940 0.000 7.320 0.700 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 8.780 0.000 9.160 0.700 ;
    END
  END N1END[3]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 24.880 0.000 25.260 0.700 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 26.260 0.000 26.640 0.700 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 28.100 0.000 28.480 0.700 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.940 0.000 30.320 0.700 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.780 0.000 32.160 0.700 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 33.620 0.000 34.000 0.700 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.460 0.000 35.840 0.700 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 36.840 0.000 37.220 0.700 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 10.620 0.000 11.000 0.700 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.460 0.000 12.840 0.700 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 14.300 0.000 14.680 0.700 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 15.680 0.000 16.060 0.700 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 17.520 0.000 17.900 0.700 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 19.360 0.000 19.740 0.700 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 21.200 0.000 21.580 0.700 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 23.040 0.000 23.420 0.700 ;
    END
  END N2MID[7]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.680 0.000 39.060 0.700 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.160 0.000 56.540 0.700 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.000 0.000 58.380 0.700 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.840 0.000 60.220 0.700 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.680 0.000 62.060 0.700 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.520 0.000 63.900 0.700 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.360 0.000 65.740 0.700 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 40.520 0.000 40.900 0.700 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 42.360 0.000 42.740 0.700 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 44.200 0.000 44.580 0.700 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 46.040 0.000 46.420 0.700 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 47.420 0.000 47.800 0.700 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 49.260 0.000 49.640 0.700 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.100 0.000 51.480 0.700 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 52.940 0.000 53.320 0.700 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.780 0.000 55.160 0.700 ;
    END
  END N4END[9]
  PIN NN4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 66.740 0.000 67.120 0.700 ;
    END
  END NN4END[0]
  PIN NN4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.680 0.000 85.060 0.700 ;
    END
  END NN4END[10]
  PIN NN4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 86.520 0.000 86.900 0.700 ;
    END
  END NN4END[11]
  PIN NN4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.900 0.000 88.280 0.700 ;
    END
  END NN4END[12]
  PIN NN4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 89.740 0.000 90.120 0.700 ;
    END
  END NN4END[13]
  PIN NN4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 91.580 0.000 91.960 0.700 ;
    END
  END NN4END[14]
  PIN NN4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 93.420 0.000 93.800 0.700 ;
    END
  END NN4END[15]
  PIN NN4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 68.580 0.000 68.960 0.700 ;
    END
  END NN4END[1]
  PIN NN4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 70.420 0.000 70.800 0.700 ;
    END
  END NN4END[2]
  PIN NN4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 72.260 0.000 72.640 0.700 ;
    END
  END NN4END[3]
  PIN NN4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.100 0.000 74.480 0.700 ;
    END
  END NN4END[4]
  PIN NN4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 75.940 0.000 76.320 0.700 ;
    END
  END NN4END[5]
  PIN NN4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.320 0.000 77.700 0.700 ;
    END
  END NN4END[6]
  PIN NN4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 79.160 0.000 79.540 0.700 ;
    END
  END NN4END[7]
  PIN NN4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.000 0.000 81.380 0.700 ;
    END
  END NN4END[8]
  PIN NN4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.840 0.000 83.220 0.700 ;
    END
  END NN4END[9]
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.640 0.000 97.020 0.700 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.480 0.000 98.860 0.700 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 100.320 0.000 100.700 0.700 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.160 0.000 102.540 0.700 ;
    END
  END S1BEG[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.000 0.000 104.380 0.700 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.840 0.000 106.220 0.700 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.220 0.000 107.600 0.700 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.060 0.000 109.440 0.700 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.900 0.000 111.280 0.700 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.740 0.000 113.120 0.700 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.580 0.000 114.960 0.700 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.420 0.000 116.800 0.700 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.800 0.000 118.180 0.700 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.640 0.000 120.020 0.700 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.480 0.000 121.860 0.700 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 123.320 0.000 123.700 0.700 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.160 0.000 125.540 0.700 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.000 0.000 127.380 0.700 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.380 0.000 128.760 0.700 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.220 0.000 130.600 0.700 ;
    END
  END S2BEGb[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.060 0.000 132.440 0.700 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.540 0.000 149.920 0.700 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.380 0.000 151.760 0.700 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 153.220 0.000 153.600 0.700 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.060 0.000 155.440 0.700 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.900 0.000 157.280 0.700 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 158.280 0.000 158.660 0.700 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.900 0.000 134.280 0.700 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.740 0.000 136.120 0.700 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 137.120 0.000 137.500 0.700 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.960 0.000 139.340 0.700 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.800 0.000 141.180 0.700 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.640 0.000 143.020 0.700 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.480 0.000 144.860 0.700 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 0.000 146.700 0.700 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 147.700 0.000 148.080 0.700 ;
    END
  END S4BEG[9]
  PIN SS4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.120 0.000 160.500 0.700 ;
    END
  END SS4BEG[0]
  PIN SS4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 177.600 0.000 177.980 0.700 ;
    END
  END SS4BEG[10]
  PIN SS4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 179.440 0.000 179.820 0.700 ;
    END
  END SS4BEG[11]
  PIN SS4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 181.280 0.000 181.660 0.700 ;
    END
  END SS4BEG[12]
  PIN SS4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 183.120 0.000 183.500 0.700 ;
    END
  END SS4BEG[13]
  PIN SS4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 184.960 0.000 185.340 0.700 ;
    END
  END SS4BEG[14]
  PIN SS4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 186.800 0.000 187.180 0.700 ;
    END
  END SS4BEG[15]
  PIN SS4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.960 0.000 162.340 0.700 ;
    END
  END SS4BEG[1]
  PIN SS4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 163.800 0.000 164.180 0.700 ;
    END
  END SS4BEG[2]
  PIN SS4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.640 0.000 166.020 0.700 ;
    END
  END SS4BEG[3]
  PIN SS4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.480 0.000 167.860 0.700 ;
    END
  END SS4BEG[4]
  PIN SS4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 168.860 0.000 169.240 0.700 ;
    END
  END SS4BEG[5]
  PIN SS4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 170.700 0.000 171.080 0.700 ;
    END
  END SS4BEG[6]
  PIN SS4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 172.540 0.000 172.920 0.700 ;
    END
  END SS4BEG[7]
  PIN SS4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 174.380 0.000 174.760 0.700 ;
    END
  END SS4BEG[8]
  PIN SS4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 176.220 0.000 176.600 0.700 ;
    END
  END SS4BEG[9]
  PIN UIO_TOP_UIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 154.140 217.300 154.520 218.000 ;
    END
  END UIO_TOP_UIN0
  PIN UIO_TOP_UIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 158.280 217.300 158.660 218.000 ;
    END
  END UIO_TOP_UIN1
  PIN UIO_TOP_UIN10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.960 217.300 162.340 218.000 ;
    END
  END UIO_TOP_UIN10
  PIN UIO_TOP_UIN11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.640 217.300 166.020 218.000 ;
    END
  END UIO_TOP_UIN11
  PIN UIO_TOP_UIN12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 169.320 217.300 169.700 218.000 ;
    END
  END UIO_TOP_UIN12
  PIN UIO_TOP_UIN13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.000 217.300 173.380 218.000 ;
    END
  END UIO_TOP_UIN13
  PIN UIO_TOP_UIN14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 176.680 217.300 177.060 218.000 ;
    END
  END UIO_TOP_UIN14
  PIN UIO_TOP_UIN15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.360 217.300 180.740 218.000 ;
    END
  END UIO_TOP_UIN15
  PIN UIO_TOP_UIN16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 184.040 217.300 184.420 218.000 ;
    END
  END UIO_TOP_UIN16
  PIN UIO_TOP_UIN17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 187.720 217.300 188.100 218.000 ;
    END
  END UIO_TOP_UIN17
  PIN UIO_TOP_UIN18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.400 217.300 191.780 218.000 ;
    END
  END UIO_TOP_UIN18
  PIN UIO_TOP_UIN19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 195.080 217.300 195.460 218.000 ;
    END
  END UIO_TOP_UIN19
  PIN UIO_TOP_UIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 198.760 217.300 199.140 218.000 ;
    END
  END UIO_TOP_UIN2
  PIN UIO_TOP_UIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 202.900 217.300 203.280 218.000 ;
    END
  END UIO_TOP_UIN3
  PIN UIO_TOP_UIN4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.580 217.300 206.960 218.000 ;
    END
  END UIO_TOP_UIN4
  PIN UIO_TOP_UIN5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 210.260 217.300 210.640 218.000 ;
    END
  END UIO_TOP_UIN5
  PIN UIO_TOP_UIN6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 213.940 217.300 214.320 218.000 ;
    END
  END UIO_TOP_UIN6
  PIN UIO_TOP_UIN7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.620 217.300 218.000 218.000 ;
    END
  END UIO_TOP_UIN7
  PIN UIO_TOP_UIN8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 221.300 217.300 221.680 218.000 ;
    END
  END UIO_TOP_UIN8
  PIN UIO_TOP_UIN9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 224.980 217.300 225.360 218.000 ;
    END
  END UIO_TOP_UIN9
  PIN UIO_TOP_UOUT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.080 217.300 80.460 218.000 ;
    END
  END UIO_TOP_UOUT0
  PIN UIO_TOP_UOUT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.760 217.300 84.140 218.000 ;
    END
  END UIO_TOP_UOUT1
  PIN UIO_TOP_UOUT10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.440 217.300 87.820 218.000 ;
    END
  END UIO_TOP_UOUT10
  PIN UIO_TOP_UOUT11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.120 217.300 91.500 218.000 ;
    END
  END UIO_TOP_UOUT11
  PIN UIO_TOP_UOUT12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.800 217.300 95.180 218.000 ;
    END
  END UIO_TOP_UOUT12
  PIN UIO_TOP_UOUT13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.480 217.300 98.860 218.000 ;
    END
  END UIO_TOP_UOUT13
  PIN UIO_TOP_UOUT14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.160 217.300 102.540 218.000 ;
    END
  END UIO_TOP_UOUT14
  PIN UIO_TOP_UOUT15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.840 217.300 106.220 218.000 ;
    END
  END UIO_TOP_UOUT15
  PIN UIO_TOP_UOUT16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.520 217.300 109.900 218.000 ;
    END
  END UIO_TOP_UOUT16
  PIN UIO_TOP_UOUT17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.200 217.300 113.580 218.000 ;
    END
  END UIO_TOP_UOUT17
  PIN UIO_TOP_UOUT18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.340 217.300 117.720 218.000 ;
    END
  END UIO_TOP_UOUT18
  PIN UIO_TOP_UOUT19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.020 217.300 121.400 218.000 ;
    END
  END UIO_TOP_UOUT19
  PIN UIO_TOP_UOUT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.700 217.300 125.080 218.000 ;
    END
  END UIO_TOP_UOUT2
  PIN UIO_TOP_UOUT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.380 217.300 128.760 218.000 ;
    END
  END UIO_TOP_UOUT3
  PIN UIO_TOP_UOUT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.060 217.300 132.440 218.000 ;
    END
  END UIO_TOP_UOUT4
  PIN UIO_TOP_UOUT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.740 217.300 136.120 218.000 ;
    END
  END UIO_TOP_UOUT5
  PIN UIO_TOP_UOUT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.420 217.300 139.800 218.000 ;
    END
  END UIO_TOP_UOUT6
  PIN UIO_TOP_UOUT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.100 217.300 143.480 218.000 ;
    END
  END UIO_TOP_UOUT7
  PIN UIO_TOP_UOUT8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.780 217.300 147.160 218.000 ;
    END
  END UIO_TOP_UOUT8
  PIN UIO_TOP_UOUT9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.460 217.300 150.840 218.000 ;
    END
  END UIO_TOP_UOUT9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 230.300 95.240 231.000 95.840 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 230.300 98.640 231.000 99.240 ;
    END
  END UserCLKo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -12.040 -11.660 -8.940 229.260 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 -11.660 242.960 -8.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 226.160 242.960 229.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.860 -11.660 242.960 229.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.580 -16.460 22.180 234.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 -16.460 175.780 234.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 21.290 247.760 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 174.470 247.760 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.840 -16.460 -13.740 234.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 -16.460 247.760 -13.360 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 230.960 247.760 234.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.660 -16.460 247.760 234.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.880 -16.460 25.480 234.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.480 -16.460 179.080 234.060 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 24.590 247.760 26.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 177.770 247.760 179.370 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 4.870 5.355 226.050 212.245 ;
      LAYER li1 ;
        RECT 5.060 5.355 225.860 212.245 ;
      LAYER met1 ;
        RECT 3.750 1.400 225.860 212.400 ;
      LAYER met2 ;
        RECT 3.780 217.020 5.280 217.300 ;
        RECT 6.220 217.020 8.960 217.300 ;
        RECT 9.900 217.020 12.640 217.300 ;
        RECT 13.580 217.020 16.320 217.300 ;
        RECT 17.260 217.020 20.000 217.300 ;
        RECT 20.940 217.020 23.680 217.300 ;
        RECT 24.620 217.020 27.360 217.300 ;
        RECT 28.300 217.020 31.500 217.300 ;
        RECT 32.440 217.020 35.180 217.300 ;
        RECT 36.120 217.020 38.860 217.300 ;
        RECT 39.800 217.020 42.540 217.300 ;
        RECT 43.480 217.020 46.220 217.300 ;
        RECT 47.160 217.020 49.900 217.300 ;
        RECT 50.840 217.020 53.580 217.300 ;
        RECT 54.520 217.020 57.260 217.300 ;
        RECT 58.200 217.020 60.940 217.300 ;
        RECT 61.880 217.020 64.620 217.300 ;
        RECT 65.560 217.020 68.300 217.300 ;
        RECT 69.240 217.020 72.440 217.300 ;
        RECT 73.380 217.020 76.120 217.300 ;
        RECT 77.060 217.020 79.800 217.300 ;
        RECT 80.740 217.020 83.480 217.300 ;
        RECT 84.420 217.020 87.160 217.300 ;
        RECT 88.100 217.020 90.840 217.300 ;
        RECT 91.780 217.020 94.520 217.300 ;
        RECT 95.460 217.020 98.200 217.300 ;
        RECT 99.140 217.020 101.880 217.300 ;
        RECT 102.820 217.020 105.560 217.300 ;
        RECT 106.500 217.020 109.240 217.300 ;
        RECT 110.180 217.020 112.920 217.300 ;
        RECT 113.860 217.020 117.060 217.300 ;
        RECT 118.000 217.020 120.740 217.300 ;
        RECT 121.680 217.020 124.420 217.300 ;
        RECT 125.360 217.020 128.100 217.300 ;
        RECT 129.040 217.020 131.780 217.300 ;
        RECT 132.720 217.020 135.460 217.300 ;
        RECT 136.400 217.020 139.140 217.300 ;
        RECT 140.080 217.020 142.820 217.300 ;
        RECT 143.760 217.020 146.500 217.300 ;
        RECT 147.440 217.020 150.180 217.300 ;
        RECT 151.120 217.020 153.860 217.300 ;
        RECT 154.800 217.020 158.000 217.300 ;
        RECT 158.940 217.020 161.680 217.300 ;
        RECT 162.620 217.020 165.360 217.300 ;
        RECT 166.300 217.020 169.040 217.300 ;
        RECT 169.980 217.020 172.720 217.300 ;
        RECT 173.660 217.020 176.400 217.300 ;
        RECT 177.340 217.020 180.080 217.300 ;
        RECT 181.020 217.020 183.760 217.300 ;
        RECT 184.700 217.020 187.440 217.300 ;
        RECT 188.380 217.020 191.120 217.300 ;
        RECT 192.060 217.020 194.800 217.300 ;
        RECT 195.740 217.020 198.480 217.300 ;
        RECT 199.420 217.020 202.620 217.300 ;
        RECT 203.560 217.020 206.300 217.300 ;
        RECT 207.240 217.020 209.980 217.300 ;
        RECT 210.920 217.020 213.660 217.300 ;
        RECT 214.600 217.020 217.340 217.300 ;
        RECT 218.280 217.020 221.020 217.300 ;
        RECT 221.960 217.020 224.700 217.300 ;
        RECT 3.780 0.980 225.300 217.020 ;
        RECT 4.380 0.270 5.280 0.980 ;
        RECT 6.220 0.270 6.660 0.980 ;
        RECT 7.600 0.270 8.500 0.980 ;
        RECT 9.440 0.270 10.340 0.980 ;
        RECT 11.280 0.270 12.180 0.980 ;
        RECT 13.120 0.270 14.020 0.980 ;
        RECT 14.960 0.270 15.400 0.980 ;
        RECT 16.340 0.270 17.240 0.980 ;
        RECT 18.180 0.270 19.080 0.980 ;
        RECT 20.020 0.270 20.920 0.980 ;
        RECT 21.860 0.270 22.760 0.980 ;
        RECT 23.700 0.270 24.600 0.980 ;
        RECT 25.540 0.270 25.980 0.980 ;
        RECT 26.920 0.270 27.820 0.980 ;
        RECT 28.760 0.270 29.660 0.980 ;
        RECT 30.600 0.270 31.500 0.980 ;
        RECT 32.440 0.270 33.340 0.980 ;
        RECT 34.280 0.270 35.180 0.980 ;
        RECT 36.120 0.270 36.560 0.980 ;
        RECT 37.500 0.270 38.400 0.980 ;
        RECT 39.340 0.270 40.240 0.980 ;
        RECT 41.180 0.270 42.080 0.980 ;
        RECT 43.020 0.270 43.920 0.980 ;
        RECT 44.860 0.270 45.760 0.980 ;
        RECT 46.700 0.270 47.140 0.980 ;
        RECT 48.080 0.270 48.980 0.980 ;
        RECT 49.920 0.270 50.820 0.980 ;
        RECT 51.760 0.270 52.660 0.980 ;
        RECT 53.600 0.270 54.500 0.980 ;
        RECT 55.440 0.270 55.880 0.980 ;
        RECT 56.820 0.270 57.720 0.980 ;
        RECT 58.660 0.270 59.560 0.980 ;
        RECT 60.500 0.270 61.400 0.980 ;
        RECT 62.340 0.270 63.240 0.980 ;
        RECT 64.180 0.270 65.080 0.980 ;
        RECT 66.020 0.270 66.460 0.980 ;
        RECT 67.400 0.270 68.300 0.980 ;
        RECT 69.240 0.270 70.140 0.980 ;
        RECT 71.080 0.270 71.980 0.980 ;
        RECT 72.920 0.270 73.820 0.980 ;
        RECT 74.760 0.270 75.660 0.980 ;
        RECT 76.600 0.270 77.040 0.980 ;
        RECT 77.980 0.270 78.880 0.980 ;
        RECT 79.820 0.270 80.720 0.980 ;
        RECT 81.660 0.270 82.560 0.980 ;
        RECT 83.500 0.270 84.400 0.980 ;
        RECT 85.340 0.270 86.240 0.980 ;
        RECT 87.180 0.270 87.620 0.980 ;
        RECT 88.560 0.270 89.460 0.980 ;
        RECT 90.400 0.270 91.300 0.980 ;
        RECT 92.240 0.270 93.140 0.980 ;
        RECT 94.080 0.270 94.980 0.980 ;
        RECT 95.920 0.270 96.360 0.980 ;
        RECT 97.300 0.270 98.200 0.980 ;
        RECT 99.140 0.270 100.040 0.980 ;
        RECT 100.980 0.270 101.880 0.980 ;
        RECT 102.820 0.270 103.720 0.980 ;
        RECT 104.660 0.270 105.560 0.980 ;
        RECT 106.500 0.270 106.940 0.980 ;
        RECT 107.880 0.270 108.780 0.980 ;
        RECT 109.720 0.270 110.620 0.980 ;
        RECT 111.560 0.270 112.460 0.980 ;
        RECT 113.400 0.270 114.300 0.980 ;
        RECT 115.240 0.270 116.140 0.980 ;
        RECT 117.080 0.270 117.520 0.980 ;
        RECT 118.460 0.270 119.360 0.980 ;
        RECT 120.300 0.270 121.200 0.980 ;
        RECT 122.140 0.270 123.040 0.980 ;
        RECT 123.980 0.270 124.880 0.980 ;
        RECT 125.820 0.270 126.720 0.980 ;
        RECT 127.660 0.270 128.100 0.980 ;
        RECT 129.040 0.270 129.940 0.980 ;
        RECT 130.880 0.270 131.780 0.980 ;
        RECT 132.720 0.270 133.620 0.980 ;
        RECT 134.560 0.270 135.460 0.980 ;
        RECT 136.400 0.270 136.840 0.980 ;
        RECT 137.780 0.270 138.680 0.980 ;
        RECT 139.620 0.270 140.520 0.980 ;
        RECT 141.460 0.270 142.360 0.980 ;
        RECT 143.300 0.270 144.200 0.980 ;
        RECT 145.140 0.270 146.040 0.980 ;
        RECT 146.980 0.270 147.420 0.980 ;
        RECT 148.360 0.270 149.260 0.980 ;
        RECT 150.200 0.270 151.100 0.980 ;
        RECT 152.040 0.270 152.940 0.980 ;
        RECT 153.880 0.270 154.780 0.980 ;
        RECT 155.720 0.270 156.620 0.980 ;
        RECT 157.560 0.270 158.000 0.980 ;
        RECT 158.940 0.270 159.840 0.980 ;
        RECT 160.780 0.270 161.680 0.980 ;
        RECT 162.620 0.270 163.520 0.980 ;
        RECT 164.460 0.270 165.360 0.980 ;
        RECT 166.300 0.270 167.200 0.980 ;
        RECT 168.140 0.270 168.580 0.980 ;
        RECT 169.520 0.270 170.420 0.980 ;
        RECT 171.360 0.270 172.260 0.980 ;
        RECT 173.200 0.270 174.100 0.980 ;
        RECT 175.040 0.270 175.940 0.980 ;
        RECT 176.880 0.270 177.320 0.980 ;
        RECT 178.260 0.270 179.160 0.980 ;
        RECT 180.100 0.270 181.000 0.980 ;
        RECT 181.940 0.270 182.840 0.980 ;
        RECT 183.780 0.270 184.680 0.980 ;
        RECT 185.620 0.270 186.520 0.980 ;
        RECT 187.460 0.270 187.900 0.980 ;
        RECT 188.840 0.270 189.740 0.980 ;
        RECT 190.680 0.270 191.580 0.980 ;
        RECT 192.520 0.270 193.420 0.980 ;
        RECT 194.360 0.270 195.260 0.980 ;
        RECT 196.200 0.270 197.100 0.980 ;
        RECT 198.040 0.270 198.480 0.980 ;
        RECT 199.420 0.270 200.320 0.980 ;
        RECT 201.260 0.270 202.160 0.980 ;
        RECT 203.100 0.270 204.000 0.980 ;
        RECT 204.940 0.270 205.840 0.980 ;
        RECT 206.780 0.270 207.680 0.980 ;
        RECT 208.620 0.270 209.060 0.980 ;
        RECT 210.000 0.270 210.900 0.980 ;
        RECT 211.840 0.270 212.740 0.980 ;
        RECT 213.680 0.270 214.580 0.980 ;
        RECT 215.520 0.270 216.420 0.980 ;
        RECT 217.360 0.270 217.800 0.980 ;
        RECT 218.740 0.270 219.640 0.980 ;
        RECT 220.580 0.270 221.480 0.980 ;
        RECT 222.420 0.270 225.300 0.980 ;
      LAYER met3 ;
        RECT 5.585 99.640 230.300 212.325 ;
        RECT 5.585 98.240 229.900 99.640 ;
        RECT 5.585 96.240 230.300 98.240 ;
        RECT 5.585 94.840 229.900 96.240 ;
        RECT 5.585 5.275 230.300 94.840 ;
      LAYER met4 ;
        RECT 99.655 6.295 173.780 126.985 ;
        RECT 176.180 6.295 177.080 126.985 ;
        RECT 179.480 6.295 192.905 126.985 ;
  END
END N_term_single
END LIBRARY

