* NGSPICE file created from LUT4AB.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
XFILLER_0_76_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_11._0_ net144 VGND VGND VPWR VPWR NN4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_2
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LG_LUT4c_frame_config_dffesr.I0mux
+ Inst_LG_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_12._0_ strobe_inbuf_12.X VGND VGND VPWR VPWR strobe_outbuf_12.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst3 net509
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.ConfigBits\[502\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[503\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit16 net57 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit6 net78 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[372\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit27 net69 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_7._0_ data_inbuf_7.X VGND VGND VPWR VPWR data_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput401 net401 VGND VGND VPWR VPWR NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput434 net434 VGND VGND VPWR VPWR S4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput412 net412 VGND VGND VPWR VPWR S2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput423 net423 VGND VGND VPWR VPWR S2BEGb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_14_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput489 net489 VGND VGND VPWR VPWR W6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput456 net456 VGND VGND VPWR VPWR SS4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput445 net445 VGND VGND VPWR VPWR SS4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput467 net467 VGND VGND VPWR VPWR W2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput478 net478 VGND VGND VPWR VPWR W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst0._0__530 VGND
+ VGND VPWR VPWR net530 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst0._0__530/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XWW4END_inbuf_3._0_ net251 VGND VGND VPWR VPWR WW4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LH_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LH_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit22 net64 net87 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[325\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._1_
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit11 net52 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[356\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit30 net73 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[608\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG3 net114 net14 net218 Inst_LUT4AB_switch_matrix.JW2BEG6
+ Inst_LUT4AB_ConfigMem.ConfigBits\[384\] Inst_LUT4AB_ConfigMem.ConfigBits\[385\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_51_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit9 net81 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[447\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput286 net286 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput275 net275 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput264 net264 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit15 net56 net90 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sCD._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._0_ sky130_fd_sc_hd__inv_2
Xoutput297 net297 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit26 net68 net90 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG1 net108 net8 net160 net246
+ Inst_LUT4AB_ConfigMem.ConfigBits\[428\] Inst_LUT4AB_ConfigMem.ConfigBits\[429\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_CD_BEG1 sky130_fd_sc_hd__mux4_2
X_200_ Inst_LUT4AB_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
X_131_ N4BEG_outbuf_11.X VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
X_062_ Inst_LUT4AB_switch_matrix.E2BEG6 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__buf_1
XFILLER_0_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix._072_ Inst_LUT4AB_switch_matrix.JS2BEG2 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit1 net61 net91 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[315\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst3 net535
+ net508 net511 Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.ConfigBits\[574\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[575\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit10 net51 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[406\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit21 net63 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[189\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG2 net541 Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1
+ Inst_LUT4AB_switch_matrix.JN2BEG1 Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[186\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[187\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LE_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LE_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XE6END_inbuf_3._0_ net29 VGND VGND VPWR VPWR E6BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ Inst_LUT4AB_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_1
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
X_045_ E6BEG_outbuf_5.X VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkbuf_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix._055_ Inst_LUT4AB_switch_matrix.JN2BEG1 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG1 sky130_fd_sc_hd__clkbuf_2
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AB._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN\[1\]
+ Inst_LUT4AB_switch_matrix.S0 VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[286\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._1_
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit14 net55 net89 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit25 net67 net89 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit22 net64 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[197\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit11 net52 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[419\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XSS4END_inbuf_5._0_ net205 VGND VGND VPWR VPWR SS4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit8 Inst_LUT4AB_switch_matrix.M_AB VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__buf_4
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit1 net61 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[397\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._107_ net509 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit4 net76 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[298\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
X_028_ data_outbuf_28.X VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit20 net62 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[191\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit31 net74 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[594\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._038_ net17 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb3
+ sky130_fd_sc_hd__clkbuf_2
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_7._0_ strobe_inbuf_7.X VGND VGND VPWR VPWR strobe_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit18 net59 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[154\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst3 net509
+ net541 net515 net542 Inst_LUT4AB_ConfigMem.ConfigBits\[538\] Inst_LUT4AB_ConfigMem.ConfigBits\[539\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst0._0_ net516 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst0 net105
+ net107 net129 net41 Inst_LUT4AB_ConfigMem.ConfigBits\[482\] Inst_LUT4AB_ConfigMem.ConfigBits\[483\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XEE4END_inbuf_4._0_ net48 VGND VGND VPWR VPWR EE4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_1._0_ net61 VGND VGND VPWR VPWR data_inbuf_1.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst1 net509 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ net538 Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[179\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[180\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
Xinput197 SS4END[1] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_2
Xinput186 S4END[6] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xinput164 S2END[6] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__buf_2
Xinput175 S4END[10] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst1 net537 net510
+ net509 net541 Inst_LUT4AB_ConfigMem.ConfigBits\[206\] Inst_LUT4AB_ConfigMem.ConfigBits\[207\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xinput153 NN4END[9] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
Xinput142 NN4END[13] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xinput120 N2MID[6] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_4
Xinput131 N4END[3] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit13 net54 net88 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit24 net66 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4BEG_outbuf_5._0_ WW4BEG_outbuf_5.A VGND VGND VPWR VPWR WW4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit7 net79 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[460\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LC_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit10 net51 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[538\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit21 net63 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[230\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst0._0__516 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst0._0__516/HI
+ net516 sky130_fd_sc_hd__conb_1
XInst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LG_LUT4c_frame_config_dffesr.I0mux
+ Inst_LG_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[254\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.WW4BEG2 sky130_fd_sc_hd__o21ai_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit30 net73 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[585\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[504\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[505\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG5
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit17 net58 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit28 net70 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit7 net79 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[401\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XE6BEG_outbuf_8._0_ E6BEG_outbuf_8.A VGND VGND VPWR VPWR E6BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[178\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.NN4BEG2 sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LA_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
Xoutput402 net402 VGND VGND VPWR VPWR NN4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput435 net435 VGND VGND VPWR VPWR S4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput457 net457 VGND VGND VPWR VPWR SS4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput413 net413 VGND VGND VPWR VPWR S2BEG[2] sky130_fd_sc_hd__clkbuf_4
XN4END_inbuf_7._0_ net124 VGND VGND VPWR VPWR N4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_2
Xoutput424 net424 VGND VGND VPWR VPWR S2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput446 net446 VGND VGND VPWR VPWR SS4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput468 net468 VGND VGND VPWR VPWR W2BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput479 net479 VGND VGND VPWR VPWR W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[198\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG2 sky130_fd_sc_hd__o21ai_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[325\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit23 net65 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[192\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit12 net53 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[344\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst0 net103
+ net109 net43 net25 Inst_LUT4AB_ConfigMem.ConfigBits\[554\] Inst_LUT4AB_ConfigMem.ConfigBits\[555\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit20 net62 net99 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit31 net74 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[596\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I0 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 Inst_LUT4AB_switch_matrix.J2END_AB_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[267\] Inst_LUT4AB_ConfigMem.ConfigBits\[268\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_59_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst0 net103 net3
+ net207 Inst_LD_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[235\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[236\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput254 net254 VGND VGND VPWR VPWR Co sky130_fd_sc_hd__buf_2
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput276 net276 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput298 net298 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput287 net287 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput265 net265 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit16 net57 net90 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit27 net69 net90 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
X_130_ N4BEG_outbuf_10.X VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG2 net110 net10 net198 net214
+ Inst_LUT4AB_ConfigMem.ConfigBits\[430\] Inst_LUT4AB_ConfigMem.ConfigBits\[431\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_CD_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_061_ Inst_LUT4AB_switch_matrix.E2BEG5 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._071_ Inst_LUT4AB_switch_matrix.JS2BEG1 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG1 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst0._0__525 VGND
+ VGND VPWR VPWR net525 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst0._0__525/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit2 net72 net91 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[314\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[576\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[577\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG7
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_62_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG3 net540 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2
+ Inst_LUT4AB_switch_matrix.JN2BEG2 Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[188\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[189\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit11 net52 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[393\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit22 net64 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[226\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LE_LUT4c_frame_config_dffesr._20_ Inst_LE_LUT4c_frame_config_dffesr._06_ Inst_LE_LUT4c_frame_config_dffesr._07_
+ Inst_LE_LUT4c_frame_config_dffesr._08_ Inst_LE_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit30 net73 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[606\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.break_comb_loop_inst0._0_ Inst_MUX8LUT_frame_config_mux.GH
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst0 net146
+ net2 net42 net22 Inst_LUT4AB_ConfigMem.ConfigBits\[518\] Inst_LUT4AB_ConfigMem.ConfigBits\[519\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix._054_ Inst_LUT4AB_switch_matrix.JN2BEG0 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG0 sky130_fd_sc_hd__clkbuf_1
X_113_ Inst_LUT4AB_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
X_044_ E6BEG_outbuf_4.X VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG0 net121 net21 net173 net225
+ Inst_LUT4AB_ConfigMem.ConfigBits\[394\] Inst_LUT4AB_ConfigMem.ConfigBits\[395\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 sky130_fd_sc_hd__mux4_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_AB._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit15 net56 net89 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[286\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit26 net68 net89 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XNN4BEG_outbuf_8._0_ NN4BEG_outbuf_8.A VGND VGND VPWR VPWR NN4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst0._0_ net525 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit12 net53 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[418\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit23 net65 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[195\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit9 Inst_LA_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__buf_4
Xdata_outbuf_10._0_ data_inbuf_10.X VGND VGND VPWR VPWR data_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit5 net77 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[309\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._106_ net510 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.D
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._037_ net16 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_027_ data_outbuf_27.X VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit10 net51 net85 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LF_LUT4c_frame_config_dffesr.I0mux
+ Inst_LF_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit21 net63 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[227\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit19 net60 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[239\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[540\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[541\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG6
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_8_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst1 net25 net159
+ net211 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[482\] Inst_LUT4AB_ConfigMem.ConfigBits\[483\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput110 N2END[4] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xinput198 SS4END[2] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_2
Xinput187 S4END[7] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xinput165 S2END[7] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__buf_2
Xinput154 S1END[0] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
Xinput176 S4END[11] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit25 net67 net88 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit14 net55 net88 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst2 net511 Inst_LH_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[206\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[207\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
Xinput132 N4END[4] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput121 N2MID[7] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_4
Xinput143 NN4END[14] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I0 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 Inst_LUT4AB_switch_matrix.J2END_CD_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[297\] Inst_LUT4AB_ConfigMem.ConfigBits\[298\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit8 net80 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[493\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit11 net52 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[520\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XW6END_inbuf_1._0_ net231 VGND VGND VPWR VPWR W6BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_5._0_ net153 VGND VGND VPWR VPWR NN4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit22 net64 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[219\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LG_LUT4c_frame_config_dffesr.I0mux
+ Inst_LG_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst0._0__529 VGND
+ VGND VPWR VPWR net529 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst0._0__529/LO
+ sky130_fd_sc_hd__conb_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[254\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit20 net62 net84 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit8 net80 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[408\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit31 net74 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[584\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit29 net71 net91 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit18 net59 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG0 net9 net199 net246 Inst_LUT4AB_switch_matrix.JN2BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[586\] Inst_LUT4AB_ConfigMem.ConfigBits\[587\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_31_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[178\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XWW4END_inbuf_11._0_ net244 VGND VGND VPWR VPWR WW4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput403 net403 VGND VGND VPWR VPWR NN4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput458 net458 VGND VGND VPWR VPWR SS4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput447 net447 VGND VGND VPWR VPWR SS4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput436 net436 VGND VGND VPWR VPWR S4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput414 net414 VGND VGND VPWR VPWR S2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput425 net425 VGND VGND VPWR VPWR S2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput469 net469 VGND VGND VPWR VPWR W2BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[198\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit13 net54 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[364\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst1 net183
+ net199 net213 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[554\] Inst_LUT4AB_ConfigMem.ConfigBits\[555\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit24 net66 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[183\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit21 net63 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[172\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit10 net51 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[512\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LF_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LF_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I1 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 Inst_LUT4AB_switch_matrix.J2END_AB_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[269\] Inst_LUT4AB_ConfigMem.ConfigBits\[270\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_59_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst1 net535 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ net539 Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[235\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[236\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput277 net277 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput299 net299 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput266 net266 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput255 net255 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit30 net73 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[615\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit17 net58 net90 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit28 net70 net90 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst0 net103
+ net111 net3 net11 Inst_LUT4AB_ConfigMem.ConfigBits\[466\] Inst_LUT4AB_ConfigMem.ConfigBits\[467\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix._070_ Inst_LUT4AB_switch_matrix.JS2BEG0 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG0 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG3 net106 net41 net158 net210
+ Inst_LUT4AB_ConfigMem.ConfigBits\[432\] Inst_LUT4AB_ConfigMem.ConfigBits\[433\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_CD_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_18_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_060_ Inst_LUT4AB_switch_matrix.E2BEG4 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG0 net120 net172 net224
+ Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[354\] Inst_LUT4AB_ConfigMem.ConfigBits\[355\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit3 net75 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_189_ SS4BEG_outbuf_1.X VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit23 net65 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[267\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit12 net53 net86 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XFILLER_0_2_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit20 net62 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[170\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit31 net74 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[605\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst1 net182
+ net198 net212 net226 Inst_LUT4AB_ConfigMem.ConfigBits\[518\] Inst_LUT4AB_ConfigMem.ConfigBits\[519\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
X_112_ Inst_LUT4AB_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_30._0_ net73 VGND VGND VPWR VPWR data_inbuf_30.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._053_ Inst_LG_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LH_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__clkbuf_1
X_043_ E6BEG_outbuf_3.X VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_1
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG1 net117 net17 net169 net221
+ Inst_LUT4AB_ConfigMem.ConfigBits\[396\] Inst_LUT4AB_ConfigMem.ConfigBits\[397\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_inbuf_21._0_ net63 VGND VGND VPWR VPWR data_inbuf_21.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I0 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 Inst_LUT4AB_switch_matrix.J2END_GH_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[327\] Inst_LUT4AB_ConfigMem.ConfigBits\[328\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit16 net57 net89 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit27 net69 net89 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit13 net54 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[414\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst0._0_ net521 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit24 net66 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[218\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_0._0_ net82 VGND VGND VPWR VPWR strobe_inbuf_0.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_12._0_ net53 VGND VGND VPWR VPWR data_inbuf_12.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit3 net75 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[413\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit6 net78 net88 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._105_ Inst_LH_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR net254 sky130_fd_sc_hd__clkbuf_1
X_026_ data_outbuf_26.X VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LF_LUT4c_frame_config_dffesr.I0mux
+ Inst_LF_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix._036_ net15 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb1
+ sky130_fd_sc_hd__buf_1
XANTENNA_7 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit22 net64 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[225\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit11 net52 net85 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst2 Inst_LB_LUT4c_frame_config_dffesr.O
+ net512 Inst_LD_LUT4c_frame_config_dffesr.O Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[482\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[483\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit30 net73 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[210\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 FrameStrobe[8] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_16
Xinput111 N2END[5] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
Xinput133 N4END[5] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput122 N4END[0] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__buf_2
Xinput144 NN4END[15] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput199 SS4END[3] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_2
Xinput188 S4END[8] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
Xinput166 S2MID[0] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__buf_2
Xinput155 S1END[1] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xinput177 S4END[12] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit15 net56 net88 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ net538 Inst_LUT4AB_ConfigMem.ConfigBits\[206\] Inst_LUT4AB_ConfigMem.ConfigBits\[207\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit26 net68 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[273\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_15._0_ strobe_inbuf_15.X VGND VGND VPWR VPWR strobe_outbuf_15.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_009_ data_outbuf_9.X VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I1 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2END_CD_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[299\] Inst_LUT4AB_ConfigMem.ConfigBits\[300\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit9 net81 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[519\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit12 net53 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[580\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit23 net65 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[215\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LG_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LG_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XWW4END_inbuf_6._0_ net239 VGND VGND VPWR VPWR WW4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit21 net63 net84 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit10 net51 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[416\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit9 net81 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[392\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit19 net60 net91 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG1 net130 net8 net217 Inst_LUT4AB_switch_matrix.JE2BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[588\] Inst_LUT4AB_ConfigMem.ConfigBits\[589\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput404 net404 VGND VGND VPWR VPWR NN4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput459 net459 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
Xoutput437 net437 VGND VGND VPWR VPWR S4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput415 net415 VGND VGND VPWR VPWR S2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput426 net426 VGND VGND VPWR VPWR S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput448 net448 VGND VGND VPWR VPWR SS4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_sCD.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.S1
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.break_comb_loop_inst0._0_ Inst_MUX8LUT_frame_config_mux.EH_GH
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit25 net67 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[182\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit14 net55 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[399\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst2 net514
+ net513 net510 Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[554\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[555\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit11 net52 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[508\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit22 net64 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[171\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LF_LUT4c_frame_config_dffesr._20_ Inst_LF_LUT4c_frame_config_dffesr._06_ Inst_LF_LUT4c_frame_config_dffesr._07_
+ Inst_LF_LUT4c_frame_config_dffesr._08_ Inst_LF_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I2 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 Inst_LUT4AB_switch_matrix.J2END_AB_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[271\] Inst_LUT4AB_ConfigMem.ConfigBits\[272\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
XFILLER_0_59_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit20 net62 net83 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput278 net278 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__buf_2
XFILLER_0_49_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput289 net289 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit31 net74 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[601\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit29 net71 net90 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit18 net59 net90 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst1 net155
+ net163 net207 net209 Inst_LUT4AB_ConfigMem.ConfigBits\[466\] Inst_LUT4AB_ConfigMem.ConfigBits\[467\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xstrobe_inbuf_12._0_ net85 VGND VGND VPWR VPWR strobe_inbuf_12.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit1 net61 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[336\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG1 net16 net168 net220 Inst_LUT4AB_switch_matrix.JE2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[356\] Inst_LUT4AB_ConfigMem.ConfigBits\[357\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XE6END_inbuf_6._0_ net32 VGND VGND VPWR VPWR E6BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit4 net76 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_188_ SS4BEG_outbuf_0.X VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit24 net66 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[288\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit13 net54 net86 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst0 net105
+ net113 net5 net13 Inst_LUT4AB_ConfigMem.ConfigBits\[506\] Inst_LUT4AB_ConfigMem.ConfigBits\[507\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst0._0_ net530 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_AH.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.EH
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit21 net63 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[181\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit10 net51 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[484\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst2 net514
+ net512 net510 Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[518\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[519\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XSS4END_inbuf_8._0_ net193 VGND VGND VPWR VPWR SS4BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_1
X_111_ Inst_LUT4AB_switch_matrix.N2BEG7 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._052_ Inst_LF_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LG_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_042_ E6BEG_outbuf_2.X VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG2 net119 net19 net171 net223
+ Inst_LUT4AB_ConfigMem.ConfigBits\[398\] Inst_LUT4AB_ConfigMem.ConfigBits\[399\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I1 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_switch_matrix.J2END_GH_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[329\] Inst_LUT4AB_ConfigMem.ConfigBits\[330\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit17 net58 net89 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit28 net70 net89 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit14 net55 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[445\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit25 net67 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[237\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit4 net76 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[462\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._104_ Inst_LC_LUT4c_frame_config_dffesr.O VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.C sky130_fd_sc_hd__clkbuf_1
XEE4END_inbuf_7._0_ net36 VGND VGND VPWR VPWR EE4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit7 net79 net88 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit12 net53 net85 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
X_025_ data_outbuf_25.X VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
XANTENNA_8 Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata_inbuf_4._0_ net76 VGND VGND VPWR VPWR data_inbuf_4.X sky130_fd_sc_hd__clkbuf_1
XInst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LF_LUT4c_frame_config_dffesr.I0mux
+ Inst_LF_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix._035_ net14 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit23 net65 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[224\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XWW4BEG_outbuf_8._0_ WW4BEG_outbuf_8.A VGND VGND VPWR VPWR WW4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[482\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[483\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit20 net62 net97 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit31 net74 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[589\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LH_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput178 S4END[13] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xinput167 S2MID[1] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_4
Xinput156 S1END[2] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_4
Xinput123 N4END[10] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput134 N4END[6] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput112 N2END[6] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_2
Xinput101 FrameStrobe[9] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_16
Xinput145 NN4END[1] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
Xinput189 S4END[9] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[208\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[209\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E6BEG1
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit16 net57 net88 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit27 net69 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[268\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_008_ data_outbuf_8.X VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEH._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[153\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit13 net54 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[554\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I2 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 Inst_LUT4AB_switch_matrix.J2END_CD_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[301\] Inst_LUT4AB_ConfigMem.ConfigBits\[302\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[237\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.SS4BEG3 sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit24 net66 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[235\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LG_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LG_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit22 net64 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[198\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit11 net52 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[394\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG2 net145 net41 net181 Inst_LUT4AB_switch_matrix.JS2BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[590\] Inst_LUT4AB_ConfigMem.ConfigBits\[591\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit30 net73 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[216\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[275\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._1_
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput405 net405 VGND VGND VPWR VPWR NN4BEG[8] sky130_fd_sc_hd__buf_2
XN4BEG_outbuf_2._0_ N4BEG_outbuf_2.A VGND VGND VPWR VPWR N4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xoutput416 net416 VGND VGND VPWR VPWR S2BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput438 net438 VGND VGND VPWR VPWR S4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput449 net449 VGND VGND VPWR VPWR SS4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput427 net427 VGND VGND VPWR VPWR S4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4BEG_outbuf_1._0_ SS4BEG_outbuf_1.A VGND VGND VPWR VPWR SS4BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit15 net56 net87 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit26 net68 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[228\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst3 Inst_LF_LUT4c_frame_config_dffesr.O
+ net511 Inst_LH_LUT4c_frame_config_dffesr.O Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[554\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[555\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit23 net65 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[180\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit12 net53 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[488\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst0 net102
+ net106 net2 net6 Inst_LUT4AB_ConfigMem.ConfigBits\[542\] Inst_LUT4AB_ConfigMem.ConfigBits\[543\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LA_I3 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 Inst_LUT4AB_switch_matrix.J2END_AB_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[273\] Inst_LUT4AB_ConfigMem.ConfigBits\[274\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_1
XW6BEG_outbuf_2._0_ W6BEG_outbuf_2.A VGND VGND VPWR VPWR W6BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput268 net268 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput257 net257 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit21 net63 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[199\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput279 net279 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit19 net60 net90 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit10 net51 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[395\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst2 net514
+ Inst_LB_LUT4c_frame_config_dffesr.O net537 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[466\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[467\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEF.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.S2
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit2 net72 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[353\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG2 net118 net18 net222 Inst_LUT4AB_switch_matrix.JS2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[358\] Inst_LUT4AB_ConfigMem.ConfigBits\[359\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit5 net77 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_187_ Inst_LUT4AB_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_31._0_ data_inbuf_31.X VGND VGND VPWR VPWR data_outbuf_31.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit14 net55 net86 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit25 net67 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[287\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst1 net155
+ net157 net165 net209 Inst_LUT4AB_ConfigMem.ConfigBits\[506\] Inst_LUT4AB_ConfigMem.ConfigBits\[507\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit11 net52 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[456\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_22._0_ data_inbuf_22.X VGND VGND VPWR VPWR data_outbuf_22.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit22 net64 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[208\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LE_LUT4c_frame_config_dffesr.I0mux
+ Inst_LE_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst3 net508
+ net511 Inst_LH_LUT4c_frame_config_dffesr.O Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[518\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[519\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
X_110_ Inst_LUT4AB_switch_matrix.N2BEG6 VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_041_ E6BEG_outbuf_1.X VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._051_ Inst_LE_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LF_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG3 net115 net15 net167 net219
+ Inst_LUT4AB_ConfigMem.ConfigBits\[400\] Inst_LUT4AB_ConfigMem.ConfigBits\[401\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_18_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_13._0_ data_inbuf_13.X VGND VGND VPWR VPWR data_outbuf_13.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_2._0_ S4BEG_outbuf_2.A VGND VGND VPWR VPWR S4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I2 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 Inst_LUT4AB_switch_matrix.J2END_GH_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[331\] Inst_LUT4AB_ConfigMem.ConfigBits\[332\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
X_239_ WW4BEG_outbuf_3.X VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit18 net59 net89 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit29 net71 net89 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst0 net104 net156
+ net208 net508 Inst_LUT4AB_ConfigMem.ConfigBits\[246\] Inst_LUT4AB_ConfigMem.ConfigBits\[247\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit26 net68 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[245\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit15 net56 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[525\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit5 net77 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[481\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4END_inbuf_0._0_ net184 VGND VGND VPWR VPWR S4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._103_ net513 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.B
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit8 net80 net88 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_024_ data_outbuf_24.X VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit13 net54 net85 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LF_LUT4c_frame_config_dffesr.I0mux
+ Inst_LF_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix._034_ Inst_LUT4AB_switch_matrix.JE2BEG7 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG7 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit24 net66 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[223\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_9 Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[484\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[485\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit21 net63 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[177\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit10 net51 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[437\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XNN4END_inbuf_8._0_ net141 VGND VGND VPWR VPWR NN4BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_4
XEE4BEG_outbuf_1._0_ EE4BEG_outbuf_1.A VGND VGND VPWR VPWR EE4BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XW6END_inbuf_4._0_ net234 VGND VGND VPWR VPWR W6BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput179 S4END[14] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
Xinput168 S2MID[2] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__buf_2
Xinput157 S1END[3] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
Xinput135 N4END[7] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xinput102 N1END[0] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__buf_4
Xinput146 NN4END[2] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_1
Xinput124 N4END[11] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
Xinput113 N2END[7] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_4
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit28 net70 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[289\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit17 net58 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LD_I3 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 Inst_LUT4AB_switch_matrix.J2END_CD_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[303\] Inst_LUT4AB_ConfigMem.ConfigBits\[304\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit14 net55 net100 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
X_007_ data_outbuf_7.X VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[153\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit25 net67 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[244\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[237\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LG_LUT4c_frame_config_dffesr._20_ Inst_LG_LUT4c_frame_config_dffesr._06_ Inst_LG_LUT4c_frame_config_dffesr._07_
+ Inst_LG_LUT4c_frame_config_dffesr._08_ Inst_LG_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit12 net53 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[410\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit23 net65 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[188\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG3 net122 net190 net226 Inst_LUT4AB_switch_matrix.JW2BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[592\] Inst_LUT4AB_ConfigMem.ConfigBits\[593\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit0 net50 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[311\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit31 net74 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[604\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit20 net62 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[550\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[275\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput406 net406 VGND VGND VPWR VPWR NN4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_0_22_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput439 net439 VGND VGND VPWR VPWR S4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput428 net428 VGND VGND VPWR VPWR S4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput417 net417 VGND VGND VPWR VPWR S2BEG[6] sky130_fd_sc_hd__clkbuf_4
XInst_LA_LUT4c_frame_config_dffesr._19_ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LA_LUT4c_frame_config_dffesr.SR Inst_LA_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit0 net50 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[322\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit16 net57 net87 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit27 net69 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[272\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[556\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[557\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG2
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit13 net54 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[540\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4BEG_outbuf_11._0_ EE4BEG_outbuf_11.A VGND VGND VPWR VPWR EE4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit24 net66 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[217\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst1 net154
+ net158 net206 net208 Inst_LUT4AB_ConfigMem.ConfigBits\[542\] Inst_LUT4AB_ConfigMem.ConfigBits\[543\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst0 net102 net2
+ net154 net513 Inst_LUT4AB_ConfigMem.ConfigBits\[196\] Inst_LUT4AB_ConfigMem.ConfigBits\[197\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit11 net52 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[411\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput269 net269 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__buf_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_AH._4_ Inst_LUT4AB_switch_matrix.S3 Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._0_
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._1_ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.AH
+ sky130_fd_sc_hd__o21ai_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LC_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit22 net64 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[196\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst3 Inst_LF_LUT4c_frame_config_dffesr.O
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.ConfigBits\[466\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[467\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit30 net73 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[186\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit3 net75 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[349\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG3 net114 net14 net166 Inst_LUT4AB_switch_matrix.JW2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[360\] Inst_LUT4AB_ConfigMem.ConfigBits\[361\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_outbuf_0._0_ data_inbuf_0.X VGND VGND VPWR VPWR data_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit6 net78 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_68_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_186_ Inst_LUT4AB_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit15 net56 net86 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_24._0_ net66 VGND VGND VPWR VPWR data_inbuf_24.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit26 net68 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[277\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst2 net514
+ net513 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[506\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[507\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit23 net65 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[206\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit12 net53 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[492\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_3._0_ net95 VGND VGND VPWR VPWR strobe_inbuf_3.X sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LE_LUT4c_frame_config_dffesr.I0mux
+ Inst_LE_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[520\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[521\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_15._0_ net56 VGND VGND VPWR VPWR data_inbuf_15.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._050_ Inst_LD_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LE_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_040_ E6BEG_outbuf_0.X VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sGH.break_comb_loop_inst0._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit19 net60 net89 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
X_169_ Inst_LUT4AB_switch_matrix.S2BEGb5 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LG_I3 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 Inst_LUT4AB_switch_matrix.J2END_GH_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[333\] Inst_LUT4AB_ConfigMem.ConfigBits\[334\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_2
X_238_ WW4BEG_outbuf_2.X VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst1 net540 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2END_GH_BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[246\] Inst_LUT4AB_ConfigMem.ConfigBits\[247\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit27 net69 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[292\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit16 net57 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[524\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit6 net78 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[473\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LH_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LH_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
X_023_ data_outbuf_23.X VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._033_ Inst_LUT4AB_switch_matrix.JE2BEG6 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG6 sky130_fd_sc_hd__buf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._102_ net514 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.A
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit9 net81 net88 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit14 net55 net85 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LF_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LF_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit25 net67 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[269\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_outbuf_18._0_ strobe_inbuf_18.X VGND VGND VPWR VPWR strobe_outbuf_18.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit22 net64 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[175\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit11 net52 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[436\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput169 S2MID[3] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
Xinput158 S2END[0] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_4
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit18 net59 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4END_inbuf_9._0_ net242 VGND VGND VPWR VPWR WW4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_1
Xinput136 N4END[8] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
Xinput114 N2MID[0] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_4
Xinput125 N4END[12] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_1
Xinput103 N1END[1] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__buf_4
Xinput147 NN4END[3] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit29 net71 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[282\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
X_006_ data_outbuf_6.X VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit26 net68 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[290\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit15 net56 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[161\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit13 net54 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[403\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit24 net66 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[187\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit1 net61 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[347\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit10 net51 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[486\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit21 net63 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[549\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_0._0_ strobe_inbuf_0.X VGND VGND VPWR VPWR strobe_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[251\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.WW4BEG1 sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput429 net429 VGND VGND VPWR VPWR S4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput418 net418 VGND VGND VPWR VPWR S2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput407 net407 VGND VGND VPWR VPWR S1BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LA_LUT4c_frame_config_dffesr._18_ Inst_LA_LUT4c_frame_config_dffesr.SR Inst_LA_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit1 net61 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[318\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit17 net58 net87 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit28 net70 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[293\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[175\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.NN4BEG1 sky130_fd_sc_hd__o21ai_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit14 net55 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[522\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit25 net67 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[236\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_15._0_ net88 VGND VGND VPWR VPWR strobe_inbuf_15.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.O
+ net532 net512 Inst_LD_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[542\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[543\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XE6END_inbuf_9._0_ net24 VGND VGND VPWR VPWR E6BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst1 net512 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_switch_matrix.J2END_CD_BEG0
+ Inst_LUT4AB_ConfigMem.ConfigBits\[196\] Inst_LUT4AB_ConfigMem.ConfigBits\[197\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AB.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.A
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[195\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG1 sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit12 net53 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[557\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput259 net259 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit23 net65 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[222\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XInst_MUX8LUT_frame_config_mux.cus_mux21_AH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN\[1\]
+ Inst_LUT4AB_switch_matrix.S3 VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[468\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[469\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG4
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_45_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit20 net62 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[500\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit31 net74 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[168\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit4 net76 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[367\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XE6BEG_outbuf_1._0_ E6BEG_outbuf_1.A VGND VGND VPWR VPWR E6BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit7 net79 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_185_ Inst_LUT4AB_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XN4END_inbuf_0._0_ net132 VGND VGND VPWR VPWR N4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit16 net57 net86 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit27 net69 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[276\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst3 net509
+ Inst_LF_LUT4c_frame_config_dffesr.O Inst_LH_LUT4c_frame_config_dffesr.O Inst_LUT4AB_switch_matrix.M_AD
+ Inst_LUT4AB_ConfigMem.ConfigBits\[506\] Inst_LUT4AB_ConfigMem.ConfigBits\[507\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit24 net66 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[204\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit13 net54 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[513\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LE_LUT4c_frame_config_dffesr.I0mux
+ Inst_LE_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG0 net512 Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3
+ Inst_LUT4AB_switch_matrix.JW2BEG3 Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[154\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[155\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[152\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_AD sky130_fd_sc_hd__o21ai_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[335\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._1_
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
Xdata_inbuf_7._0_ net79 VGND VGND VPWR VPWR data_inbuf_7.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_168_ Inst_LUT4AB_switch_matrix.S2BEGb4 VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_1
X_237_ WW4BEG_outbuf_1.X VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__clkbuf_1
X_099_ Inst_LUT4AB_switch_matrix.EE4BEG3 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit30 net73 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[265\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit17 net58 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[541\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit28 net70 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[281\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit7 net79 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[472\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LH_LUT4c_frame_config_dffesr._20_ Inst_LH_LUT4c_frame_config_dffesr._06_ Inst_LH_LUT4c_frame_config_dffesr._07_
+ Inst_LH_LUT4c_frame_config_dffesr._08_ Inst_LH_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
X_022_ data_outbuf_22.X VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._032_ Inst_LUT4AB_switch_matrix.JE2BEG5 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG5 sky130_fd_sc_hd__buf_1
XFILLER_0_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix._101_ net225 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb7
+ sky130_fd_sc_hd__buf_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit15 net56 net85 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit26 net68 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[266\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit23 net65 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[174\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit12 net53 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[458\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XFILLER_0_52_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput126 N4END[13] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_1
Xinput115 N2MID[1] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xinput104 N1END[2] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__buf_4
Xinput159 S2END[1] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit19 net60 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput148 NN4END[4] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput137 N4END[9] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
XInst_LB_LUT4c_frame_config_dffesr._19_ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LB_LUT4c_frame_config_dffesr.SR Inst_LB_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ data_outbuf_5.X VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit16 net57 net100 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit27 net69 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[286\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XNN4BEG_outbuf_1._0_ NN4BEG_outbuf_1.A VGND VGND VPWR VPWR NN4BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XN4BEG_outbuf_5._0_ N4BEG_outbuf_5.A VGND VGND VPWR VPWR N4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XSS4BEG_outbuf_4._0_ SS4BEG_outbuf_4.A VGND VGND VPWR VPWR SS4BEG_outbuf_4.X sky130_fd_sc_hd__buf_2
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[296\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._1_
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit25 net67 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[201\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit14 net55 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[521\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit2 net72 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[420\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit22 net64 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[532\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit11 net52 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[482\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[251\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput408 net408 VGND VGND VPWR VPWR S1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput419 net419 VGND VGND VPWR VPWR S2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XW6BEG_outbuf_5._0_ W6BEG_outbuf_5.A VGND VGND VPWR VPWR W6BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_2
XInst_LA_LUT4c_frame_config_dffesr._17_ Inst_LA_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit2 net72 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[296\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit18 net59 net87 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit29 net71 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[291\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[175\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit15 net56 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[582\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit26 net68 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[280\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst3 Inst_LE_LUT4c_frame_config_dffesr.O
+ net508 net511 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[542\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[543\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst0 net102
+ net108 net130 net8 Inst_LUT4AB_ConfigMem.ConfigBits\[486\] Inst_LUT4AB_ConfigMem.ConfigBits\[487\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LD_LUT4c_frame_config_dffesr.I0mux
+ Inst_LD_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[195\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit24 net66 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[221\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit13 net54 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[581\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AH._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit21 net63 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[547\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit10 net51 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[438\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit5 net77 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[431\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_25._0_ data_inbuf_25.X VGND VGND VPWR VPWR data_outbuf_25.X sky130_fd_sc_hd__clkbuf_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit8 net80 net91 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_184_ Inst_LUT4AB_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_16._0_ data_inbuf_16.X VGND VGND VPWR VPWR data_outbuf_16.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS4BEG_outbuf_5._0_ S4BEG_outbuf_5.A VGND VGND VPWR VPWR S4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit17 net58 net86 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit28 net70 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[592\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[508\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[509\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG6
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG1 net510 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0
+ Inst_LUT4AB_switch_matrix.JW2BEG0 Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[156\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[157\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_CD.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.C
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LE_LUT4c_frame_config_dffesr.I0mux
+ Inst_LE_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit25 net67 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[231\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit14 net55 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[490\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XS4END_inbuf_3._0_ net187 VGND VGND VPWR VPWR S4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[152\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[335\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._1_
+ sky130_fd_sc_hd__nand2_1
X_098_ Inst_LUT4AB_switch_matrix.EE4BEG2 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_167_ Inst_LUT4AB_switch_matrix.S2BEGb3 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_1
X_236_ WW4BEG_outbuf_0.X VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit20 net62 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[536\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit18 net59 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[556\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit31 net74 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[264\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit29 net71 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[591\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst0 net104
+ net110 net10 net22 Inst_LUT4AB_ConfigMem.ConfigBits\[558\] Inst_LUT4AB_ConfigMem.ConfigBits\[559\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit8 net80 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[502\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4BEG_outbuf_4._0_ EE4BEG_outbuf_4.A VGND VGND VPWR VPWR EE4BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XW6END_inbuf_7._0_ net237 VGND VGND VPWR VPWR W6BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._100_ net224 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
X_021_ data_outbuf_21.X VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit0 net50 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[354\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit16 net57 net85 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit27 net69 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[593\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit24 net66 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[173\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit13 net54 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[457\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_219_ Inst_LUT4AB_switch_matrix.W2BEGb3 VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit0 net50 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[305\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput149 NN4END[5] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xinput138 NN4END[0] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_1
Xinput127 N4END[14] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput116 N2MID[2] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_4
Xinput105 N1END[3] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__buf_4
XInst_LB_LUT4c_frame_config_dffesr._18_ Inst_LB_LUT4c_frame_config_dffesr.SR Inst_LB_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[612\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_SR_BEG0 sky130_fd_sc_hd__o21ai_4
X_004_ data_outbuf_4.X VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit17 net58 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[194\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit28 net70 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[607\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit30 net73 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[250\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst0 net147
+ net3 net9 net25 Inst_LUT4AB_ConfigMem.ConfigBits\[522\] Inst_LUT4AB_ConfigMem.ConfigBits\[523\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit15 net56 net84 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[296\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit26 net68 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[234\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit3 net75 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[433\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit12 net53 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[469\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEH.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.S1
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit23 net65 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[165\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput409 net409 VGND VGND VPWR VPWR S1BEG[2] sky130_fd_sc_hd__buf_2
XInst_LA_LUT4c_frame_config_dffesr._16_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit3 net75 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[332\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4END_inbuf_11._0_ net128 VGND VGND VPWR VPWR N4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit19 net60 net87 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSS4END_inbuf_10._0_ net195 VGND VGND VPWR VPWR SS4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit16 net57 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[555\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit27 net69 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[590\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_3._0_ data_inbuf_3.X VGND VGND VPWR VPWR data_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[544\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[545\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG7
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst1 net22 net160
+ net212 net247 Inst_LUT4AB_ConfigMem.ConfigBits\[486\] Inst_LUT4AB_ConfigMem.ConfigBits\[487\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LD_LUT4c_frame_config_dffesr.I0mux
+ Inst_LD_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit14 net55 net83 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit25 net67 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[220\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_27._0_ net69 VGND VGND VPWR VPWR data_inbuf_27.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit22 net64 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[546\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit11 net52 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[465\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit6 net78 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[430\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst0._0_ net517 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
Xstrobe_inbuf_6._0_ net98 VGND VGND VPWR VPWR strobe_inbuf_6.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_18._0_ net59 VGND VGND VPWR VPWR data_inbuf_18.X sky130_fd_sc_hd__clkbuf_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit9 net81 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_183_ S4BEG_outbuf_11.X VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit18 net59 net86 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit29 net71 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[613\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit15 net56 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[507\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG2 net509 Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1
+ Inst_LUT4AB_switch_matrix.JW2BEG1 Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[158\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[159\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_2
XInst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LE_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LE_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit26 net68 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[214\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_52_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_235_ Inst_LUT4AB_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkbuf_1
X_097_ Inst_LUT4AB_switch_matrix.EE4BEG1 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkbuf_1
X_166_ Inst_LUT4AB_switch_matrix.S2BEGb2 VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit21 net63 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[535\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LC_LUT4c_frame_config_dffesr._19_ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LC_LUT4c_frame_config_dffesr.SR Inst_LC_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit10 net51 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[483\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XS4END_inbuf_11._0_ net180 VGND VGND VPWR VPWR S4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit19 net60 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[583\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst1 net162
+ net174 net214 net246 Inst_LUT4AB_ConfigMem.ConfigBits\[558\] Inst_LUT4AB_ConfigMem.ConfigBits\[559\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit9 net81 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[558\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_MUX8LUT_frame_config_mux.cus_mux21_EF.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.E
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit17 net58 net85 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
X_020_ data_outbuf_20.X VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit1 net61 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[350\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit28 net70 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[587\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_149_ Inst_LUT4AB_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit25 net67 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[185\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit14 net55 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[516\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
X_218_ Inst_LUT4AB_switch_matrix.W2BEGb2 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst0 net104
+ net112 net4 net12 Inst_LUT4AB_ConfigMem.ConfigBits\[470\] Inst_LUT4AB_ConfigMem.ConfigBits\[471\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit1 net61 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[303\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSS4END_inbuf_1._0_ net201 VGND VGND VPWR VPWR SS4BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_1
XEE4END_inbuf_10._0_ net39 VGND VGND VPWR VPWR EE4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_2
Xinput139 NN4END[10] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xinput117 N2MID[3] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
Xinput128 N4END[15] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xinput106 N2END[0] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_4
XInst_LB_LUT4c_frame_config_dffesr._17_ Inst_LB_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[612\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_90 NN4BEG_outbuf_0.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit20 net62 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[572\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst0._0__522 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst0._0__522/HI
+ net522 sky130_fd_sc_hd__conb_1
X_003_ data_outbuf_3.X VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit18 net59 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[193\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit31 net74 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[249\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit29 net71 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[600\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_3._0_ strobe_inbuf_3.X VGND VGND VPWR VPWR strobe_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst1 net161
+ net183 net213 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[522\] Inst_LUT4AB_ConfigMem.ConfigBits\[523\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit16 net57 net84 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[234\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.SS4BEG2 sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit27 net69 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[233\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4END_inbuf_0._0_ net44 VGND VGND VPWR VPWR EE4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit4 net76 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[449\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit13 net54 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[468\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit24 net66 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[152\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_18._0_ net91 VGND VGND VPWR VPWR strobe_inbuf_18.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XWW4BEG_outbuf_1._0_ WW4BEG_outbuf_1.A VGND VGND VPWR VPWR WW4BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_2
XInst_LA_LUT4c_frame_config_dffesr._15_ Inst_LA_LUT4c_frame_config_dffesr._01_ Inst_LA_LUT4c_frame_config_dffesr._02_
+ Inst_LA_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit4 net76 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[331\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst0._0_ net526 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit17 net58 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[552\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit28 net70 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[588\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XE6BEG_outbuf_4._0_ E6BEG_outbuf_4.A VGND VGND VPWR VPWR E6BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst2 net543
+ net512 Inst_LD_LUT4c_frame_config_dffesr.O net535 Inst_LUT4AB_ConfigMem.ConfigBits\[486\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[487\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LD_LUT4c_frame_config_dffesr.I0mux
+ Inst_LD_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst0._0__531 VGND
+ VGND VPWR VPWR net531 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst0._0__531/LO
+ sky130_fd_sc_hd__conb_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit15 net56 net83 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit26 net68 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[200\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XN4END_inbuf_3._0_ net135 VGND VGND VPWR VPWR N4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit12 net53 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[477\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit23 net65 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[545\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG0 net108 net129 net25 net509 Inst_LUT4AB_ConfigMem.ConfigBits\[162\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[163\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit7 net79 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[451\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_251_ Inst_LUT4AB_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkbuf_1
X_182_ S4BEG_outbuf_10.X VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XFILLER_0_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit19 net60 net86 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit16 net57 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[553\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit27 net69 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[213\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N1BEG3 net541 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2
+ Inst_LUT4AB_switch_matrix.JW2BEG2 Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[160\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[161\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_73_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_234_ Inst_LUT4AB_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_1
X_165_ Inst_LUT4AB_switch_matrix.S2BEGb1 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr._18_ Inst_LC_LUT4c_frame_config_dffesr.SR Inst_LC_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
X_096_ Inst_LUT4AB_switch_matrix.EE4BEG0 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit11 net52 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[475\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit22 net64 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[531\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.O
+ Inst_LB_LUT4c_frame_config_dffesr.O net512 Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[558\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[559\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.break_comb_loop_inst0._0_ Inst_MUX8LUT_frame_config_mux.CD
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit2 net72 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[341\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit18 net59 net85 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit29 net71 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[612\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput390 net390 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ Inst_LUT4AB_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit26 net68 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[178\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit15 net56 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[511\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_217_ Inst_LUT4AB_switch_matrix.W2BEGb1 VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._089_ Inst_LUT4AB_switch_matrix.JW2BEG3 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG3 sky130_fd_sc_hd__clkbuf_1
X_079_ strobe_outbuf_15.X VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst1 net156
+ net164 net206 net208 Inst_LUT4AB_ConfigMem.ConfigBits\[470\] Inst_LUT4AB_ConfigMem.ConfigBits\[471\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4BEG_outbuf_4._0_ NN4BEG_outbuf_4.A VGND VGND VPWR VPWR NN4BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XN4BEG_outbuf_8._0_ N4BEG_outbuf_8.A VGND VGND VPWR VPWR N4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit2 net72 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[323\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XSS4BEG_outbuf_7._0_ SS4BEG_outbuf_7.A VGND VGND VPWR VPWR SS4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_2
Xinput107 N2END[1] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__buf_2
Xinput118 N2MID[4] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__buf_2
Xinput129 N4END[1] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__buf_2
XInst_LB_LUT4c_frame_config_dffesr._16_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XS4BEG_outbuf_11._0_ S4BEG_outbuf_11.A VGND VGND VPWR VPWR S4BEG_outbuf_11.X sky130_fd_sc_hd__buf_2
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XANTENNA_91 NN4BEG_outbuf_8.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit21 net63 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[571\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
X_002_ data_outbuf_2.X VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_80 net543 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit10 net51 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[526\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_GH.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.G
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit19 net60 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[209\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst0 net102
+ net106 net2 net6 Inst_LUT4AB_ConfigMem.ConfigBits\[510\] Inst_LUT4AB_ConfigMem.ConfigBits\[511\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.O
+ Inst_LB_LUT4c_frame_config_dffesr.O Inst_LD_LUT4c_frame_config_dffesr.O Inst_LE_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_ConfigMem.ConfigBits\[522\] Inst_LUT4AB_ConfigMem.ConfigBits\[523\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AD.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.CD
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XW6BEG_outbuf_8._0_ W6BEG_outbuf_8.A VGND VGND VPWR VPWR W6BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit17 net58 net84 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit28 net70 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[610\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[234\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LC_LUT4c_frame_config_dffesr.I0mux
+ Inst_LC_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit5 net77 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[425\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit14 net55 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[466\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit25 net67 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[176\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst0._0__517 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst0._0__517/HI
+ net517 sky130_fd_sc_hd__conb_1
XFILLER_0_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4END_inbuf_1._0_ net149 VGND VGND VPWR VPWR NN4BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_4
XInst_LA_LUT4c_frame_config_dffesr._14_ Inst_LA_LUT4c_frame_config_dffesr.I\[1\] Inst_LA_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LA_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LH_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit5 net77 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[355\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit20 net62 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[259\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit18 net59 net99 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst0._0_ net522 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit29 net71 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[609\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_28._0_ data_inbuf_28.X VGND VGND VPWR VPWR data_outbuf_28.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst3 net508
+ net511 Inst_LH_LUT4c_frame_config_dffesr.O net542 Inst_LUT4AB_ConfigMem.ConfigBits\[486\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[487\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LD_LUT4c_frame_config_dffesr.I0mux
+ Inst_LD_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit16 net57 net83 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_19._0_ data_inbuf_19.X VGND VGND VPWR VPWR data_outbuf_19.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LF_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit27 net69 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[232\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_8._0_ S4BEG_outbuf_8.A VGND VGND VPWR VPWR S4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit13 net54 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[476\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit24 net66 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[533\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit8 net80 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[450\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr._19_ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LD_LUT4c_frame_config_dffesr.SR Inst_LD_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG1 net109 net130 net22 net508 Inst_LUT4AB_ConfigMem.ConfigBits\[164\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[165\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG1
+ sky130_fd_sc_hd__mux4_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_250_ Inst_LUT4AB_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkbuf_1
X_181_ S4BEG_outbuf_9.X VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XS4END_inbuf_6._0_ net175 VGND VGND VPWR VPWR S4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[285\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._1_
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit17 net58 net98 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit28 net70 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[212\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst0._0__526 VGND
+ VGND VPWR VPWR net526 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst0._0__526/LO
+ sky130_fd_sc_hd__conb_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit0 net50 net90 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[304\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4BEG_outbuf_7._0_ EE4BEG_outbuf_7.A VGND VGND VPWR VPWR EE4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG0 net113 net42 net165 net217
+ Inst_LUT4AB_ConfigMem.ConfigBits\[434\] Inst_LUT4AB_ConfigMem.ConfigBits\[435\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 sky130_fd_sc_hd__mux4_2
X_095_ EE4BEG_outbuf_11.X VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_1
X_233_ W6BEG_outbuf_9.X VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_164_ Inst_LUT4AB_switch_matrix.S2BEGb0 VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr._17_ Inst_LC_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit12 net53 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[474\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit23 net65 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[561\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.ConfigBits\[558\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[559\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_MUX8LUT_frame_config_mux.cus_mux21_GH._4_ Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.GH sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit3 net75 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[328\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput391 net391 VGND VGND VPWR VPWR NN4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput380 net380 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit19 net60 net85 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit27 net69 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[205\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit16 net57 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[510\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
X_078_ strobe_outbuf_14.X VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__clkbuf_1
X_147_ NN4BEG_outbuf_11.X VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_216_ Inst_LUT4AB_switch_matrix.W2BEGb0 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._088_ Inst_LUT4AB_switch_matrix.JW2BEG2 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG2 sky130_fd_sc_hd__buf_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst2 net514
+ net532 net537 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[470\] Inst_LUT4AB_ConfigMem.ConfigBits\[471\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit3 net75 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[320\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_28_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 N2END[2] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_2
XFILLER_0_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LB_LUT4c_frame_config_dffesr._15_ Inst_LB_LUT4c_frame_config_dffesr._01_ Inst_LB_LUT4c_frame_config_dffesr._02_
+ Inst_LB_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
Xinput119 N2MID[5] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_4
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit22 net64 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[570\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
X_001_ data_outbuf_1.X VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_1
XANTENNA_81 E6BEG_outbuf_7.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_92 S4BEG_outbuf_4.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit11 net52 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[543\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_70 net224 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XNN4BEG_outbuf_11._0_ NN4BEG_outbuf_11.A VGND VGND VPWR VPWR NN4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst1 net154
+ net156 net190 net238 Inst_LUT4AB_ConfigMem.ConfigBits\[510\] Inst_LUT4AB_ConfigMem.ConfigBits\[511\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst3 net508
+ net511 Inst_LH_LUT4c_frame_config_dffesr.O Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.ConfigBits\[522\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[523\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_10._0_ net143 VGND VGND VPWR VPWR NN4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit18 net59 net84 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit29 net71 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[602\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit6 net78 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[424\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
Xinput90 FrameStrobe[17] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_8
XFILLER_0_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit26 net68 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[184\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LC_LUT4c_frame_config_dffesr.I0mux
+ Inst_LC_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit15 net56 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[517\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.break_comb_loop_inst0._0_ net531 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_54_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_11._0_ strobe_inbuf_11.X VGND VGND VPWR VPWR strobe_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_6._0_ data_inbuf_6.X VGND VGND VPWR VPWR data_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst0 net105 net157
+ net209 net514 Inst_LUT4AB_ConfigMem.ConfigBits\[249\] Inst_LUT4AB_ConfigMem.ConfigBits\[250\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux41_buf_inst0 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[610\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[611\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit6 net78 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[339\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit21 net63 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[248\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit10 net51 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[577\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit19 net60 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[160\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[248\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.WW4BEG0 sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XWW4END_inbuf_2._0_ net250 VGND VGND VPWR VPWR WW4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[488\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[489\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG1
+ sky130_fd_sc_hd__mux4_2
Xstrobe_inbuf_9._0_ net101 VGND VGND VPWR VPWR strobe_inbuf_9.X sky130_fd_sc_hd__clkbuf_1
XInst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LD_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LD_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[172\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.NN4BEG0 sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit17 net58 net83 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit28 net70 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[271\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LD_LUT4c_frame_config_dffesr._18_ Inst_LD_LUT4c_frame_config_dffesr.SR Inst_LD_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit25 net67 net95 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit9 net81 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[446\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit14 net55 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[497\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG2 net106 net131 net229 net540 Inst_LUT4AB_ConfigMem.ConfigBits\[166\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[167\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG2
+ sky130_fd_sc_hd__mux4_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[192\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG0 sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_180_ S4BEG_outbuf_8.X VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit18 net59 net98 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[285\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit29 net71 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[211\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit1 net61 net90 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[299\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XE6END_inbuf_2._0_ net28 VGND VGND VPWR VPWR E6BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG1 net109 net9 net161 net245
+ Inst_LUT4AB_ConfigMem.ConfigBits\[436\] Inst_LUT4AB_ConfigMem.ConfigBits\[437\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_EF_BEG1 sky130_fd_sc_hd__mux4_2
X_232_ W6BEG_outbuf_8.X VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_094_ EE4BEG_outbuf_10.X VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_1
X_163_ Inst_LUT4AB_switch_matrix.S2BEG7 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_1
XInst_LC_LUT4c_frame_config_dffesr._16_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit24 net66 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[564\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit13 net54 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[494\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[560\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[561\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG3
+ sky130_fd_sc_hd__mux4_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_GH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN\[1\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XSS4END_inbuf_4._0_ net204 VGND VGND VPWR VPWR SS4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit4 net76 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[368\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput392 net392 VGND VGND VPWR VPWR NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput381 net381 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__buf_2
Xoutput370 net370 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst0 net103 net3
+ net155 Inst_LD_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[199\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[200\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit17 net58 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[506\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit28 net70 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[229\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
X_215_ Inst_LUT4AB_switch_matrix.W2BEG7 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_1
X_146_ NN4BEG_outbuf_10.X VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
X_077_ strobe_outbuf_13.X VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst3 net509
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[470\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[471\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix._087_ Inst_LUT4AB_switch_matrix.JW2BEG1 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LE_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_6._0_ strobe_inbuf_6.X VGND VGND VPWR VPWR strobe_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit4 net76 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[316\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG0 net121 net21 net173 net225
+ Inst_LUT4AB_ConfigMem.ConfigBits\[402\] Inst_LUT4AB_ConfigMem.ConfigBits\[403\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput109 N2END[3] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
XInst_LB_LUT4c_frame_config_dffesr._14_ Inst_LB_LUT4c_frame_config_dffesr.I\[1\] Inst_LB_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LB_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XEE4END_inbuf_3._0_ net47 VGND VGND VPWR VPWR EE4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_000_ data_outbuf_0.X VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_0._0_ net50 VGND VGND VPWR VPWR data_inbuf_0.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit23 net65 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[569\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_82 EE4BEG_outbuf_1.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 net238 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit12 net53 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[542\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_93 SS4BEG_outbuf_5.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst2 net514
+ net513 net512 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[510\] Inst_LUT4AB_ConfigMem.ConfigBits\[511\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XWW4BEG_outbuf_4._0_ WW4BEG_outbuf_4.A VGND VGND VPWR VPWR WW4BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[524\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[525\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG2
+ sky130_fd_sc_hd__mux4_2
X_129_ N4BEG_outbuf_9.X VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LC_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit19 net60 net84 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput80 FrameData[8] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_8
Xinput91 FrameStrobe[18] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_8
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit7 net79 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[487\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LC_LUT4c_frame_config_dffesr.I0mux
+ Inst_LC_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit27 net69 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[179\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit16 net57 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[515\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst1 net515 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 Inst_LUT4AB_switch_matrix.J2END_EF_BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[249\] Inst_LUT4AB_ConfigMem.ConfigBits\[250\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XE6BEG_outbuf_7._0_ E6BEG_outbuf_7.A VGND VGND VPWR VPWR E6BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr._19_ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LE_LUT4c_frame_config_dffesr.SR Inst_LE_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_22_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr._12_ Inst_LA_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XFILLER_0_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix.JN2BEG1
+ Inst_LUT4AB_switch_matrix.JE2BEG1 Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_switch_matrix.JW2BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[610\] Inst_LUT4AB_ConfigMem.ConfigBits\[611\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit7 net79 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[387\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XN4END_inbuf_6._0_ net123 VGND VGND VPWR VPWR N4BEG_outbuf_6.A sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit22 net64 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[247\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit11 net52 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[576\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LD_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[248\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[172\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit18 net59 net83 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit29 net71 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[270\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit26 net68 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[166\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit15 net56 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[496\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr._17_ Inst_LD_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_N4BEG3 net107 net122 net226 net515 Inst_LUT4AB_ConfigMem.ConfigBits\[168\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[169\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N4BEG3
+ sky130_fd_sc_hd__mux4_2
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[192\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.GH
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit19 net60 net98 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit2 net72 net90 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[325\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst0 net107
+ net129 net5 net7 Inst_LUT4AB_ConfigMem.ConfigBits\[450\] Inst_LUT4AB_ConfigMem.ConfigBits\[451\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG2 net111 net11 net197 net215
+ Inst_LUT4AB_ConfigMem.ConfigBits\[438\] Inst_LUT4AB_ConfigMem.ConfigBits\[439\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_EF_BEG2 sky130_fd_sc_hd__mux4_2
X_231_ W6BEG_outbuf_7.X VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_162_ Inst_LUT4AB_switch_matrix.S2BEG6 VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ EE4BEG_outbuf_9.X VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr._15_ Inst_LC_LUT4c_frame_config_dffesr._01_ Inst_LC_LUT4c_frame_config_dffesr._02_
+ Inst_LC_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit25 net67 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[167\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit14 net55 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[503\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_GH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_GH._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG0 net20 net172 net224 Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[362\] Inst_LUT4AB_ConfigMem.ConfigBits\[363\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_46_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4BEG_outbuf_7._0_ NN4BEG_outbuf_7.A VGND VGND VPWR VPWR NN4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
Xinput1 Ci VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit5 net77 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[384\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput371 net371 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput360 net360 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput393 net393 VGND VGND VPWR VPWR NN4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput382 net382 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst1 net535 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 Inst_LUT4AB_switch_matrix.J2END_AB_BEG0
+ Inst_LUT4AB_ConfigMem.ConfigBits\[199\] Inst_LUT4AB_ConfigMem.ConfigBits\[200\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_145_ NN4BEG_outbuf_9.X VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit29 net71 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[202\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit18 net59 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[551\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_214_ Inst_LUT4AB_switch_matrix.W2BEG6 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_1
X_076_ strobe_outbuf_12.X VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._086_ Inst_LUT4AB_switch_matrix.JW2BEG0 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG0 sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[472\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[473\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG5
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit5 net77 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[312\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LB_LUT4c_frame_config_dffesr.I0mux
+ Inst_LB_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG1 net117 net17 net169 net221
+ Inst_LUT4AB_ConfigMem.ConfigBits\[404\] Inst_LUT4AB_ConfigMem.ConfigBits\[405\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_11_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_83 EE4BEG_outbuf_1.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_72 net539 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_50 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit13 net54 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[537\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit24 net66 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[565\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_94 W6BEG_outbuf_6.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst3 net509
+ net508 net511 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[510\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[511\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ N4BEG_outbuf_8.X VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._069_ net121 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb7
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_059_ Inst_LUT4AB_switch_matrix.E2BEG3 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkbuf_1
XNN4END_inbuf_4._0_ net152 VGND VGND VPWR VPWR NN4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XW6END_inbuf_0._0_ net230 VGND VGND VPWR VPWR W6BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[345\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._1_
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
Xinput70 FrameData[28] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_8
Xinput81 FrameData[9] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_8
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit8 net80 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[459\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput92 FrameStrobe[19] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_8
XInst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LC_LUT4c_frame_config_dffesr.I0mux
+ Inst_LC_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit28 net70 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[169\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit17 net58 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[514\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LE_LUT4c_frame_config_dffesr._18_ Inst_LE_LUT4c_frame_config_dffesr.SR Inst_LE_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XInst_LA_LUT4c_frame_config_dffesr._11_ Inst_LA_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit8 net80 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[400\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XWW4END_inbuf_10._0_ net243 VGND VGND VPWR VPWR WW4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S0 Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_switch_matrix.JE2BEG4 Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_switch_matrix.JW2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[346\] Inst_LUT4AB_ConfigMem.ConfigBits\[347\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S0 sky130_fd_sc_hd__mux4_2
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4BEG_outbuf_11._0_ N4BEG_outbuf_11.A VGND VGND VPWR VPWR N4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit12 net53 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[568\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit23 net65 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[243\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG0 net131 net9 net213 Inst_LUT4AB_switch_matrix.JN2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[594\] Inst_LUT4AB_ConfigMem.ConfigBits\[595\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4END_inbuf_9._0_ net178 VGND VGND VPWR VPWR S4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit19 net60 net83 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit27 net69 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[164\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit16 net57 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[495\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr._16_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[306\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._1_
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I0 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 Inst_LUT4AB_switch_matrix.J2END_AB_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[277\] Inst_LUT4AB_ConfigMem.ConfigBits\[278\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LB_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AD._4_ Inst_LUT4AB_switch_matrix.S1 Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._0_
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._1_ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.AD
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit3 net75 net90 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst1 net25 net197
+ net211 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[450\] Inst_LUT4AB_ConfigMem.ConfigBits\[451\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG3 net146 net7 net159 net211
+ Inst_LUT4AB_ConfigMem.ConfigBits\[440\] Inst_LUT4AB_ConfigMem.ConfigBits\[441\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_161_ Inst_LUT4AB_switch_matrix.S2BEG5 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_230_ W6BEG_outbuf_6.X VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkbuf_1
X_092_ EE4BEG_outbuf_8.X VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr._14_ Inst_LC_LUT4c_frame_config_dffesr.I\[1\] Inst_LC_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LC_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit26 net68 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[163\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit15 net56 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[499\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_20._0_ net62 VGND VGND VPWR VPWR data_inbuf_20.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG1 net116 net16 net220 Inst_LUT4AB_switch_matrix.JE2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[364\] Inst_LUT4AB_ConfigMem.ConfigBits\[365\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 E1END[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst0 net103
+ net109 net131 net9 Inst_LUT4AB_ConfigMem.ConfigBits\[490\] Inst_LUT4AB_ConfigMem.ConfigBits\[491\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_inbuf_11._0_ net52 VGND VGND VPWR VPWR data_inbuf_11.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput350 net350 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput361 net361 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit6 net78 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[383\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput394 net394 VGND VGND VPWR VPWR NN4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput383 net383 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput372 net372 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_075_ strobe_outbuf_11.X VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_1
X_144_ NN4BEG_outbuf_8.X VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit19 net60 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[548\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._085_ net173 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb7
+ sky130_fd_sc_hd__clkbuf_1
X_213_ Inst_LUT4AB_switch_matrix.W2BEG5 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG2 net119 net19 net171 net223
+ Inst_LUT4AB_ConfigMem.ConfigBits\[406\] Inst_LUT4AB_ConfigMem.ConfigBits\[407\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit6 net78 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[310\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_28_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LB_LUT4c_frame_config_dffesr.I0mux
+ Inst_LB_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LF_LUT4c_frame_config_dffesr._19_ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LF_LUT4c_frame_config_dffesr.SR Inst_LF_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr._12_ Inst_LB_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_95 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 net542 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit14 net55 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[534\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit25 net67 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[563\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_40 W6BEG_outbuf_8.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 Inst_LB_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_62 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_14._0_ strobe_inbuf_14.X VGND VGND VPWR VPWR strobe_outbuf_14.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[512\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[513\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG7
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix._068_ net120 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
X_127_ N4BEG_outbuf_7.X VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_9._0_ data_inbuf_9.X VGND VGND VPWR VPWR data_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
X_058_ Inst_LUT4AB_switch_matrix.E2BEG2 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkbuf_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[345\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput71 FrameData[29] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_8
Xinput60 FrameData[19] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_8
XInst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LC_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LC_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
Xinput93 FrameStrobe[1] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_16
Xinput82 FrameStrobe[0] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_8
XInst_LUT4AB_ConfigMem.Inst_Frame6_bit9 net81 net98 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[485\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame6_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit18 net59 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[509\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit29 net71 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[203\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XWW4END_inbuf_5._0_ net253 VGND VGND VPWR VPWR WW4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._2_ Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O._0_ sky130_fd_sc_hd__inv_2
XInst_LE_LUT4c_frame_config_dffesr._17_ Inst_LE_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst0 net103
+ net111 net3 net11 Inst_LUT4AB_ConfigMem.ConfigBits\[562\] Inst_LUT4AB_ConfigMem.ConfigBits\[563\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I0 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 Inst_LUT4AB_switch_matrix.J2END_EF_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[307\] Inst_LUT4AB_ConfigMem.ConfigBits\[308\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame11_bit9 net81 net84 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[417\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame11_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[231\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.SS4BEG1 sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1 Inst_LUT4AB_switch_matrix.JN2BEG5
+ Inst_LUT4AB_switch_matrix.JE2BEG5 Inst_LUT4AB_switch_matrix.JS2BEG5 Inst_LUT4AB_switch_matrix.JW2BEG5
+ Inst_LUT4AB_ConfigMem.ConfigBits\[348\] Inst_LUT4AB_ConfigMem.ConfigBits\[349\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1 sky130_fd_sc_hd__mux4_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit13 net54 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[159\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit24 net66 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[242\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG1 net146 net8 net182 Inst_LUT4AB_switch_matrix.JE2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[596\] Inst_LUT4AB_ConfigMem.ConfigBits\[597\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_62_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput250 WW4END[6] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit28 net70 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[162\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit17 net58 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[491\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr._15_ Inst_LD_LUT4c_frame_config_dffesr._01_ Inst_LD_LUT4c_frame_config_dffesr._02_
+ Inst_LD_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_11._0_ net84 VGND VGND VPWR VPWR strobe_inbuf_11.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst0 net110
+ net4 net10 net22 Inst_LUT4AB_ConfigMem.ConfigBits\[526\] Inst_LUT4AB_ConfigMem.ConfigBits\[527\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6END_inbuf_5._0_ net31 VGND VGND VPWR VPWR E6BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[306\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit1 net61 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[348\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I1 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 Inst_LUT4AB_switch_matrix.J2END_AB_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[279\] Inst_LUT4AB_ConfigMem.ConfigBits\[280\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_AD._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN\[1\]
+ Inst_LUT4AB_switch_matrix.S1 VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit4 net76 net90 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst2 net513
+ net537 net510 net509 Inst_LUT4AB_ConfigMem.ConfigBits\[450\] Inst_LUT4AB_ConfigMem.ConfigBits\[451\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AH.break_comb_loop_inst0._0_ Inst_MUX8LUT_frame_config_mux.AD
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG0 net508 Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3
+ Inst_LUT4AB_switch_matrix.JS2BEG3 Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[238\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[239\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_2
XSS4END_inbuf_7._0_ net192 VGND VGND VPWR VPWR SS4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_091_ EE4BEG_outbuf_7.X VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
X_160_ Inst_LUT4AB_switch_matrix.S2BEG4 VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit16 net57 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[498\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit27 net69 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[257\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG2 net118 net18 net170 Inst_LUT4AB_switch_matrix.JS2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[366\] Inst_LUT4AB_ConfigMem.ConfigBits\[367\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_23_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_9._0_ strobe_inbuf_9.X VGND VGND VPWR VPWR strobe_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
Xinput3 E1END[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst1 net25 net161
+ net213 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[490\] Inst_LUT4AB_ConfigMem.ConfigBits\[491\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit7 net79 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[382\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput373 net373 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput362 net362 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput340 net340 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput351 net351 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput395 net395 VGND VGND VPWR VPWR NN4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput384 net384 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__clkbuf_4
XEE4END_inbuf_6._0_ net35 VGND VGND VPWR VPWR EE4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_212_ Inst_LUT4AB_switch_matrix.W2BEG4 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
X_143_ NN4BEG_outbuf_7.X VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_1
X_074_ strobe_outbuf_10.X VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_3._0_ net75 VGND VGND VPWR VPWR data_inbuf_3.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._084_ net172 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
XWW4BEG_outbuf_7._0_ WW4BEG_outbuf_7.A VGND VGND VPWR VPWR WW4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I0 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 Inst_LUT4AB_switch_matrix.J2END_GH_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[337\] Inst_LUT4AB_ConfigMem.ConfigBits\[338\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit7 net79 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[308\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG3 net115 net15 net167 net219
+ Inst_LUT4AB_ConfigMem.ConfigBits\[408\] Inst_LUT4AB_ConfigMem.ConfigBits\[409\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 sky130_fd_sc_hd__mux4_2
XInst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LB_LUT4c_frame_config_dffesr.I0mux
+ Inst_LB_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LF_LUT4c_frame_config_dffesr._18_ Inst_LF_LUT4c_frame_config_dffesr.SR Inst_LF_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LB_LUT4c_frame_config_dffesr._11_ Inst_LB_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[615\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_EN_BEG0 sky130_fd_sc_hd__o21ai_4
XANTENNA_96 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit15 net56 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[530\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_85 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit26 net68 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[262\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_30 S4BEG_outbuf_3.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_74 net542 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 WW4BEG_outbuf_2.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinst_clk_buf UserCLK VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix._067_ net119 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb5
+ sky130_fd_sc_hd__clkbuf_1
X_126_ N4BEG_outbuf_6.X VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
X_057_ Inst_LUT4AB_switch_matrix.E2BEG1 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkbuf_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR._0_ sky130_fd_sc_hd__inv_2
Xinput50 FrameData[0] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_6
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput72 FrameData[2] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_8
Xinput61 FrameData[1] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_8
XFILLER_0_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XN4END_inbuf_9._0_ net126 VGND VGND VPWR VPWR N4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_2
Xinput83 FrameStrobe[10] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_16
Xinput94 FrameStrobe[2] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit19 net60 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[489\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LE_LUT4c_frame_config_dffesr._16_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst1 net155
+ net157 net163 net207 Inst_LUT4AB_ConfigMem.ConfigBits\[562\] Inst_LUT4AB_ConfigMem.ConfigBits\[563\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XN4BEG_outbuf_1._0_ N4BEG_outbuf_1.A VGND VGND VPWR VPWR N4BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I1 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 Inst_LUT4AB_switch_matrix.J2END_EF_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[309\] Inst_LUT4AB_ConfigMem.ConfigBits\[310\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[231\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
X_109_ Inst_LUT4AB_switch_matrix.N2BEG5 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S2 Inst_LUT4AB_switch_matrix.JN2BEG6
+ Inst_LUT4AB_switch_matrix.JE2BEG6 Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_switch_matrix.JW2BEG6
+ Inst_LUT4AB_ConfigMem.ConfigBits\[350\] Inst_LUT4AB_ConfigMem.ConfigBits\[351\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2 sky130_fd_sc_hd__mux4_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4BEG_outbuf_0._0_ SS4BEG_outbuf_0.A VGND VGND VPWR VPWR SS4BEG_outbuf_0.X sky130_fd_sc_hd__buf_2
XFILLER_0_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit14 net55 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[158\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst0 net105
+ net113 net5 net13 Inst_LUT4AB_ConfigMem.ConfigBits\[474\] Inst_LUT4AB_ConfigMem.ConfigBits\[475\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG2 net129 net197 net214 Inst_LUT4AB_switch_matrix.JS2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[598\] Inst_LUT4AB_ConfigMem.ConfigBits\[599\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput240 WW4END[11] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
Xinput251 WW4END[7] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkbuf_1
XW6BEG_outbuf_1._0_ W6BEG_outbuf_1.A VGND VGND VPWR VPWR W6BEG_outbuf_1.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit29 net71 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[153\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit18 net59 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[505\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr._14_ Inst_LD_LUT4c_frame_config_dffesr.I\[1\] Inst_LD_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LD_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst1 net162
+ net174 net214 net246 Inst_LUT4AB_ConfigMem.ConfigBits\[526\] Inst_LUT4AB_ConfigMem.ConfigBits\[527\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I2 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 Inst_LUT4AB_switch_matrix.J2END_AB_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[281\] Inst_LUT4AB_ConfigMem.ConfigBits\[282\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
Xdata_outbuf_30._0_ data_inbuf_30.X VGND VGND VPWR VPWR data_outbuf_30.X sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AD._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AD._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit5 net77 net90 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst3 Inst_LF_LUT4c_frame_config_dffesr.O
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AB Inst_LUT4AB_ConfigMem.ConfigBits\[450\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[451\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG1 net511 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0
+ Inst_LUT4AB_switch_matrix.JS2BEG0 Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[240\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[241\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_1
Xoutput500 net500 VGND VGND VPWR VPWR WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xdata_outbuf_21._0_ data_inbuf_21.X VGND VGND VPWR VPWR data_outbuf_21.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LG_LUT4c_frame_config_dffesr._19_ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LG_LUT4c_frame_config_dffesr.SR Inst_LG_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_090_ EE4BEG_outbuf_6.X VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LC_LUT4c_frame_config_dffesr._12_ Inst_LC_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LA_LUT4c_frame_config_dffesr.I0mux
+ Inst_LA_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xdata_outbuf_12._0_ data_inbuf_12.X VGND VGND VPWR VPWR data_outbuf_12.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit28 net70 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[251\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit17 net58 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[529\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_1._0_ S4BEG_outbuf_1.A VGND VGND VPWR VPWR S4BEG_outbuf_1.X sky130_fd_sc_hd__buf_2
XFILLER_0_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG3 net114 net166 net218
+ Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.ConfigBits\[368\] Inst_LUT4AB_ConfigMem.ConfigBits\[369\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 E1END[2] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.O
+ net532 Inst_LD_LUT4c_frame_config_dffesr.O net535 Inst_LUT4AB_ConfigMem.ConfigBits\[490\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[491\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit8 net80 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[379\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput341 net341 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput385 net385 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput374 net374 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput363 net363 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput352 net352 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput396 net396 VGND VGND VPWR VPWR NN4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput330 net330 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__buf_2
X_142_ NN4BEG_outbuf_6.X VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_211_ Inst_LUT4AB_switch_matrix.W2BEG3 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_073_ strobe_outbuf_9.X VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._083_ net171 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb5
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I1 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_switch_matrix.J2END_GH_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[339\] Inst_LUT4AB_ConfigMem.ConfigBits\[340\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XInst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LB_LUT4c_frame_config_dffesr.I0mux
+ Inst_LB_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit8 net80 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[307\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LF_LUT4c_frame_config_dffesr._17_ Inst_LF_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4END_inbuf_7._0_ net140 VGND VGND VPWR VPWR NN4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XEE4BEG_outbuf_0._0_ EE4BEG_outbuf_0.A VGND VGND VPWR VPWR EE4BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XW6END_inbuf_3._0_ net233 VGND VGND VPWR VPWR W6BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[615\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_20 N4BEG_outbuf_9.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_31 S4BEG_outbuf_3.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_75 net542 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit27 net69 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[260\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_97 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit16 net57 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[560\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_42 WW4BEG_outbuf_7.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst0._0_ net518 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
X_125_ N4BEG_outbuf_5.X VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix._066_ net118 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_056_ Inst_LUT4AB_switch_matrix.E2BEG0 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_1
XFILLER_0_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput73 FrameData[30] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_8
XFILLER_0_71_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput62 FrameData[20] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_8
Xinput51 FrameData[10] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_8
Xmax_cap510 Inst_LD_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_12
Xinput40 EE4END[15] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput84 FrameStrobe[11] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_16
Xinput95 FrameStrobe[3] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst2 net514
+ Inst_LB_LUT4c_frame_config_dffesr.O Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[562\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[563\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LE_LUT4c_frame_config_dffesr._15_ Inst_LE_LUT4c_frame_config_dffesr._01_ Inst_LE_LUT4c_frame_config_dffesr._02_
+ Inst_LE_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
X_108_ Inst_LUT4AB_switch_matrix.N2BEG4 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix._049_ Inst_LC_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LD_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S3 Inst_LUT4AB_switch_matrix.JN2BEG7
+ Inst_LUT4AB_switch_matrix.JE2BEG7 Inst_LUT4AB_switch_matrix.JS2BEG7 Inst_LUT4AB_switch_matrix.JW2BEG7
+ Inst_LUT4AB_ConfigMem.ConfigBits\[352\] Inst_LUT4AB_ConfigMem.ConfigBits\[353\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S3 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I2 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 Inst_LUT4AB_switch_matrix.J2END_EF_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[311\] Inst_LUT4AB_ConfigMem.ConfigBits\[312\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
X_039_ Inst_LUT4AB_switch_matrix.E2BEGb7 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit0 net50 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[359\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit15 net56 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[157\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst1 net157
+ net165 net207 net209 Inst_LUT4AB_ConfigMem.ConfigBits\[474\] Inst_LUT4AB_ConfigMem.ConfigBits\[475\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit0 net50 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[330\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4BEG_outbuf_10._0_ EE4BEG_outbuf_10.A VGND VGND VPWR VPWR EE4BEG_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG3 net43 net174 net245 Inst_LUT4AB_switch_matrix.JW2BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[600\] Inst_LUT4AB_ConfigMem.ConfigBits\[601\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_65_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput241 WW4END[12] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
Xinput252 WW4END[8] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkbuf_1
Xinput230 W6END[2] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame3_bit19 net60 net95 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[501\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame3_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.O
+ Inst_LB_LUT4c_frame_config_dffesr.O net512 Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[526\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[527\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LB_I3 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 Inst_LUT4AB_switch_matrix.J2END_AB_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[283\] Inst_LUT4AB_ConfigMem.ConfigBits\[284\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_1
Xdata_inbuf_23._0_ net65 VGND VGND VPWR VPWR data_inbuf_23.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit6 net78 net90 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst0 net104 net4
+ net208 net541 Inst_LUT4AB_ConfigMem.ConfigBits\[170\] Inst_LUT4AB_ConfigMem.ConfigBits\[171\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[452\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[453\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG0
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG2 net515 Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1
+ Inst_LUT4AB_switch_matrix.JS2BEG1 Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[242\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[243\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_1
Xoutput501 net501 VGND VGND VPWR VPWR WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_2._0_ net94 VGND VGND VPWR VPWR strobe_inbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_14._0_ net55 VGND VGND VPWR VPWR data_inbuf_14.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LG_LUT4c_frame_config_dffesr._18_ Inst_LG_LUT4c_frame_config_dffesr.SR Inst_LG_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XInst_LC_LUT4c_frame_config_dffesr._11_ Inst_LC_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LA_LUT4c_frame_config_dffesr.I0mux
+ Inst_LA_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_110 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit18 net59 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[528\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XWW4BEG_outbuf_11._0_ WW4BEG_outbuf_11.A VGND VGND VPWR VPWR WW4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_2
Xinput5 E1END[3] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst3 net508
+ net511 Inst_LH_LUT4c_frame_config_dffesr.O Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[490\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[491\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit9 net81 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[378\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
Xoutput353 net353 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput397 net397 VGND VGND VPWR VPWR NN4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput375 net375 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput386 net386 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput364 net364 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput320 net320 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__clkbuf_4
X_141_ NN4BEG_outbuf_5.X VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix._082_ net170 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
X_210_ Inst_LUT4AB_switch_matrix.W2BEG2 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_1
X_072_ strobe_outbuf_8.X VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst0._0_ net527 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_17._0_ strobe_inbuf_17.X VGND VGND VPWR VPWR strobe_outbuf_17.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I2 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 Inst_LUT4AB_switch_matrix.J2END_GH_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[341\] Inst_LUT4AB_ConfigMem.ConfigBits\[342\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
XInst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LB_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LB_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit9 net81 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[334\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LF_LUT4c_frame_config_dffesr._16_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XANTENNA_21 NN4BEG_outbuf_1.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_65 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 WW4BEG_outbuf_8.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 S4BEG_outbuf_6.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_98 net102 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit17 net58 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[559\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_76 net543 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit28 net70 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[256\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[295\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._1_
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XWW4END_inbuf_8._0_ net241 VGND VGND VPWR VPWR WW4BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_1
X_124_ N4BEG_outbuf_4.X VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst0 net5 net209
+ net514 net532 Inst_LUT4AB_ConfigMem.ConfigBits\[258\] Inst_LUT4AB_ConfigMem.ConfigBits\[259\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
X_055_ Inst_LUT4AB_switch_matrix.E1BEG3 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._065_ net117 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb3
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput74 FrameData[31] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_8
Xinput52 FrameData[11] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_8
Xinput63 FrameData[21] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_8
Xmax_cap511 Inst_LG_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkbuf_8
Xinput30 E6END[6] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput41 EE4END[1] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput96 FrameStrobe[4] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_12
XFILLER_0_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput85 FrameStrobe[12] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LE_LUT4c_frame_config_dffesr._14_ Inst_LE_LUT4c_frame_config_dffesr.I\[1\] Inst_LE_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LE_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst3 net508
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[562\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[563\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ Inst_LUT4AB_switch_matrix.N2BEG3 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit1 net61 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[346\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
X_038_ Inst_LUT4AB_switch_matrix.E2BEGb6 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LE_I3 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 Inst_LUT4AB_switch_matrix.J2END_EF_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[313\] Inst_LUT4AB_ConfigMem.ConfigBits\[314\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_21_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._048_ Inst_LB_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LC_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__buf_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit16 net57 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[241\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst2 net514
+ net513 net537 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[474\] Inst_LUT4AB_ConfigMem.ConfigBits\[475\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit1 net61 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[338\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_14._0_ net87 VGND VGND VPWR VPWR strobe_inbuf_14.X sky130_fd_sc_hd__clkbuf_1
Xinput242 WW4END[13] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
Xinput253 WW4END[9] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkbuf_1
Xinput231 W6END[3] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
Xinput220 W2MID[2] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_4
XE6END_inbuf_8._0_ net23 VGND VGND VPWR VPWR E6BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_2
XInst_LH_LUT4c_frame_config_dffesr._19_ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LH_LUT4c_frame_config_dffesr.SR Inst_LH_LUT4c_frame_config_dffesr.EN VGND VGND
+ VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._09_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LD_LUT4c_frame_config_dffesr._12_ Inst_LD_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6BEG_outbuf_0._0_ E6BEG_outbuf_0.A VGND VGND VPWR VPWR E6BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[526\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[527\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit4 net76 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[366\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst1 net540 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2END_GH_BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[170\] Inst_LUT4AB_ConfigMem.ConfigBits\[171\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit7 net79 net90 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput502 net502 VGND VGND VPWR VPWR WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_W1BEG3 net543 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2
+ Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[244\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[245\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_49_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst0 net102 net154
+ net206 net532 Inst_LUT4AB_ConfigMem.ConfigBits\[252\] Inst_LUT4AB_ConfigMem.ConfigBits\[253\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_LG_LUT4c_frame_config_dffesr._17_ Inst_LG_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LA_LUT4c_frame_config_dffesr.I0mux
+ Inst_LA_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit19 net60 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[544\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_100 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XEE4END_inbuf_9._0_ net38 VGND VGND VPWR VPWR EE4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_6._0_ net78 VGND VGND VPWR VPWR data_inbuf_6.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 E2END[0] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[492\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[493\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_6_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput343 net343 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__buf_2
Xoutput321 net321 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput310 net310 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput332 net332 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
XInst_MUX8LUT_frame_config_mux.cus_mux21_sGH._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[152\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.S sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput387 net387 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput376 net376 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput365 net365 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput398 net398 VGND VGND VPWR VPWR NN4BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_071_ strobe_outbuf_7.X VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_1
X_140_ NN4BEG_outbuf_4.X VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix._081_ net169 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb3
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst0._0_ net523 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LH_I3 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 Inst_LUT4AB_switch_matrix.J2END_GH_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[343\] Inst_LUT4AB_ConfigMem.ConfigBits\[344\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_2
XFILLER_0_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LF_LUT4c_frame_config_dffesr._15_ Inst_LF_LUT4c_frame_config_dffesr._01_ Inst_LF_LUT4c_frame_config_dffesr._02_
+ Inst_LF_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_63_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_22 NN4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 Inst_LUT4AB_switch_matrix.N1BEG0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit18 net59 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[578\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_55 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 SS4BEG_outbuf_0.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 net543 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_88 Inst_LUT4AB_switch_matrix.W2BEGb7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 WW4BEG_outbuf_8.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[295\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit29 net71 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[255\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst0 net104 net4
+ net208 net541 Inst_LUT4AB_ConfigMem.ConfigBits\[226\] Inst_LUT4AB_ConfigMem.ConfigBits\[227\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_123_ N4BEG_outbuf_3.X VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._064_ net116 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst1 net537 net510
+ net509 net508 Inst_LUT4AB_ConfigMem.ConfigBits\[258\] Inst_LUT4AB_ConfigMem.ConfigBits\[259\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
X_054_ Inst_LUT4AB_switch_matrix.E1BEG2 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4BEG_outbuf_0._0_ NN4BEG_outbuf_0.A VGND VGND VPWR VPWR NN4BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XN4BEG_outbuf_4._0_ N4BEG_outbuf_4.A VGND VGND VPWR VPWR N4BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput31 E6END[7] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 E2MID[6] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 FrameData[22] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_8
Xinput53 FrameData[12] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_8
Xmax_cap512 Inst_LC_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_8
Xinput75 FrameData[3] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_8
Xinput42 EE4END[2] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput86 FrameStrobe[13] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_8
Xinput97 FrameStrobe[5] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4BEG_outbuf_3._0_ SS4BEG_outbuf_3.A VGND VGND VPWR VPWR SS4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst0._0__523 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_SR.break_comb_loop_inst0._0__523/HI
+ net523 sky130_fd_sc_hd__conb_1
XFILLER_0_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[564\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[565\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG4
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_30_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XSS4BEG_outbuf_11._0_ SS4BEG_outbuf_11.A VGND VGND VPWR VPWR SS4BEG_outbuf_11.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_106_ Inst_LUT4AB_switch_matrix.N2BEG2 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_1
X_037_ Inst_LUT4AB_switch_matrix.E2BEGb5 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit2 net72 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[421\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._047_ Inst_LA_LUT4c_frame_config_dffesr.Co VGND VGND VPWR
+ VPWR Inst_LB_LUT4c_frame_config_dffesr.Ci sky130_fd_sc_hd__clkbuf_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XW6BEG_outbuf_4._0_ W6BEG_outbuf_4.A VGND VGND VPWR VPWR W6BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit17 net58 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[240\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst3 net509
+ Inst_LF_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[474\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[475\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit2 net72 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[391\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput232 W6END[4] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
Xinput243 WW4END[14] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
Xinput221 W2MID[3] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__buf_2
Xinput210 W2END[0] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_58_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LH_LUT4c_frame_config_dffesr._18_ Inst_LH_LUT4c_frame_config_dffesr.SR Inst_LH_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._08_ sky130_fd_sc_hd__or2b_1
XFILLER_0_53_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr._11_ Inst_LD_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_24._0_ data_inbuf_24.X VGND VGND VPWR VPWR data_outbuf_24.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[528\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[529\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_35_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_15._0_ data_inbuf_15.X VGND VGND VPWR VPWR data_outbuf_15.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit5 net77 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[374\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_4._0_ S4BEG_outbuf_4.A VGND VGND VPWR VPWR S4BEG_outbuf_4.X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit8 net80 net90 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput503 net503 VGND VGND VPWR VPWR WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst1 net512 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_switch_matrix.J2END_CD_BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[252\] Inst_LUT4AB_ConfigMem.ConfigBits\[253\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LG_LUT4c_frame_config_dffesr._16_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LA_LUT4c_frame_config_dffesr.I0mux
+ Inst_LA_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XS4END_inbuf_2._0_ net186 VGND VGND VPWR VPWR S4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_1
XANTENNA_112 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 net170 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 E2END[1] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput366 net366 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput344 net344 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput377 net377 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput322 net322 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput311 net311 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput333 net333 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__clkbuf_4
XInst_MUX8LUT_frame_config_mux.cus_mux21_sGH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[152\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._1_
+ sky130_fd_sc_hd__nand2_1
Xoutput300 net300 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_0_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XW6END_inbuf_6._0_ net236 VGND VGND VPWR VPWR W6BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_1
Xoutput399 net399 VGND VGND VPWR VPWR NN4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput388 net388 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__clkbuf_4
XEE4BEG_outbuf_3._0_ EE4BEG_outbuf_3.A VGND VGND VPWR VPWR EE4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
X_070_ strobe_outbuf_6.X VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix._080_ net168 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LF_LUT4c_frame_config_dffesr._14_ Inst_LF_LUT4c_frame_config_dffesr.I\[1\] Inst_LF_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LF_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit0 net50 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[351\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_199_ SS4BEG_outbuf_11.X VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_23 NN4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 Inst_LUT4AB_switch_matrix.N1BEG3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 NN4BEG_outbuf_0.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit19 net60 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[573\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_67 net209 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 SS4BEG_outbuf_0.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 net543 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst1 net540 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2END_GH_BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[226\] Inst_LUT4AB_ConfigMem.ConfigBits\[227\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst2 net540 net515
+ net542 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[258\] Inst_LUT4AB_ConfigMem.ConfigBits\[259\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit0 net50 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[302\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
X_122_ N4BEG_outbuf_2.X VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
X_053_ Inst_LUT4AB_switch_matrix.E1BEG1 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__buf_1
XFILLER_0_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix._063_ net115 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb1
+ sky130_fd_sc_hd__clkbuf_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EF._4_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_EF sky130_fd_sc_hd__o21ai_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst0 net108
+ net130 net2 net8 Inst_LUT4AB_ConfigMem.ConfigBits\[454\] Inst_LUT4AB_ConfigMem.ConfigBits\[455\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput54 FrameData[13] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_8
XFILLER_0_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 E6END[8] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 EE4END[3] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput21 E2MID[7] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xinput10 E2END[4] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
Xinput65 FrameData[23] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_8
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput76 FrameData[4] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_8
Xinput87 FrameStrobe[14] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_8
Xinput98 FrameStrobe[6] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
Xmax_cap513 Inst_LB_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LE_LUT4c_frame_config_dffesr._12_ Inst_LE_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEH.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.S3
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LE_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
X_105_ Inst_LUT4AB_switch_matrix.N2BEG1 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit3 net75 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[429\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
X_036_ Inst_LUT4AB_switch_matrix.E2BEGb4 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix._046_ net1 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.Ci
+ sky130_fd_sc_hd__buf_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit18 net59 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[263\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XN4END_inbuf_10._0_ net127 VGND VGND VPWR VPWR N4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[476\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[477\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG6
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[228\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.SS4BEG0 sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst0._0__518 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_SR.break_comb_loop_inst0._0__518/HI
+ net518 sky130_fd_sc_hd__conb_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit3 net75 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[390\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput200 SS4END[4] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_2._0_ data_inbuf_2.X VGND VGND VPWR VPWR data_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xinput233 W6END[5] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
Xinput244 WW4END[15] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
Xinput222 W2MID[4] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_4
Xinput211 W2END[1] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_4
XInst_LH_LUT4c_frame_config_dffesr._17_ Inst_LH_LUT4c_frame_config_dffesr.EN VGND
+ VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._07_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_019_ data_outbuf_19.X VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_26._0_ net68 VGND VGND VPWR VPWR data_inbuf_26.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_inbuf_5._0_ net97 VGND VGND VPWR VPWR strobe_inbuf_5.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_inbuf_17._0_ net58 VGND VGND VPWR VPWR data_inbuf_17.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit6 net78 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[423\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit9 net81 net90 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput504 net504 VGND VGND VPWR VPWR WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LG_LUT4c_frame_config_dffesr._15_ Inst_LG_LUT4c_frame_config_dffesr._01_ Inst_LG_LUT4c_frame_config_dffesr._02_
+ Inst_LG_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst4 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3 Inst_LA_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LA_LUT4c_frame_config_dffesr.I\[3\] VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.LUT_out
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_113 EE4BEG_outbuf_2.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 E2END[2] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XS4END_inbuf_10._0_ net179 VGND VGND VPWR VPWR S4BEG_outbuf_10.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst0._0__527 VGND
+ VGND VPWR VPWR net527 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_EN.break_comb_loop_inst0._0__527/LO
+ sky130_fd_sc_hd__conb_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sGH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput345 net345 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput378 net378 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput389 net389 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput367 net367 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput356 net356 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput323 net323 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput312 net312 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput334 net334 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__buf_2
Xoutput301 net301 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit1 net61 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[329\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_198_ SS4BEG_outbuf_10.X VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 Inst_LUT4AB_switch_matrix.N2BEG1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[316\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._1_
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_24 NN4BEG_outbuf_2.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_57 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_35 SS4BEG_outbuf_1.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 net543 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XSS4END_inbuf_0._0_ net200 VGND VGND VPWR VPWR SS4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_1
X_121_ N4BEG_outbuf_1.X VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._062_ net114 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.N2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit1 net61 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[326\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[258\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[259\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
X_052_ Inst_LUT4AB_switch_matrix.E1BEG0 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EF._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN\[1\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst1 net22 net160
+ net212 net226 Inst_LUT4AB_ConfigMem.ConfigBits\[454\] Inst_LUT4AB_ConfigMem.ConfigBits\[455\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_2._0_ strobe_inbuf_2.X VGND VGND VPWR VPWR strobe_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xinput66 FrameData[24] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_8
Xinput55 FrameData[14] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_8
Xinput77 FrameData[5] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_16
Xinput33 E6END[9] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput22 E6END[0] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_4
Xinput44 EE4END[4] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput11 E2END[5] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap514 Inst_LA_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_12
XFILLER_0_3_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput88 FrameStrobe[15] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_8
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput99 FrameStrobe[7] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_12
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LE_LUT4c_frame_config_dffesr._11_ Inst_LE_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_104_ Inst_LUT4AB_switch_matrix.N2BEG0 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._045_ net515 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.H
+ sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_17._0_ net90 VGND VGND VPWR VPWR strobe_inbuf_17.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_035_ Inst_LUT4AB_switch_matrix.E2BEGb3 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XWW4BEG_outbuf_0._0_ WW4BEG_outbuf_0.A VGND VGND VPWR VPWR WW4BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst0 net104
+ net110 net122 net10 Inst_LUT4AB_ConfigMem.ConfigBits\[494\] Inst_LUT4AB_ConfigMem.ConfigBits\[495\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit4 net76 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[454\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit19 net60 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[261\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[228\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit4 net76 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[381\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput201 SS4END[5] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XE6BEG_outbuf_3._0_ E6BEG_outbuf_3.A VGND VGND VPWR VPWR E6BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
Xinput234 W6END[6] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
Xinput212 W2END[2] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__buf_2
Xinput223 W2MID[5] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_2
Xinput245 WW4END[1] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_2
XInst_LH_LUT4c_frame_config_dffesr._16_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._06_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_018_ data_outbuf_18.X VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XN4END_inbuf_2._0_ net134 VGND VGND VPWR VPWR N4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_2
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit7 net79 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[439\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_inbuf_9._0_ net81 VGND VGND VPWR VPWR data_inbuf_9.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput505 net505 VGND VGND VPWR VPWR WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst0 net104
+ net112 net4 net12 Inst_LUT4AB_ConfigMem.ConfigBits\[566\] Inst_LUT4AB_ConfigMem.ConfigBits\[567\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LG_LUT4c_frame_config_dffesr._14_ Inst_LG_LUT4c_frame_config_dffesr.I\[1\] Inst_LG_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LG_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 EE4BEG_outbuf_4.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 net208 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 E2END[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput346 net346 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput379 net379 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput368 net368 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput357 net357 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput324 net324 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput302 net302 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LF_LUT4c_frame_config_dffesr._12_ Inst_LF_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit2 net72 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[369\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_197_ SS4BEG_outbuf_9.X VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XNN4BEG_outbuf_3._0_ NN4BEG_outbuf_3.A VGND VGND VPWR VPWR NN4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XN4BEG_outbuf_7._0_ N4BEG_outbuf_7.A VGND VGND VPWR VPWR N4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_14 Inst_LUT4AB_switch_matrix.N2BEG2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 NN4BEG_outbuf_3.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst0 net103
+ net111 net3 net11 Inst_LUT4AB_ConfigMem.ConfigBits\[530\] Inst_LUT4AB_ConfigMem.ConfigBits\[531\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[316\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_36 SS4BEG_outbuf_2.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_69 net222 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XSS4BEG_outbuf_6._0_ SS4BEG_outbuf_6.A VGND VGND VPWR VPWR SS4BEG_outbuf_6.X sky130_fd_sc_hd__buf_2
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XS4BEG_outbuf_10._0_ S4BEG_outbuf_10.A VGND VGND VPWR VPWR S4BEG_outbuf_10.X sky130_fd_sc_hd__buf_2
X_120_ N4BEG_outbuf_0.X VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._061_ Inst_LUT4AB_switch_matrix.JN2BEG7 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_051_ Inst_LUT4AB_switch_matrix.E6BEG1 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit2 net72 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[321\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[260\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[261\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W6BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EF._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EF._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst2 net514
+ net512 net510 net509 Inst_LUT4AB_ConfigMem.ConfigBits\[454\] Inst_LUT4AB_ConfigMem.ConfigBits\[455\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput67 FrameData[25] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_8
Xmax_cap515 Inst_LH_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_8
Xinput56 FrameData[15] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_8
Xinput78 FrameData[6] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_8
Xinput23 E6END[10] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput45 EE4END[5] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 EE4END[0] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput12 E2END[6] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput89 FrameStrobe[16] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_8
X_249_ Inst_LUT4AB_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_AD.break_comb_loop_inst0._0_ net542 VGND
+ VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AD.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XW6BEG_outbuf_7._0_ W6BEG_outbuf_7.A VGND VGND VPWR VPWR W6BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_103_ Inst_LUT4AB_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit5 net77 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[453\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._044_ net540 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.G
+ sky130_fd_sc_hd__clkbuf_1
X_034_ Inst_LUT4AB_switch_matrix.E2BEGb2 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst1 net22 net162
+ net214 net226 Inst_LUT4AB_ConfigMem.ConfigBits\[494\] Inst_LUT4AB_ConfigMem.ConfigBits\[495\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LH_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XNN4END_inbuf_0._0_ net148 VGND VGND VPWR VPWR NN4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit5 net77 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[380\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput202 SS4END[6] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_27._0_ data_inbuf_27.X VGND VGND VPWR VPWR data_outbuf_27.X sky130_fd_sc_hd__clkbuf_1
Xinput235 W6END[7] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_1
Xinput224 W2MID[6] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_4
Xinput213 W2END[3] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput246 WW4END[2] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__buf_2
XInst_LH_LUT4c_frame_config_dffesr._15_ Inst_LH_LUT4c_frame_config_dffesr._01_ Inst_LH_LUT4c_frame_config_dffesr._02_
+ Inst_LH_LUT4c_frame_config_dffesr._05_ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.Co
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_18._0_ data_inbuf_18.X VGND VGND VPWR VPWR data_outbuf_18.X sky130_fd_sc_hd__clkbuf_1
X_017_ data_outbuf_17.X VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XS4BEG_outbuf_7._0_ S4BEG_outbuf_7.A VGND VGND VPWR VPWR S4BEG_outbuf_7.X sky130_fd_sc_hd__clkbuf_2
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XS4END_inbuf_5._0_ net189 VGND VGND VPWR VPWR S4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit8 net80 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[464\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput506 net506 VGND VGND VPWR VPWR WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_72_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst1 net154
+ net156 net164 net208 Inst_LUT4AB_ConfigMem.ConfigBits\[566\] Inst_LUT4AB_ConfigMem.ConfigBits\[567\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XEE4BEG_outbuf_6._0_ EE4BEG_outbuf_6.A VGND VGND VPWR VPWR EE4BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XW6END_inbuf_9._0_ net228 VGND VGND VPWR VPWR W6BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit0 net50 net89 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[335\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_104 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 EE4BEG_outbuf_4.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst0 net102
+ net106 net2 net34 Inst_LUT4AB_ConfigMem.ConfigBits\[478\] Inst_LUT4AB_ConfigMem.ConfigBits\[479\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xoutput325 net325 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput314 net314 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput303 net303 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput369 net369 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput347 net347 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput336 net336 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG0 net113 net13 net165 net238
+ Inst_LUT4AB_ConfigMem.ConfigBits\[442\] Inst_LUT4AB_ConfigMem.ConfigBits\[443\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_GH_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_68_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LF_LUT4c_frame_config_dffesr._11_ Inst_LF_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_196_ SS4BEG_outbuf_8.X VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit3 net75 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[432\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_15 Inst_LUT4AB_switch_matrix.N4BEG3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 NN4BEG_outbuf_5.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_59 net158 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst1 net155
+ net163 net207 net209 Inst_LUT4AB_ConfigMem.ConfigBits\[530\] Inst_LUT4AB_ConfigMem.ConfigBits\[531\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_48 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_37 SS4BEG_outbuf_7.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._060_ Inst_LUT4AB_switch_matrix.JN2BEG6 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG6 sky130_fd_sc_hd__clkbuf_1
X_050_ Inst_LUT4AB_switch_matrix.E6BEG0 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit3 net75 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[313\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XNN4BEG_outbuf_10._0_ NN4BEG_outbuf_10.A VGND VGND VPWR VPWR NN4BEG_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[454\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[455\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput13 E2END[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_0_33_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput68 FrameData[26] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_8
Xinput57 FrameData[16] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_8
Xinput79 FrameData[7] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_8
XFILLER_0_58_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput24 E6END[11] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput35 EE4END[10] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput46 EE4END[6] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_179_ S4BEG_outbuf_7.X VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_1
X_248_ Inst_LUT4AB_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG0 net121 net21 net173 net225
+ Inst_LUT4AB_ConfigMem.ConfigBits\[410\] Inst_LUT4AB_ConfigMem.ConfigBits\[411\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG0 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix._112_ Inst_LUT4AB_switch_matrix.JE2BEG4 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG4 sky130_fd_sc_hd__buf_1
Xstrobe_outbuf_10._0_ strobe_inbuf_10.X VGND VGND VPWR VPWR strobe_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
X_102_ Inst_LUT4AB_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._043_ Inst_LF_LUT4c_frame_config_dffesr.O VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.F sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_033_ Inst_LUT4AB_switch_matrix.E2BEGb1 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit6 net78 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[448\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst2 Inst_LA_LUT4c_frame_config_dffesr.O
+ net513 net512 net535 Inst_LUT4AB_ConfigMem.ConfigBits\[494\] Inst_LUT4AB_ConfigMem.ConfigBits\[495\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
Xdata_outbuf_5._0_ data_inbuf_5.X VGND VGND VPWR VPWR data_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_29._0_ net71 VGND VGND VPWR VPWR data_inbuf_29.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XWW4END_inbuf_1._0_ net249 VGND VGND VPWR VPWR WW4BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit6 net78 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[377\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput203 SS4END[7] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_8._0_ net100 VGND VGND VPWR VPWR strobe_inbuf_8.X sky130_fd_sc_hd__clkbuf_1
Xinput236 W6END[8] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
Xinput225 W2MID[7] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__buf_2
Xinput214 W2END[4] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_4
Xinput247 WW4END[3] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LH_LUT4c_frame_config_dffesr._14_ Inst_LH_LUT4c_frame_config_dffesr.I\[1\] Inst_LH_LUT4c_frame_config_dffesr.I\[2\]
+ Inst_LH_LUT4c_frame_config_dffesr.Ci VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._05_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_016_ data_outbuf_16.X VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame2_bit9 net81 net94 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[461\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame2_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput507 net507 VGND VGND VPWR VPWR WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst2 net514
+ net532 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[566\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[567\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LG_LUT4c_frame_config_dffesr._12_ Inst_LG_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit1 net61 net89 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[345\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_105 net216 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 W6BEG_outbuf_0.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XE6END_inbuf_1._0_ net27 VGND VGND VPWR VPWR E6BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux41_buf_inst0 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[613\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[614\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LG_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput348 net348 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__clkbuf_4
Xoutput359 net359 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput337 net337 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput326 net326 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__clkbuf_4
Xoutput315 net315 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput304 net304 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst1 net154
+ net158 net206 net208 Inst_LUT4AB_ConfigMem.ConfigBits\[478\] Inst_LUT4AB_ConfigMem.ConfigBits\[479\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XSS4END_inbuf_3._0_ net203 VGND VGND VPWR VPWR SS4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG1 net109 net9 net190 net213
+ Inst_LUT4AB_ConfigMem.ConfigBits\[444\] Inst_LUT4AB_ConfigMem.ConfigBits\[445\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_GH_BEG1 sky130_fd_sc_hd__mux4_2
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit4 net76 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[427\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
X_195_ SS4BEG_outbuf_7.X VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_5._0_ strobe_inbuf_5.X VGND VGND VPWR VPWR strobe_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LE_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_49 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 N4BEG_outbuf_0.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_27 NN4BEG_outbuf_6.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst2 net514
+ net513 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[530\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[531\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XANTENNA_38 W6BEG_outbuf_1.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit4 net76 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[306\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG0 net120 net20 net224 Inst_LUT4AB_switch_matrix.JN2BEG5
+ Inst_LUT4AB_ConfigMem.ConfigBits\[370\] Inst_LUT4AB_ConfigMem.ConfigBits\[371\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0 sky130_fd_sc_hd__mux4_2
XEE4END_inbuf_2._0_ net46 VGND VGND VPWR VPWR EE4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst0 net105 net5
+ net209 net514 Inst_LUT4AB_ConfigMem.ConfigBits\[173\] Inst_LUT4AB_ConfigMem.ConfigBits\[174\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG0 net535 Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3
+ Inst_LUT4AB_switch_matrix.JE2BEG3 Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[210\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[211\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[456\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[457\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput25 E6END[1] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_4
Xinput36 EE4END[11] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 E2MID[0] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
X_247_ WW4BEG_outbuf_11.X VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkbuf_1
XWW4BEG_outbuf_3._0_ WW4BEG_outbuf_3.A VGND VGND VPWR VPWR WW4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_2
Xinput69 FrameData[27] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_8
Xinput58 FrameData[17] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_8
Xinput47 EE4END[7] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
X_178_ S4BEG_outbuf_6.X VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_101_ Inst_LUT4AB_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix._042_ net21 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb7
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._111_ Inst_LUT4AB_switch_matrix.JE2BEG3 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG3 sky130_fd_sc_hd__buf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG1 net117 net17 net169 net221
+ Inst_LUT4AB_ConfigMem.ConfigBits\[412\] Inst_LUT4AB_ConfigMem.ConfigBits\[413\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit7 net79 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[444\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
X_032_ Inst_LUT4AB_switch_matrix.E2BEGb0 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[494\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[495\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XE6BEG_outbuf_6._0_ E6BEG_outbuf_6.A VGND VGND VPWR VPWR E6BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XN4END_inbuf_5._0_ net137 VGND VGND VPWR VPWR N4BEG_outbuf_5.A sky130_fd_sc_hd__buf_2
XFILLER_0_18_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_115 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit7 net79 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[376\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput204 SS4END[8] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
Xinput237 W6END[9] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkbuf_1
Xinput226 W6END[0] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput215 W2END[5] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_2
Xinput248 WW4END[4] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_1
X_015_ data_outbuf_15.X VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[305\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._1_
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst0 net4 net208
+ net514 net532 Inst_LUT4AB_ConfigMem.ConfigBits\[262\] Inst_LUT4AB_ConfigMem.ConfigBits\[263\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH.break_comb_loop_inst0._0_ Inst_LUT4AB_switch_matrix.M_EF
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst0._0_ net519 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_39_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst3 net509
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[566\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[567\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LG_LUT4c_frame_config_dffesr._11_ Inst_LG_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 EE4BEG_outbuf_0.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 WW4BEG_outbuf_9.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit2 net72 net89 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix.JN2BEG2
+ Inst_LUT4AB_switch_matrix.JE2BEG2 Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_switch_matrix.JW2BEG2
+ Inst_LUT4AB_ConfigMem.ConfigBits\[613\] Inst_LUT4AB_ConfigMem.ConfigBits\[614\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_EN_BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput349 net349 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput338 net338 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput327 net327 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput305 net305 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst2 net514
+ net532 net537 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[478\] Inst_LUT4AB_ConfigMem.ConfigBits\[479\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4BEG_outbuf_6._0_ NN4BEG_outbuf_6.A VGND VGND VPWR VPWR NN4BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[266\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._1_
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4BEG_outbuf_9._0_ SS4BEG_outbuf_9.A VGND VGND VPWR VPWR SS4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[152\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.EH_GH sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG2 net145 net11 net163 net215
+ Inst_LUT4AB_ConfigMem.ConfigBits\[446\] Inst_LUT4AB_ConfigMem.ConfigBits\[447\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_GH_BEG2 sky130_fd_sc_hd__mux4_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit5 net77 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[426\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
X_194_ SS4BEG_outbuf_6.X VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_17 N4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst3 net508
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[530\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[531\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_39 W6BEG_outbuf_5.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 S4BEG_outbuf_0.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit5 net77 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[343\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst1 net515 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 Inst_LUT4AB_switch_matrix.J2END_EF_BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[173\] Inst_LUT4AB_ConfigMem.ConfigBits\[174\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG1 net116 net16 net168 Inst_LUT4AB_switch_matrix.JE2BEG5
+ Inst_LUT4AB_ConfigMem.ConfigBits\[372\] Inst_LUT4AB_ConfigMem.ConfigBits\[373\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG1 net508 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0
+ Inst_LUT4AB_switch_matrix.JE2BEG0 Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[212\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[213\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_1
Xinput59 FrameData[18] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_8
XFILLER_0_64_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput26 E6END[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 EE4END[12] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput48 EE4END[8] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xinput15 E2MID[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_246_ WW4BEG_outbuf_10.X VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkbuf_1
X_177_ S4BEG_outbuf_5.X VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst0 net103 net155
+ net207 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[255\] Inst_LUT4AB_ConfigMem.ConfigBits\[256\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XNN4END_inbuf_3._0_ net151 VGND VGND VPWR VPWR NN4BEG_outbuf_3.A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG2 net119 net19 net171 net223
+ Inst_LUT4AB_ConfigMem.ConfigBits\[414\] Inst_LUT4AB_ConfigMem.ConfigBits\[415\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG2 sky130_fd_sc_hd__mux4_1
X_031_ data_outbuf_31.X VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
X_100_ Inst_LUT4AB_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG0 net112 net12 net199 net216
+ Inst_LUT4AB_ConfigMem.ConfigBits\[418\] Inst_LUT4AB_ConfigMem.ConfigBits\[419\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_AB_BEG0 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix._041_ net20 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[496\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[497\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG3
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix._110_ Inst_LUT4AB_switch_matrix.JE2BEG2 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG2 sky130_fd_sc_hd__buf_1
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit8 net80 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[441\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_229_ W6BEG_outbuf_5.X VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4BEG_outbuf_10._0_ N4BEG_outbuf_10.A VGND VGND VPWR VPWR N4BEG_outbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit8 net80 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[360\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
Xinput205 SS4END[9] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xinput227 W6END[10] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
Xinput216 W2END[6] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_2
Xinput238 WW4END[0] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_2
Xinput249 WW4END[5] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr._12_ Inst_LH_LUT4c_frame_config_dffesr.I\[2\] VGND
+ VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._02_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst0 net105
+ net107 net7 net25 Inst_LUT4AB_ConfigMem.ConfigBits\[546\] Inst_LUT4AB_ConfigMem.ConfigBits\[547\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_014_ data_outbuf_14.X VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XS4END_inbuf_8._0_ net177 VGND VGND VPWR VPWR S4BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[305\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst0._0_ net528 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LD_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst0 net105 net5
+ net209 net543 Inst_LUT4AB_ConfigMem.ConfigBits\[229\] Inst_LUT4AB_ConfigMem.ConfigBits\[230\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst1 net512 net510
+ net509 net508 Inst_LUT4AB_ConfigMem.ConfigBits\[262\] Inst_LUT4AB_ConfigMem.ConfigBits\[263\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XEE4BEG_outbuf_9._0_ EE4BEG_outbuf_9.A VGND VGND VPWR VPWR EE4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG0 net131 net34 net183 Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[602\] Inst_LUT4AB_ConfigMem.ConfigBits\[603\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_GH_BEG0 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LB_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[568\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[569\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG5
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_118 E6BEG_outbuf_0.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 EE4BEG_outbuf_9.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit3 net75 net89 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput339 net339 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput317 net317 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst3 net509
+ net541 net540 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[478\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[479\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xoutput306 net306 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput328 net328 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_10._0_ net51 VGND VGND VPWR VPWR data_inbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[266\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[152\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG3 net107 net43 net159 net211
+ Inst_LUT4AB_ConfigMem.ConfigBits\[448\] Inst_LUT4AB_ConfigMem.ConfigBits\[449\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_GH_BEG3 sky130_fd_sc_hd__mux4_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit6 net78 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[443\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ SS4BEG_outbuf_5.X VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_18 N4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[532\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[533\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG4
+ sky130_fd_sc_hd__mux4_2
XANTENNA_29 S4BEG_outbuf_2.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit6 net78 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[365\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG2 net118 net170 net222
+ Inst_LUT4AB_switch_matrix.JS2BEG5 Inst_LUT4AB_ConfigMem.ConfigBits\[374\] Inst_LUT4AB_ConfigMem.ConfigBits\[375\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG2 net511 Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1
+ Inst_LUT4AB_switch_matrix.JE2BEG1 Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[214\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[215\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst1 net535 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ net539 Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[255\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[256\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
Xstrobe_outbuf_13._0_ strobe_inbuf_13.X VGND VGND VPWR VPWR strobe_outbuf_13.X sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_8._0_ data_inbuf_8.X VGND VGND VPWR VPWR data_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
Xinput27 E6END[3] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput38 EE4END[13] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput49 EE4END[9] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput16 E2MID[2] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
Xmax_cap508 Inst_LF_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__buf_6
X_245_ WW4BEG_outbuf_9.X VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_176_ S4BEG_outbuf_4.X VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG3 net115 net15 net167 net219
+ Inst_LUT4AB_ConfigMem.ConfigBits\[416\] Inst_LUT4AB_ConfigMem.ConfigBits\[417\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG3 sky130_fd_sc_hd__mux4_1
XWW4END_inbuf_4._0_ net252 VGND VGND VPWR VPWR WW4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_1
X_030_ data_outbuf_30.X VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._040_ net19 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb5
+ sky130_fd_sc_hd__buf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG1 net138 net8 net160 net212
+ Inst_LUT4AB_ConfigMem.ConfigBits\[420\] Inst_LUT4AB_ConfigMem.ConfigBits\[421\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_AB_BEG1 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame5_bit9 net81 net97 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[440\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame5_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_228_ W6BEG_outbuf_4.X VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkbuf_1
X_159_ Inst_LUT4AB_switch_matrix.S2BEG3 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame10_bit9 net81 net83 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[398\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame10_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput206 W1END[0] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__buf_4
XFILLER_0_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput217 W2END[7] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst1 net159
+ net181 net211 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[546\] Inst_LUT4AB_ConfigMem.ConfigBits\[547\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xinput228 W6END[11] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
Xinput239 WW4END[10] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr._11_ Inst_LH_LUT4c_frame_config_dffesr.I\[1\] VGND
+ VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr._01_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR._0_ sky130_fd_sc_hd__inv_2
X_013_ data_outbuf_13.X VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst1 Inst_LH_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2
+ Inst_LUT4AB_switch_matrix.J2END_EF_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[229\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[230\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst2 net511 net515
+ Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[262\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[263\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst0 net109
+ net131 net3 net9 Inst_LUT4AB_ConfigMem.ConfigBits\[458\] Inst_LUT4AB_ConfigMem.ConfigBits\[459\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_10._0_ net83 VGND VGND VPWR VPWR strobe_inbuf_10.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XE6END_inbuf_4._0_ net30 VGND VGND VPWR VPWR E6BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG1 net130 net198 net212 Inst_LUT4AB_switch_matrix.JE2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[604\] Inst_LUT4AB_ConfigMem.ConfigBits\[605\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_GH_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_41_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 E6BEG_outbuf_0.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 SS4BEG_outbuf_2.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit4 net76 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XSS4END_inbuf_6._0_ net191 VGND VGND VPWR VPWR SS4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput307 net307 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[480\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[481\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG7
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput318 net318 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput329 net329 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I0 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG0 Inst_LUT4AB_switch_matrix.J2END_CD_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[287\] Inst_LUT4AB_ConfigMem.ConfigBits\[288\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_8._0_ strobe_inbuf_8.X VGND VGND VPWR VPWR strobe_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN._0_ sky130_fd_sc_hd__inv_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH._0_ sky130_fd_sc_hd__inv_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XEE4END_inbuf_5._0_ net49 VGND VGND VPWR VPWR EE4BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit7 net79 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[518\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
X_192_ SS4BEG_outbuf_4.X VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_2._0_ net72 VGND VGND VPWR VPWR data_inbuf_2.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG0 net25 net160 net181 net543 Inst_LUT4AB_ConfigMem.ConfigBits\[218\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[219\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 N4BEG_outbuf_6.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XWW4BEG_outbuf_6._0_ WW4BEG_outbuf_6.A VGND VGND VPWR VPWR WW4BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit7 net79 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[373\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG3 net14 net166 net218 Inst_LUT4AB_switch_matrix.JW2BEG5
+ Inst_LUT4AB_ConfigMem.ConfigBits\[376\] Inst_LUT4AB_ConfigMem.ConfigBits\[377\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S1BEG3 Inst_LH_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 Inst_LUT4AB_switch_matrix.JE2BEG2 Inst_LUT4AB_switch_matrix.J_l_AB_BEG0
+ Inst_LUT4AB_ConfigMem.ConfigBits\[216\] Inst_LUT4AB_ConfigMem.ConfigBits\[217\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S1BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_244_ WW4BEG_outbuf_8.X VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XE6BEG_outbuf_9._0_ E6BEG_outbuf_9.A VGND VGND VPWR VPWR E6BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
Xinput28 E6END[4] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput39 EE4END[14] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput17 E2MID[3] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
Xmax_cap509 Inst_LE_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_6
X_175_ S4BEG_outbuf_3.X VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEF._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[153\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S sky130_fd_sc_hd__o21ai_2
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LF_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LA_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4END_inbuf_8._0_ net125 VGND VGND VPWR VPWR N4BEG_outbuf_8.A sky130_fd_sc_hd__buf_2
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XFILLER_0_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG2 net110 net34 net162 net214
+ Inst_LUT4AB_ConfigMem.ConfigBits\[422\] Inst_LUT4AB_ConfigMem.ConfigBits\[423\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_AB_BEG2 sky130_fd_sc_hd__mux4_2
Xoutput490 net490 VGND VGND VPWR VPWR W6BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_227_ W6BEG_outbuf_3.X VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XN4BEG_outbuf_0._0_ N4BEG_outbuf_0.A VGND VGND VPWR VPWR N4BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_089_ EE4BEG_outbuf_5.X VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkbuf_1
X_158_ Inst_LUT4AB_switch_matrix.S2BEG2 VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix._099_ net223 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb5
+ sky130_fd_sc_hd__buf_1
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput229 W6END[1] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__buf_4
Xinput207 W1END[1] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_4
Xinput218 W2MID[0] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst2 Inst_LB_LUT4c_frame_config_dffesr.O
+ net537 net510 net509 Inst_LUT4AB_ConfigMem.ConfigBits\[546\] Inst_LUT4AB_ConfigMem.ConfigBits\[547\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit2 net72 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[396\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[326\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._1_
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
X_012_ data_outbuf_12.X VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XW6BEG_outbuf_0._0_ W6BEG_outbuf_0.A VGND VGND VPWR VPWR W6BEG_outbuf_0.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I0 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG0
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0 Inst_LUT4AB_switch_matrix.J2END_EF_BEG0
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[317\] Inst_LUT4AB_ConfigMem.ConfigBits\[318\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.I\[0\] sky130_fd_sc_hd__mux4_1
XFILLER_0_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ net539 Inst_LUT4AB_ConfigMem.ConfigBits\[262\] Inst_LUT4AB_ConfigMem.ConfigBits\[263\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst1 net25 net161
+ net213 net245 Inst_LUT4AB_ConfigMem.ConfigBits\[458\] Inst_LUT4AB_ConfigMem.ConfigBits\[459\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.EH
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH_GH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG2 net25 net181 net247 Inst_LUT4AB_switch_matrix.JS2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[606\] Inst_LUT4AB_ConfigMem.ConfigBits\[607\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_GH_BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XNN4BEG_outbuf_9._0_ NN4BEG_outbuf_9.A VGND VGND VPWR VPWR NN4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst0 net103
+ net111 net3 net11 Inst_LUT4AB_ConfigMem.ConfigBits\[498\] Inst_LUT4AB_ConfigMem.ConfigBits\[499\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst0._0__520 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst0._0__520/HI
+ net520 sky130_fd_sc_hd__conb_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit2 net72 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[388\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_20._0_ data_inbuf_20.X VGND VGND VPWR VPWR data_outbuf_20.X sky130_fd_sc_hd__clkbuf_1
XANTENNA_109 W6BEG_outbuf_2.X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit5 net77 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_11._0_ data_inbuf_11.X VGND VGND VPWR VPWR data_outbuf_11.X sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_0._0_ S4BEG_outbuf_0.A VGND VGND VPWR VPWR S4BEG_outbuf_0.X sky130_fd_sc_hd__buf_2
XFILLER_0_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput319 net319 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput308 net308 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I1 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2END_CD_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[289\] Inst_LUT4AB_ConfigMem.ConfigBits\[290\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
XFILLER_0_22_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit8 net80 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[523\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
X_191_ SS4BEG_outbuf_3.X VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG0 net147 net183 net238 Inst_LUT4AB_switch_matrix.JN2BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[578\] Inst_LUT4AB_ConfigMem.ConfigBits\[579\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_AB_BEG0 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG1 net22 net161 net182 net532 Inst_LUT4AB_ConfigMem.ConfigBits\[220\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[221\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XNN4END_inbuf_6._0_ net139 VGND VGND VPWR VPWR NN4BEG_outbuf_6.A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XW6END_inbuf_2._0_ net232 VGND VGND VPWR VPWR W6BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit8 net80 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[409\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 E2MID[4] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
X_243_ WW4BEG_outbuf_7.X VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst0 net105
+ net113 net5 net13 Inst_LUT4AB_ConfigMem.ConfigBits\[570\] Inst_LUT4AB_ConfigMem.ConfigBits\[571\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEF._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[153\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._1_
+ sky130_fd_sc_hd__nand2_1
Xinput29 E6END[5] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
X_174_ S4BEG_outbuf_2.X VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG3 net106 net6 net158 net247
+ Inst_LUT4AB_ConfigMem.ConfigBits\[424\] Inst_LUT4AB_ConfigMem.ConfigBits\[425\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_AB_BEG3 sky130_fd_sc_hd__mux4_2
Xoutput491 net491 VGND VGND VPWR VPWR W6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput480 net480 VGND VGND VPWR VPWR W6BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_226_ W6BEG_outbuf_2.X VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkbuf_1
X_157_ Inst_LUT4AB_switch_matrix.S2BEG1 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_1
X_088_ EE4BEG_outbuf_4.X VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._098_ net222 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit0 net50 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[358\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG0 net121 net21 net173 net225
+ Inst_LUT4AB_ConfigMem.ConfigBits\[386\] Inst_LUT4AB_ConfigMem.ConfigBits\[387\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG0 sky130_fd_sc_hd__mux4_1
Xinput219 W2MID[1] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_2
Xinput208 W1END[2] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst3 Inst_LF_LUT4c_frame_config_dffesr.O
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.ConfigBits\[546\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[547\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[326\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._1_
+ sky130_fd_sc_hd__nand2_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_CD._4_ Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.CD sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit3 net75 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[412\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
X_011_ data_outbuf_11.X VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst0 net104
+ net112 net4 net12 Inst_LUT4AB_ConfigMem.ConfigBits\[534\] Inst_LUT4AB_ConfigMem.ConfigBits\[535\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I1 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1 Inst_LUT4AB_switch_matrix.J2END_EF_BEG1
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[319\] Inst_LUT4AB_ConfigMem.ConfigBits\[320\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.I\[1\] sky130_fd_sc_hd__mux4_2
X_209_ Inst_LUT4AB_switch_matrix.W2BEG1 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[264\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[265\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W6BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst2 net514
+ net513 net510 net509 Inst_LUT4AB_ConfigMem.ConfigBits\[458\] Inst_LUT4AB_ConfigMem.ConfigBits\[459\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_31._0_ net74 VGND VGND VPWR VPWR data_inbuf_31.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG3 net138 net22 net210 Inst_LUT4AB_switch_matrix.JW2BEG4
+ Inst_LUT4AB_ConfigMem.ConfigBits\[608\] Inst_LUT4AB_ConfigMem.ConfigBits\[609\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_GH_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LA_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_22._0_ net64 VGND VGND VPWR VPWR data_inbuf_22.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst1 net155
+ net157 net163 net207 Inst_LUT4AB_ConfigMem.ConfigBits\[498\] Inst_LUT4AB_ConfigMem.ConfigBits\[499\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit3 net75 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[386\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_inbuf_1._0_ net93 VGND VGND VPWR VPWR strobe_inbuf_1.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_13._0_ net54 VGND VGND VPWR VPWR data_inbuf_13.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit6 net78 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_63_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput309 net309 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I2 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG2 Inst_LUT4AB_switch_matrix.J2END_CD_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[291\] Inst_LUT4AB_ConfigMem.ConfigBits\[292\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
XWW4BEG_outbuf_10._0_ WW4BEG_outbuf_10.A VGND VGND VPWR VPWR WW4BEG_outbuf_10.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit20 net62 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[238\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ SS4BEG_outbuf_2.X VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit9 net81 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[539\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG2 net158 net183 net229 net512 Inst_LUT4AB_ConfigMem.ConfigBits\[222\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[223\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG2
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG1 net42 net182 net217 Inst_LUT4AB_switch_matrix.JE2BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[580\] Inst_LUT4AB_ConfigMem.ConfigBits\[581\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_AB_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_63_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_16._0_ strobe_inbuf_16.X VGND VGND VPWR VPWR strobe_outbuf_16.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit9 net81 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[407\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XWW4END_inbuf_7._0_ net240 VGND VGND VPWR VPWR WW4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 E2MID[5] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
X_173_ S4BEG_outbuf_1.X VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_1
X_242_ WW4BEG_outbuf_6.X VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst1 net155
+ net157 net165 net209 Inst_LUT4AB_ConfigMem.ConfigBits\[570\] Inst_LUT4AB_ConfigMem.ConfigBits\[571\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEF._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit30 net73 net91 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[294\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sCD.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.S0
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.AH
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_J_SR_BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
Xoutput470 net470 VGND VGND VPWR VPWR W2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput481 net481 VGND VGND VPWR VPWR W6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput492 net492 VGND VGND VPWR VPWR WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ EE4BEG_outbuf_3.X VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ W6BEG_outbuf_1.X VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_1
X_156_ Inst_LUT4AB_switch_matrix.S2BEG0 VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__buf_1
XFILLER_0_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix._097_ net221 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb3
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst0._0__524 VGND
+ VGND VPWR VPWR net524 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst0._0__524/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit1 net61 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[352\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput209 W1END[3] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_8
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG1 net117 net17 net169 net221
+ Inst_LUT4AB_ConfigMem.ConfigBits\[388\] Inst_LUT4AB_ConfigMem.ConfigBits\[389\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[548\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[549\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN._0_ sky130_fd_sc_hd__inv_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_CD._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN\[1\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit4 net76 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[405\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
X_010_ data_outbuf_10.X VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_13._0_ net86 VGND VGND VPWR VPWR strobe_inbuf_13.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst1 net156
+ net164 net206 net208 Inst_LUT4AB_ConfigMem.ConfigBits\[534\] Inst_LUT4AB_ConfigMem.ConfigBits\[535\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XE6END_inbuf_7._0_ net33 VGND VGND VPWR VPWR E6BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I2 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG2
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG2 Inst_LUT4AB_switch_matrix.J2END_EF_BEG2
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[321\] Inst_LUT4AB_ConfigMem.ConfigBits\[322\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.I\[2\] sky130_fd_sc_hd__mux4_2
X_139_ NN4BEG_outbuf_3.X VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst0 net104 net4
+ net156 net541 Inst_LUT4AB_ConfigMem.ConfigBits\[190\] Inst_LUT4AB_ConfigMem.ConfigBits\[191\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
X_208_ Inst_LUT4AB_switch_matrix.W2BEG0 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst0._0__519 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LD_SR.break_comb_loop_inst0._0__519/HI
+ net519 sky130_fd_sc_hd__conb_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[458\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[459\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4END_inbuf_9._0_ net194 VGND VGND VPWR VPWR SS4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit4 net76 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[422\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst2 net514
+ Inst_LB_LUT4c_frame_config_dffesr.O Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[498\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[499\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit7 net79 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XEE4END_inbuf_8._0_ net37 VGND VGND VPWR VPWR EE4BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_5._0_ net77 VGND VGND VPWR VPWR data_inbuf_5.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LC_I3 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 Inst_LUT4AB_switch_matrix.J2END_CD_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_CD_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[293\] Inst_LUT4AB_ConfigMem.ConfigBits\[294\]
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_2
XWW4BEG_outbuf_9._0_ WW4BEG_outbuf_9.A VGND VGND VPWR VPWR WW4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit10 net51 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[467\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit21 net63 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[258\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_S4BEG3 net159 net174 net226 Inst_LD_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_ConfigMem.ConfigBits\[224\] Inst_LUT4AB_ConfigMem.ConfigBits\[225\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG2 net129 net25 net229 Inst_LUT4AB_switch_matrix.JS2BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[582\] Inst_LUT4AB_ConfigMem.ConfigBits\[583\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_AB_BEG2 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst0._0__528 VGND
+ VGND VPWR VPWR net528 Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_EN.break_comb_loop_inst0._0__528/LO
+ sky130_fd_sc_hd__conb_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_172_ S4BEG_outbuf_0.X VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_1
X_241_ WW4BEG_outbuf_5.X VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst2 net514
+ net513 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[570\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[571\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4BEG_outbuf_3._0_ N4BEG_outbuf_3.A VGND VGND VPWR VPWR N4BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit20 net62 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit31 net74 net91 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[284\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XSS4BEG_outbuf_2._0_ SS4BEG_outbuf_2.A VGND VGND VPWR VPWR SS4BEG_outbuf_2.X sky130_fd_sc_hd__buf_2
XFILLER_0_64_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput482 net482 VGND VGND VPWR VPWR W6BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput460 net460 VGND VGND VPWR VPWR W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput471 net471 VGND VGND VPWR VPWR W2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput493 net493 VGND VGND VPWR VPWR WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
XSS4BEG_outbuf_10._0_ SS4BEG_outbuf_10.A VGND VGND VPWR VPWR SS4BEG_outbuf_10.X sky130_fd_sc_hd__buf_2
XFILLER_0_49_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_224_ W6BEG_outbuf_0.X VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_1
X_086_ EE4BEG_outbuf_2.X VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_1
X_155_ Inst_LUT4AB_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._096_ net220 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XW6BEG_outbuf_3._0_ W6BEG_outbuf_3.A VGND VGND VPWR VPWR W6BEG_outbuf_3.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit2 net72 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[363\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_CD._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_CD._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG2 net119 net19 net171 net223
+ Inst_LUT4AB_ConfigMem.ConfigBits\[390\] Inst_LUT4AB_ConfigMem.ConfigBits\[391\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG2 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit5 net77 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[404\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sEF.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.S0
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sEF.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst2 net514
+ net513 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[534\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[535\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
Xoutput290 net290 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit30 net73 net90 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[295\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst1 net540 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2END_GH_BEG0
+ Inst_LUT4AB_ConfigMem.ConfigBits\[190\] Inst_LUT4AB_ConfigMem.ConfigBits\[191\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_LF_I3 Inst_LUT4AB_switch_matrix.J2MID_EFa_BEG3
+ Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG3 Inst_LUT4AB_switch_matrix.J2END_EF_BEG3
+ Inst_LUT4AB_switch_matrix.J_l_EF_BEG3 Inst_LUT4AB_ConfigMem.ConfigBits\[323\] Inst_LUT4AB_ConfigMem.ConfigBits\[324\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.I\[3\] sky130_fd_sc_hd__mux4_1
X_207_ Inst_LUT4AB_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_1
X_069_ strobe_outbuf_5.X VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkbuf_1
X_138_ NN4BEG_outbuf_2.X VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix._079_ net167 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb1
+ sky130_fd_sc_hd__clkbuf_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst0 net102 net2
+ net206 net513 Inst_LUT4AB_ConfigMem.ConfigBits\[176\] Inst_LUT4AB_ConfigMem.ConfigBits\[177\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst0 net5 net209
+ net514 net513 Inst_LUT4AB_ConfigMem.ConfigBits\[202\] Inst_LUT4AB_ConfigMem.ConfigBits\[203\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[460\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[461\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_outbuf_23._0_ data_inbuf_23.X VGND VGND VPWR VPWR data_outbuf_23.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_outbuf_14._0_ data_inbuf_14.X VGND VGND VPWR VPWR data_outbuf_14.X sky130_fd_sc_hd__clkbuf_1
XInst_LA_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LA_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XS4BEG_outbuf_3._0_ S4BEG_outbuf_3.A VGND VGND VPWR VPWR S4BEG_outbuf_3.X sky130_fd_sc_hd__buf_2
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit5 net77 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[463\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst3 net508
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[498\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[499\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit8 net80 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XS4END_inbuf_1._0_ net185 VGND VGND VPWR VPWR S4BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsplit1 Inst_LB_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__buf_6
XFILLER_0_42_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[315\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._1_
+ VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.SR sky130_fd_sc_hd__o21ai_1
XNN4END_inbuf_9._0_ net142 VGND VGND VPWR VPWR NN4BEG_outbuf_9.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XEE4BEG_outbuf_2._0_ EE4BEG_outbuf_2.A VGND VGND VPWR VPWR EE4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XW6END_inbuf_5._0_ net235 VGND VGND VPWR VPWR W6BEG_outbuf_5.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit22 net64 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[254\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit11 net52 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[575\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG3 net122 net22 net174 Inst_LUT4AB_switch_matrix.JW2BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[584\] Inst_LUT4AB_ConfigMem.ConfigBits\[585\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J_l_AB_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput190 SS4END[0] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit0 net50 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[340\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_240_ WW4BEG_outbuf_4.X VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst3 net509
+ Inst_LF_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[570\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[571\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_171_ Inst_LUT4AB_switch_matrix.S2BEGb7 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit0 net50 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[327\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xrebuffer1 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__dlygate4sd1_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit21 net63 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.break_comb_loop_inst0._0_ net524 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LA_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit10 net51 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput483 net483 VGND VGND VPWR VPWR W6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput450 net450 VGND VGND VPWR VPWR SS4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput461 net461 VGND VGND VPWR VPWR W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput472 net472 VGND VGND VPWR VPWR W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput494 net494 VGND VGND VPWR VPWR WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_223_ Inst_LUT4AB_switch_matrix.W2BEGb7 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ EE4BEG_outbuf_1.X VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkbuf_1
X_154_ Inst_LUT4AB_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[276\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._1_
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_switch_matrix._095_ net219 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst1._0_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit3 net75 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[375\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG3 net115 net15 net167 net219
+ Inst_LUT4AB_ConfigMem.ConfigBits\[392\] Inst_LUT4AB_ConfigMem.ConfigBits\[393\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG3 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit6 net78 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[479\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_outbuf_1._0_ data_inbuf_1.X VGND VGND VPWR VPWR data_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst3 net509
+ Inst_LG_LUT4c_frame_config_dffesr.O net515 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[534\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[535\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xoutput280 net280 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput291 net291 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit20 net62 net90 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit31 net74 net90 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[285\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
X_137_ NN4BEG_outbuf_1.X VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_206_ Inst_LUT4AB_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_068_ strobe_outbuf_4.X VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix._078_ net166 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.S2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst1 net537 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_switch_matrix.J2END_CD_BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[176\] Inst_LUT4AB_ConfigMem.ConfigBits\[177\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_25._0_ net67 VGND VGND VPWR VPWR data_inbuf_25.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst1 net537 net510
+ net509 net541 Inst_LUT4AB_ConfigMem.ConfigBits\[202\] Inst_LUT4AB_ConfigMem.ConfigBits\[203\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_4._0_ net96 VGND VGND VPWR VPWR strobe_inbuf_4.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_16._0_ net57 VGND VGND VPWR VPWR data_inbuf_16.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LA_LUT4c_frame_config_dffesr._20_ Inst_LA_LUT4c_frame_config_dffesr._06_ Inst_LA_LUT4c_frame_config_dffesr._07_
+ Inst_LA_LUT4c_frame_config_dffesr._08_ Inst_LA_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_sGH.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.S
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sGH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[500\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[501\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JE2BEG4
+ sky130_fd_sc_hd__mux4_2
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit9 net81 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit30 net73 net89 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[283\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_outbuf_19._0_ strobe_inbuf_19.X VGND VGND VPWR VPWR strobe_outbuf_19.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst0 net102
+ net108 net8 net22 Inst_LUT4AB_ConfigMem.ConfigBits\[550\] Inst_LUT4AB_ConfigMem.ConfigBits\[551\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[315\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit23 net65 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[253\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit12 net53 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[574\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst0 net102 net2
+ net206 net532 Inst_LUT4AB_ConfigMem.ConfigBits\[232\] Inst_LUT4AB_ConfigMem.ConfigBits\[233\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput180 S4END[15] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput191 SS4END[10] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit1 net61 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[385\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_170_ Inst_LUT4AB_switch_matrix.S2BEGb6 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[572\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[573\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG6
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_1._0_ strobe_inbuf_1.X VGND VGND VPWR VPWR strobe_outbuf_1.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit1 net61 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[297\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
Xrebuffer2 Inst_LUT4AB_switch_matrix.JW2BEG5 VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__buf_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit22 net64 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit11 net52 net91 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst0 net145
+ net5 net7 net25 Inst_LUT4AB_ConfigMem.ConfigBits\[514\] Inst_LUT4AB_ConfigMem.ConfigBits\[515\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.break_comb_loop_inst0._0_ net520 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput484 net484 VGND VGND VPWR VPWR W6BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput495 net495 VGND VGND VPWR VPWR WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput451 net451 VGND VGND VPWR VPWR SS4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput440 net440 VGND VGND VPWR VPWR S4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput462 net462 VGND VGND VPWR VPWR W1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput473 net473 VGND VGND VPWR VPWR W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_153_ Inst_LUT4AB_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[276\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix._094_ net218 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
X_222_ Inst_LUT4AB_switch_matrix.W2BEGb6 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_16._0_ net89 VGND VGND VPWR VPWR strobe_inbuf_16.X sky130_fd_sc_hd__clkbuf_1
X_084_ EE4BEG_outbuf_0.X VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_AB.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.B
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_AB.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit4 net76 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[371\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LB_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit7 net79 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[478\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[536\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[537\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG5
+ sky130_fd_sc_hd__mux4_2
Xoutput270 net270 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput281 net281 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__clkbuf_4
XE6BEG_outbuf_2._0_ E6BEG_outbuf_2.A VGND VGND VPWR VPWR E6BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
Xoutput292 net292 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit21 net63 net90 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit10 net51 net90 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
X_136_ NN4BEG_outbuf_0.X VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix._077_ Inst_LUT4AB_switch_matrix.JS2BEG7 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG7 sky130_fd_sc_hd__clkbuf_1
X_205_ Inst_LUT4AB_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_067_ strobe_outbuf_3.X VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__clkbuf_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XN4END_inbuf_1._0_ net133 VGND VGND VPWR VPWR N4BEG_outbuf_1.A sky130_fd_sc_hd__buf_2
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst2 net540 net515
+ net542 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[202\] Inst_LUT4AB_ConfigMem.ConfigBits\[203\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_inbuf_8._0_ net80 VGND VGND VPWR VPWR data_inbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_119_ Inst_LUT4AB_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit7 net79 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[480\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit20 net62 net89 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit31 net74 net89 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[274\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._4_ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.I0mux sky130_fd_sc_hd__o21ai_4
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst1 net160
+ net182 net212 net226 Inst_LUT4AB_ConfigMem.ConfigBits\[550\] Inst_LUT4AB_ConfigMem.ConfigBits\[551\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LE_SR._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit13 net54 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[567\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit24 net66 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[252\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst1 net512 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_switch_matrix.J2END_CD_BEG3
+ Inst_LUT4AB_ConfigMem.ConfigBits\[232\] Inst_LUT4AB_ConfigMem.ConfigBits\[233\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[257\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o21ai_1
Xinput181 S4END[1] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xinput170 S2MID[4] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_4
Xinput192 SS4END[11] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst0 net110
+ net122 net4 net10 Inst_LUT4AB_ConfigMem.ConfigBits\[462\] Inst_LUT4AB_ConfigMem.ConfigBits\[463\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XNN4BEG_outbuf_2._0_ NN4BEG_outbuf_2.A VGND VGND VPWR VPWR NN4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_1
XN4BEG_outbuf_6._0_ N4BEG_outbuf_6.A VGND VGND VPWR VPWR N4BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.break_comb_loop_inst0._0_ net529 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_EN.AIN\[0\] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit30 net73 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[279\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit2 net72 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[415\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4BEG_outbuf_5._0_ SS4BEG_outbuf_5.A VGND VGND VPWR VPWR SS4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_2
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[181\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.NN4BEG3 sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit2 net72 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[337\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit12 net53 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
Xrebuffer3 net536 VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__buf_6
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit23 net65 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[13\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[201\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.EE4BEG3 sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst1 net159
+ net181 net211 net229 Inst_LUT4AB_ConfigMem.ConfigBits\[514\] Inst_LUT4AB_ConfigMem.ConfigBits\[515\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XW6BEG_outbuf_6._0_ W6BEG_outbuf_6.A VGND VGND VPWR VPWR W6BEG_outbuf_6.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput452 net452 VGND VGND VPWR VPWR SS4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput441 net441 VGND VGND VPWR VPWR S4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput430 net430 VGND VGND VPWR VPWR S4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput485 net485 VGND VGND VPWR VPWR W6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput496 net496 VGND VGND VPWR VPWR WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput463 net463 VGND VGND VPWR VPWR W1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput474 net474 VGND VGND VPWR VPWR W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_083_ strobe_outbuf_19.X VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ Inst_LUT4AB_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_EN._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix._093_ Inst_LUT4AB_switch_matrix.JW2BEG7 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG7 sky130_fd_sc_hd__clkbuf_1
X_221_ Inst_LUT4AB_switch_matrix.W2BEGb5 VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LH_LUT4c_frame_config_dffesr.I0mux
+ Inst_LH_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit5 net77 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[370\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr._20_ Inst_LB_LUT4c_frame_config_dffesr._06_ Inst_LB_LUT4c_frame_config_dffesr._07_
+ Inst_LB_LUT4c_frame_config_dffesr._08_ Inst_LB_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit8 net80 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[471\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_26._0_ data_inbuf_26.X VGND VGND VPWR VPWR data_outbuf_26.X sky130_fd_sc_hd__clkbuf_1
Xoutput282 net282 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput293 net293 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput271 net271 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput260 net260 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit22 net64 net90 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit11 net52 net90 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_204_ Inst_LUT4AB_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_1
X_066_ strobe_outbuf_2.X VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_1
X_135_ Inst_LUT4AB_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._076_ Inst_LUT4AB_switch_matrix.JS2BEG6 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG6 sky130_fd_sc_hd__buf_1
XFILLER_0_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_17._0_ data_inbuf_17.X VGND VGND VPWR VPWR data_outbuf_17.X sky130_fd_sc_hd__clkbuf_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XS4BEG_outbuf_6._0_ S4BEG_outbuf_6.A VGND VGND VPWR VPWR S4BEG_outbuf_6.X sky130_fd_sc_hd__buf_2
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix.J2MID_ABb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG1 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG1
+ Inst_LUT4AB_switch_matrix.J2MID_GHb_BEG1 Inst_LUT4AB_ConfigMem.ConfigBits\[202\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[203\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_CD.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.D
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XS4END_inbuf_4._0_ net188 VGND VGND VPWR VPWR S4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_118_ Inst_LUT4AB_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._059_ Inst_LUT4AB_switch_matrix.JN2BEG5 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG5 sky130_fd_sc_hd__buf_1
X_049_ E6BEG_outbuf_9.X VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit8 net80 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[504\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit21 net63 net89 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit10 net51 net89 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XEE4BEG_outbuf_5._0_ EE4BEG_outbuf_5.A VGND VGND VPWR VPWR EE4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XW6END_inbuf_8._0_ net227 VGND VGND VPWR VPWR W6BEG_outbuf_8.A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._3_ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\]
+ Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[17\] VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit4 Inst_LE_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__buf_6
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[336\]
+ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._0_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._1_
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.EN sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.A0 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit0 net50 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[301\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XANTENNA_1 E6BEG_outbuf_3.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst2 net514
+ net512 net510 Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[550\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[551\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit14 net55 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[566\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit25 net67 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[246\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH._4_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.EH sky130_fd_sc_hd__o21ai_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[257\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
Xinput182 S4END[2] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_2
Xinput160 S2END[2] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
Xinput171 S2MID[5] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xinput193 SS4END[12] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit20 net62 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst1 net22 net162
+ net214 net226 Inst_LUT4AB_ConfigMem.ConfigBits\[462\] Inst_LUT4AB_ConfigMem.ConfigBits\[463\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LG_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit31 net74 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[275\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit3 net75 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[402\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[181\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LC_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LC_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst0 net104
+ net112 net4 net12 Inst_LUT4AB_ConfigMem.ConfigBits\[502\] Inst_LUT4AB_ConfigMem.ConfigBits\[503\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit13 net54 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[9\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
Xrebuffer4 Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlymetal6s2s_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit24 net66 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit3 net75 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[333\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[201\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst2 Inst_LB_LUT4c_frame_config_dffesr.O
+ net512 Inst_LD_LUT4c_frame_config_dffesr.O Inst_LE_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[514\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[515\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput486 net486 VGND VGND VPWR VPWR W6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput431 net431 VGND VGND VPWR VPWR S4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput453 net453 VGND VGND VPWR VPWR SS4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput442 net442 VGND VGND VPWR VPWR S4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput420 net420 VGND VGND VPWR VPWR S2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput464 net464 VGND VGND VPWR VPWR W2BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput475 net475 VGND VGND VPWR VPWR W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XSS4END_inbuf_11._0_ net196 VGND VGND VPWR VPWR SS4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_1
Xoutput497 net497 VGND VGND VPWR VPWR WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_220_ Inst_LUT4AB_switch_matrix.W2BEGb4 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_1
X_082_ strobe_outbuf_18.X VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkbuf_1
X_151_ Inst_LUT4AB_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix._092_ Inst_LUT4AB_switch_matrix.JW2BEG6 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG6 sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst1 Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[5\] Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[7\] Inst_LH_LUT4c_frame_config_dffesr.I0mux
+ Inst_LH_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xdata_outbuf_4._0_ data_inbuf_4.X VGND VGND VPWR VPWR data_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit30 net73 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[278\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG0 net120 net20 net172 Inst_LUT4AB_switch_matrix.JN2BEG6
+ Inst_LUT4AB_ConfigMem.ConfigBits\[378\] Inst_LUT4AB_ConfigMem.ConfigBits\[379\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit6 net78 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[428\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_28._0_ net70 VGND VGND VPWR VPWR data_inbuf_28.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit9 net81 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[470\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XWW4END_inbuf_0._0_ net248 VGND VGND VPWR VPWR WW4BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LB_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
Xoutput283 net283 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput294 net294 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__buf_2
Xoutput272 net272 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput261 net261 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__buf_2
Xstrobe_inbuf_7._0_ net99 VGND VGND VPWR VPWR strobe_inbuf_7.X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_19._0_ net60 VGND VGND VPWR VPWR data_inbuf_19.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit12 net53 net90 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit23 net65 net90 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_203_ Inst_LUT4AB_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_1
X_065_ strobe_outbuf_1.X VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_1
X_134_ Inst_LUT4AB_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix._075_ Inst_LUT4AB_switch_matrix.JS2BEG5 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG5 sky130_fd_sc_hd__buf_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[204\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[205\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E6BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst0 net102
+ net138 net2 net6 Inst_LUT4AB_ConfigMem.ConfigBits\[574\] Inst_LUT4AB_ConfigMem.ConfigBits\[575\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ Inst_LUT4AB_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix._058_ Inst_LUT4AB_switch_matrix.JN2BEG4 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG4 sky130_fd_sc_hd__clkbuf_1
X_048_ E6BEG_outbuf_8.X VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkbuf_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame1_bit9 net81 net93 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[527\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame1_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit22 net64 net89 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit11 net52 net89 VGND VGND VPWR VPWR Inst_LA_LUT4c_frame_config_dffesr.ConfigBits\[18\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_EF.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.F
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EF.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._2_ Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux._0_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit30 net73 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[603\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XE6END_inbuf_0._0_ net26 VGND VGND VPWR VPWR E6BEG_outbuf_0.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsplit5 Inst_LG_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__buf_4
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._3_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[336\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit1 net61 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[300\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LG_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_2 E6BEG_outbuf_3.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[550\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[551\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst0 net105
+ net113 net5 net13 Inst_LUT4AB_ConfigMem.ConfigBits\[538\] Inst_LUT4AB_ConfigMem.ConfigBits\[539\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit15 net56 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[562\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4END_inbuf_2._0_ net202 VGND VGND VPWR VPWR SS4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_1
XEE4END_inbuf_11._0_ net40 VGND VGND VPWR VPWR EE4BEG_outbuf_11.A sky130_fd_sc_hd__clkbuf_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN\[1\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.S VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput183 S4END[3] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__buf_2
Xinput194 SS4END[13] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
Xinput172 S2MID[6] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xinput161 S2END[3] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit21 net63 net88 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst2 net514
+ Inst_LB_LUT4c_frame_config_dffesr.O net512 net509 Inst_LUT4AB_ConfigMem.ConfigBits\[462\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[463\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
Xinput150 NN4END[6] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit10 net51 net88 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_4._0_ strobe_inbuf_4.X VGND VGND VPWR VPWR strobe_outbuf_4.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit4 net76 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[442\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
XEE4END_inbuf_1._0_ net45 VGND VGND VPWR VPWR EE4BEG_outbuf_1.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LC_LUT4c_frame_config_dffesr._20_ Inst_LC_LUT4c_frame_config_dffesr._06_ Inst_LC_LUT4c_frame_config_dffesr._07_
+ Inst_LC_LUT4c_frame_config_dffesr._08_ Inst_LC_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit4 net76 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[342\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst1 net154
+ net156 net164 net208 Inst_LUT4AB_ConfigMem.ConfigBits\[502\] Inst_LUT4AB_ConfigMem.ConfigBits\[503\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XWW4BEG_outbuf_2._0_ WW4BEG_outbuf_2.A VGND VGND VPWR VPWR WW4BEG_outbuf_2.X sky130_fd_sc_hd__clkbuf_2
Xstrobe_inbuf_19._0_ net92 VGND VGND VPWR VPWR strobe_inbuf_19.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit14 net55 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux21_inst._0_
+ sky130_fd_sc_hd__inv_2
Xrebuffer5 Inst_LUT4AB_switch_matrix.S0 VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit25 net67 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.ConfigBits\[514\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[515\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput487 net487 VGND VGND VPWR VPWR W6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput498 net498 VGND VGND VPWR VPWR WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput454 net454 VGND VGND VPWR VPWR SS4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput443 net443 VGND VGND VPWR VPWR SS4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput432 net432 VGND VGND VPWR VPWR S4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput410 net410 VGND VGND VPWR VPWR S1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput421 net421 VGND VGND VPWR VPWR S2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput465 net465 VGND VGND VPWR VPWR W2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput476 net476 VGND VGND VPWR VPWR W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
X_150_ Inst_LUT4AB_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_EN_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LC_EN.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_081_ strobe_outbuf_17.X VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit20 net62 net87 VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix._091_ net533 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.W2BEG5
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit31 net74 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[614\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst2 Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[8\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[9\] Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[11\] Inst_LH_LUT4c_frame_config_dffesr.I0mux
+ Inst_LH_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XE6BEG_outbuf_5._0_ E6BEG_outbuf_5.A VGND VGND VPWR VPWR E6BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG1 net116 net168 net220
+ Inst_LUT4AB_switch_matrix.JE2BEG6 Inst_LUT4AB_ConfigMem.ConfigBits\[380\] Inst_LUT4AB_ConfigMem.ConfigBits\[381\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit7 net79 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[455\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XN4END_inbuf_4._0_ net136 VGND VGND VPWR VPWR N4BEG_outbuf_4.A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_sCD._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[152\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._1_
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_CD.S sky130_fd_sc_hd__o21ai_1
Xoutput284 net284 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput295 net295 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput273 net273 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput262 net262 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit13 net54 net90 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit24 net66 net90 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
X_133_ Inst_LUT4AB_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._074_ Inst_LUT4AB_switch_matrix.JS2BEG4 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG4 sky130_fd_sc_hd__buf_1
X_202_ Inst_LUT4AB_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_1
X_064_ strobe_outbuf_0.X VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkbuf_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._4_ Inst_LUT4AB_ConfigMem.ConfigBits\[153\]
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._0_ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._1_
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_AH sky130_fd_sc_hd__o21ai_4
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.break_comb_loop_inst0._0_ Inst_LB_LUT4c_frame_config_dffesr.LUT_out
+ VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst1 net154
+ net156 net158 net206 Inst_LUT4AB_ConfigMem.ConfigBits\[574\] Inst_LUT4AB_ConfigMem.ConfigBits\[575\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit30 net73 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[611\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG0 Inst_LD_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_switch_matrix.J2MID_CDb_BEG3 Inst_LUT4AB_switch_matrix.JN2BEG3 Inst_LUT4AB_switch_matrix.J_l_CD_BEG1
+ Inst_LUT4AB_ConfigMem.ConfigBits\[182\] Inst_LUT4AB_ConfigMem.ConfigBits\[183\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_116_ Inst_LUT4AB_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._057_ Inst_LUT4AB_switch_matrix.JN2BEG3 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG3 sky130_fd_sc_hd__clkbuf_2
X_047_ E6BEG_outbuf_7.X VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkbuf_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit12 net53 net89 VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.break_comb_loop_inst1._0_ Inst_MUX8LUT_frame_config_mux.AD
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AD.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit23 net65 net89 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._4_ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._0_ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.O sky130_fd_sc_hd__o21ai_4
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit20 net62 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[579\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit31 net74 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[599\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsplit6 Inst_LC_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__buf_6
XFILLER_0_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._2_ Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LH_EN._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit2 net72 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[319\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr._21_ UserCLK Inst_LD_LUT4c_frame_config_dffesr._04_
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.LUT_flop sky130_fd_sc_hd__dfxtp_1
XANTENNA_3 EE4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._109_ Inst_LUT4AB_switch_matrix.JE2BEG1 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG1 sky130_fd_sc_hd__buf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[552\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[553\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JW2BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_21_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XNN4BEG_outbuf_5._0_ NN4BEG_outbuf_5.A VGND VGND VPWR VPWR NN4BEG_outbuf_5.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit16 net57 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[156\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XN4BEG_outbuf_9._0_ N4BEG_outbuf_9.A VGND VGND VPWR VPWR N4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst1 net157
+ net165 net207 net209 Inst_LUT4AB_ConfigMem.ConfigBits\[538\] Inst_LUT4AB_ConfigMem.ConfigBits\[539\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XSS4BEG_outbuf_8._0_ SS4BEG_outbuf_8.A VGND VGND VPWR VPWR SS4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst0 net105 net5
+ net157 net543 Inst_LUT4AB_ConfigMem.ConfigBits\[193\] Inst_LUT4AB_ConfigMem.ConfigBits\[194\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux.cus_mux21_GH.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.H
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_GH.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
Xinput162 S2END[4] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
XInst_MUX8LUT_frame_config_mux.cus_mux21_EH._2_ Inst_MUX8LUT_frame_config_mux.cus_mux21_EH.AIN\[0\]
+ VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_EH._0_ sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst3 net508
+ net511 net515 Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.ConfigBits\[462\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[463\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xinput151 NN4END[7] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xinput140 NN4END[11] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xinput184 S4END[4] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xinput173 S2MID[7] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_2
Xinput195 SS4END[14] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit22 net64 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[17\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit11 net52 net88 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit5 net77 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[435\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit30 net73 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[598\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XW6BEG_outbuf_9._0_ W6BEG_outbuf_9.A VGND VGND VPWR VPWR W6BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_2
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst0 Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[0\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[1\] Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[2\]
+ Inst_LG_LUT4c_frame_config_dffesr.ConfigBits\[3\] Inst_LG_LUT4c_frame_config_dffesr.I0mux
+ Inst_LG_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit15 net56 net91 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[16\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit5 net77 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[362\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst2 net514
+ net513 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[502\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[503\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit26 net68 net91 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[10\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[516\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[517\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JS2BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_64_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XNN4END_inbuf_2._0_ net150 VGND VGND VPWR VPWR NN4BEG_outbuf_2.A sky130_fd_sc_hd__clkbuf_2
Xoutput400 net400 VGND VGND VPWR VPWR NN4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput411 net411 VGND VGND VPWR VPWR S2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput488 net488 VGND VGND VPWR VPWR W6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput433 net433 VGND VGND VPWR VPWR S4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput422 net422 VGND VGND VPWR VPWR S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput444 net444 VGND VGND VPWR VPWR SS4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput455 net455 VGND VGND VPWR VPWR SS4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput466 net466 VGND VGND VPWR VPWR W2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput499 net499 VGND VGND VPWR VPWR WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput477 net477 VGND VGND VPWR VPWR W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
X_080_ strobe_outbuf_16.X VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.break_comb_loop_inst1._0_ Inst_LUT4AB_switch_matrix.J_SR_BEG0
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LG_SR.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix._090_ Inst_LUT4AB_switch_matrix.JW2BEG4 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.W2BEG4 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_29._0_ data_inbuf_29.X VGND VGND VPWR VPWR data_outbuf_29.X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit21 net63 net87 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[11\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame14_bit10 net51 net87 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[357\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame14_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_inst3 Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[12\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[13\] Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[14\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[15\] Inst_LH_LUT4c_frame_config_dffesr.I0mux
+ Inst_LH_LUT4c_frame_config_dffesr.I\[1\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG2 net18 net170 net222 Inst_LUT4AB_switch_matrix.JS2BEG6
+ Inst_LUT4AB_ConfigMem.ConfigBits\[382\] Inst_LUT4AB_ConfigMem.ConfigBits\[383\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2MID_GHa_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_51_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame4_bit8 net80 net96 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[452\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame4_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst1._0_ Inst_LF_LUT4c_frame_config_dffesr.Ci
+ VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[1\] sky130_fd_sc_hd__clkbuf_1
XS4BEG_outbuf_9._0_ S4BEG_outbuf_9.A VGND VGND VPWR VPWR S4BEG_outbuf_9.X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_MUX8LUT_frame_config_mux.cus_mux21_sCD._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[152\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_sCD._1_
+ sky130_fd_sc_hd__nand2_1
Xoutput285 net285 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput296 net296 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput263 net263 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_0_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit14 net55 net90 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[6\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem.Inst_Frame17_bit25 net67 net90 VGND VGND VPWR VPWR Inst_LE_LUT4c_frame_config_dffesr.ConfigBits\[7\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame17_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
X_132_ Inst_LUT4AB_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG0 net147 net12 net164 net216
+ Inst_LUT4AB_ConfigMem.ConfigBits\[426\] Inst_LUT4AB_ConfigMem.ConfigBits\[427\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.J2END_CD_BEG0 sky130_fd_sc_hd__mux4_2
X_063_ Inst_LUT4AB_switch_matrix.E2BEG7 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._073_ Inst_LUT4AB_switch_matrix.JS2BEG3 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.S2BEG3 sky130_fd_sc_hd__buf_1
X_201_ Inst_LUT4AB_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_1
XS4END_inbuf_7._0_ net176 VGND VGND VPWR VPWR S4BEG_outbuf_7.A sky130_fd_sc_hd__clkbuf_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._3_ Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH.AIN\[1\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[153\] VGND VGND VPWR VPWR Inst_MUX8LUT_frame_config_mux.cus_mux21_M_AH._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.break_comb_loop_inst0._0_ Inst_LD_LUT4c_frame_config_dffesr.I\[0\]
+ VGND VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr.cus_mux21_I0mux.AIN\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem.Inst_Frame18_bit0 net50 net91 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[324\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame18_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit20 net62 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[190\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame13_bit31 net74 net86 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[595\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame13_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst2 net543
+ net532 net512 Inst_LD_LUT4c_frame_config_dffesr.O Inst_LUT4AB_ConfigMem.ConfigBits\[574\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[575\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix.inst_cus_mux41_buf_E1BEG1 net535 Inst_LUT4AB_switch_matrix.J2MID_EFb_BEG0
+ Inst_LUT4AB_switch_matrix.JN2BEG0 Inst_LUT4AB_switch_matrix.J_l_EF_BEG2 Inst_LUT4AB_ConfigMem.ConfigBits\[184\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[185\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E1BEG1
+ sky130_fd_sc_hd__mux4_1
XEE4BEG_outbuf_8._0_ EE4BEG_outbuf_8.A VGND VGND VPWR VPWR EE4BEG_outbuf_8.X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_115_ Inst_LUT4AB_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
X_046_ E6BEG_outbuf_6.X VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix._056_ Inst_LUT4AB_switch_matrix.JN2BEG2 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.N2BEG2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux.cus_mux21_AB._4_ net534 Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._0_
+ Inst_MUX8LUT_frame_config_mux.cus_mux21_AB._1_ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.M_AB
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit13 net54 net89 VGND VGND VPWR VPWR Inst_LC_LUT4c_frame_config_dffesr.ConfigBits\[5\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame16_bit24 net66 net89 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[1\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame16_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._3_ Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O.AIN\[1\]
+ Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[16\] VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.cus_mux21_O._1_
+ sky130_fd_sc_hd__nand2_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit21 net63 net101 VGND VGND VPWR VPWR Inst_LH_LUT4c_frame_config_dffesr.ConfigBits\[3\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame9_bit10 net51 net101 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[361\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame9_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsplit7 Inst_LF_LUT4c_frame_config_dffesr.O VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__buf_6
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem.Inst_Frame0_bit0 net50 net82 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[389\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame0_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit3 net75 net88 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[317\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_029_ data_outbuf_29.X VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkbuf_1
XInst_LD_LUT4c_frame_config_dffesr._20_ Inst_LD_LUT4c_frame_config_dffesr._06_ Inst_LD_LUT4c_frame_config_dffesr._07_
+ Inst_LD_LUT4c_frame_config_dffesr._08_ Inst_LD_LUT4c_frame_config_dffesr._09_ VGND
+ VGND VPWR VPWR Inst_LD_LUT4c_frame_config_dffesr._04_ sky130_fd_sc_hd__a22oi_1
XANTENNA_4 EE4BEG_outbuf_10.A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem.Inst_Frame12_bit30 net73 net85 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[586\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame12_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix._039_ net18 VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.E2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst0._0__521 VGND
+ VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux21_LF_SR.break_comb_loop_inst0._0__521/HI
+ net521 sky130_fd_sc_hd__conb_1
XFILLER_0_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix._108_ Inst_LUT4AB_switch_matrix.JE2BEG0 VGND VGND VPWR
+ VPWR Inst_LUT4AB_switch_matrix.E2BEG0 sky130_fd_sc_hd__clkbuf_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem.Inst_Frame19_bit17 net58 net92 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[155\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame19_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst2 net514
+ net513 Inst_LC_LUT4c_frame_config_dffesr.O net510 Inst_LUT4AB_ConfigMem.ConfigBits\[538\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[539\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst1 Inst_LH_LUT4c_frame_config_dffesr.O
+ Inst_LUT4AB_switch_matrix.J2MID_ABa_BEG2 Inst_LUT4AB_switch_matrix.J2MID_CDa_BEG2
+ Inst_LUT4AB_switch_matrix.J2END_EF_BEG0 Inst_LUT4AB_ConfigMem.ConfigBits\[193\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[194\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux21_inst.A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst0 net103 net3
+ net207 net510 Inst_LUT4AB_ConfigMem.ConfigBits\[179\] Inst_LUT4AB_ConfigMem.ConfigBits\[180\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux21_inst.A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput185 S4END[5] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xinput174 S4END[0] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__buf_2
Xinput163 S2END[5] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_2
Xinput196 SS4END[15] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst0 net4 net208
+ net514 net513 Inst_LUT4AB_ConfigMem.ConfigBits\[206\] Inst_LUT4AB_ConfigMem.ConfigBits\[207\]
+ VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1 Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2
+ Inst_LUT4AB_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3 Inst_LUT4AB_ConfigMem.ConfigBits\[464\]
+ Inst_LUT4AB_ConfigMem.ConfigBits\[465\] VGND VGND VPWR VPWR Inst_LUT4AB_switch_matrix.JN2BEG3
+ sky130_fd_sc_hd__mux4_2
Xinput152 NN4END[8] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xinput141 NN4END[12] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
Xinput130 N4END[2] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__buf_2
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit23 net65 net88 VGND VGND VPWR VPWR Inst_LF_LUT4c_frame_config_dffesr.ConfigBits\[15\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame15_bit12 net53 net88 VGND VGND VPWR VPWR Inst_LB_LUT4c_frame_config_dffesr.ConfigBits\[4\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame15_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame7_bit6 net78 net99 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[434\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame7_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit20 net62 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[207\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem.Inst_Frame8_bit31 net74 net100 VGND VGND VPWR VPWR Inst_LUT4AB_ConfigMem.ConfigBits\[597\]
+ Inst_LUT4AB_ConfigMem.Inst_Frame8_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
+ Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.A1 VGND VGND
+ VPWR VPWR Inst_LUT4AB_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux21_inst.AIN\[1\]
+ sky130_fd_sc_hd__clkbuf_1
.ends

