VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO summer_school_top_wrapper
  CLASS BLOCK ;
  FOREIGN summer_school_top_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 85.720 2920.000 86.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2216.370 3516.000 2216.650 3520.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1892.070 3516.000 1892.350 3520.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1567.770 3516.000 1568.050 3520.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1243.470 3516.000 1243.750 3520.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 919.170 3516.000 919.450 3520.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 594.870 3516.000 595.150 3520.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 270.570 3516.000 270.850 3520.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3459.880 4.000 3460.480 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3211.000 4.000 3211.600 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2962.120 4.000 2962.720 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 522.280 2920.000 522.880 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2713.240 4.000 2713.840 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2464.360 4.000 2464.960 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2215.480 4.000 2216.080 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1966.600 4.000 1967.200 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1717.720 4.000 1718.320 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.840 4.000 1469.440 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1219.960 4.000 1220.560 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 958.840 2920.000 959.440 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_in[30]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1395.400 2920.000 1396.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1831.960 2920.000 1832.560 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2268.520 2920.000 2269.120 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2705.080 2920.000 2705.680 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3141.640 2920.000 3142.240 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 2864.970 3516.000 2865.250 3520.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2540.670 3516.000 2540.950 3520.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 376.760 2920.000 377.360 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2000.170 3516.000 2000.450 3520.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1675.870 3516.000 1676.150 3520.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1351.570 3516.000 1351.850 3520.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1027.270 3516.000 1027.550 3520.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 702.970 3516.000 703.250 3520.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 378.670 3516.000 378.950 3520.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 54.370 3516.000 54.650 3520.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3293.960 4.000 3294.560 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3045.080 4.000 3045.680 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2796.200 4.000 2796.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 813.320 2920.000 813.920 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2547.320 4.000 2547.920 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2298.440 4.000 2299.040 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2049.560 4.000 2050.160 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1800.680 4.000 1801.280 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1551.800 4.000 1552.400 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.920 4.000 1303.520 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1249.880 2920.000 1250.480 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END io_oeb[30]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1686.440 2920.000 1687.040 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2123.000 2920.000 2123.600 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2559.560 2920.000 2560.160 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2996.120 2920.000 2996.720 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3432.680 2920.000 3433.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2648.770 3516.000 2649.050 3520.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2324.470 3516.000 2324.750 3520.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 231.240 2920.000 231.840 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2108.270 3516.000 2108.550 3520.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1783.970 3516.000 1784.250 3520.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1459.670 3516.000 1459.950 3520.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1135.370 3516.000 1135.650 3520.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 811.070 3516.000 811.350 3520.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 486.770 3516.000 487.050 3520.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.470 3516.000 162.750 3520.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3376.920 4.000 3377.520 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3128.040 4.000 3128.640 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2879.160 4.000 2879.760 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 667.800 2920.000 668.400 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2630.280 4.000 2630.880 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2381.400 4.000 2382.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2132.520 4.000 2133.120 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1883.640 4.000 1884.240 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1634.760 4.000 1635.360 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.880 4.000 1386.480 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1104.360 2920.000 1104.960 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END io_out[30]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1540.920 2920.000 1541.520 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1977.480 2920.000 1978.080 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2414.040 2920.000 2414.640 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2850.600 2920.000 2851.200 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3287.160 2920.000 3287.760 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2756.870 3516.000 2757.150 3520.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2432.570 3516.000 2432.850 3520.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.710 0.000 2413.990 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.650 0.000 2431.930 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2449.590 0.000 2449.870 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 2467.530 0.000 2467.810 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2485.470 0.000 2485.750 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2503.410 0.000 2503.690 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2521.350 0.000 2521.630 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2539.290 0.000 2539.570 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2557.230 0.000 2557.510 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.170 0.000 2575.450 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.110 0.000 799.390 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.110 0.000 2593.390 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2611.050 0.000 2611.330 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2628.990 0.000 2629.270 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2646.930 0.000 2647.210 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2664.870 0.000 2665.150 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.810 0.000 2683.090 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2700.750 0.000 2701.030 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2718.690 0.000 2718.970 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.630 0.000 2736.910 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2754.570 0.000 2754.850 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2772.510 0.000 2772.790 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2790.450 0.000 2790.730 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2808.390 0.000 2808.670 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2826.330 0.000 2826.610 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2844.270 0.000 2844.550 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2862.210 0.000 2862.490 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2880.150 0.000 2880.430 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.090 0.000 2898.370 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.930 0.000 853.210 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 0.000 907.030 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 0.000 978.790 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 0.000 996.730 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.210 0.000 1068.490 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 0.000 1086.430 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.030 0.000 1122.310 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 0.000 1158.190 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 0.000 1176.130 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 0.000 1194.070 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 0.000 1212.010 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.670 0.000 1229.950 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 0.000 1247.890 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.490 0.000 1283.770 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 0.000 1301.710 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1337.310 0.000 1337.590 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1355.250 0.000 1355.530 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1409.070 0.000 1409.350 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1427.010 0.000 1427.290 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1444.950 0.000 1445.230 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1462.890 0.000 1463.170 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1480.830 0.000 1481.110 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1498.770 0.000 1499.050 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 0.000 691.750 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1516.710 0.000 1516.990 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1534.650 0.000 1534.930 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1552.590 0.000 1552.870 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1570.530 0.000 1570.810 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1588.470 0.000 1588.750 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1606.410 0.000 1606.690 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1624.350 0.000 1624.630 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1660.230 0.000 1660.510 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1678.170 0.000 1678.450 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1696.110 0.000 1696.390 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1714.050 0.000 1714.330 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1731.990 0.000 1732.270 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1749.930 0.000 1750.210 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1767.870 0.000 1768.150 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1785.810 0.000 1786.090 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1803.750 0.000 1804.030 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1821.690 0.000 1821.970 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1839.630 0.000 1839.910 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1857.570 0.000 1857.850 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1875.510 0.000 1875.790 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1893.450 0.000 1893.730 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1911.390 0.000 1911.670 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1929.330 0.000 1929.610 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1947.270 0.000 1947.550 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1965.210 0.000 1965.490 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1983.150 0.000 1983.430 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2001.090 0.000 2001.370 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2036.970 0.000 2037.250 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2054.910 0.000 2055.190 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2072.850 0.000 2073.130 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2090.790 0.000 2091.070 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2108.730 0.000 2109.010 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.670 0.000 2126.950 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.610 0.000 2144.890 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.550 0.000 2162.830 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.490 0.000 2180.770 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.430 0.000 2198.710 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2216.370 0.000 2216.650 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2234.310 0.000 2234.590 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2252.250 0.000 2252.530 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 0.000 2270.470 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2288.130 0.000 2288.410 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.070 0.000 2306.350 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.010 0.000 2324.290 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.950 0.000 2342.230 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2359.890 0.000 2360.170 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.830 0.000 2378.110 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.770 0.000 2396.050 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.690 0.000 2419.970 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.630 0.000 2437.910 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.570 0.000 2455.850 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.510 0.000 2473.790 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.450 0.000 2491.730 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2509.390 0.000 2509.670 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.330 0.000 2527.610 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2545.270 0.000 2545.550 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.210 0.000 2563.490 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2581.150 0.000 2581.430 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.090 0.000 2599.370 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2617.030 0.000 2617.310 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2634.970 0.000 2635.250 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2652.910 0.000 2653.190 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2670.850 0.000 2671.130 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2688.790 0.000 2689.070 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2706.730 0.000 2707.010 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2724.670 0.000 2724.950 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2742.610 0.000 2742.890 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2760.550 0.000 2760.830 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 823.030 0.000 823.310 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2778.490 0.000 2778.770 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2796.430 0.000 2796.710 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2814.370 0.000 2814.650 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2832.310 0.000 2832.590 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2850.250 0.000 2850.530 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2868.190 0.000 2868.470 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2886.130 0.000 2886.410 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2904.070 0.000 2904.350 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 840.970 0.000 841.250 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 912.730 0.000 913.010 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.670 0.000 930.950 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 0.000 966.830 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.490 0.000 984.770 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.370 0.000 1020.650 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 0.000 1038.590 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.190 0.000 1074.470 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 0.000 1110.350 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 0.000 1146.230 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 661.570 0.000 661.850 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 0.000 1164.170 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 0.000 1182.110 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.770 0.000 1200.050 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1217.710 0.000 1217.990 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.650 0.000 1235.930 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1253.590 0.000 1253.870 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1289.470 0.000 1289.750 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1307.410 0.000 1307.690 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.290 0.000 1343.570 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1361.230 0.000 1361.510 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.050 0.000 1415.330 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 0.000 1433.270 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.930 0.000 1451.210 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.870 0.000 1469.150 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.810 0.000 1487.090 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.750 0.000 1505.030 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.690 0.000 1522.970 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.630 0.000 1540.910 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.510 0.000 1576.790 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.450 0.000 1594.730 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.390 0.000 1612.670 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.330 0.000 1630.610 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.270 0.000 1648.550 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 0.000 1666.490 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 0.000 1684.430 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.090 0.000 1702.370 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.030 0.000 1720.310 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.970 0.000 1738.250 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.910 0.000 1756.190 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.850 0.000 1774.130 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.790 0.000 1792.070 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.730 0.000 1810.010 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.670 0.000 1827.950 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.610 0.000 1845.890 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.550 0.000 1863.830 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.490 0.000 1881.770 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.430 0.000 1899.710 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.370 0.000 1917.650 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.310 0.000 1935.590 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.250 0.000 1953.530 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.190 0.000 1971.470 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.130 0.000 1989.410 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.070 0.000 2007.350 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.010 0.000 2025.290 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.950 0.000 2043.230 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.890 0.000 2061.170 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.830 0.000 2079.110 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.770 0.000 2097.050 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2114.710 0.000 2114.990 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2132.650 0.000 2132.930 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2150.590 0.000 2150.870 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.530 0.000 2168.810 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.470 0.000 2186.750 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.410 0.000 2204.690 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2222.350 0.000 2222.630 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 769.210 0.000 769.490 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.290 0.000 2240.570 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2258.230 0.000 2258.510 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.170 0.000 2276.450 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2294.110 0.000 2294.390 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 0.000 2312.330 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.990 0.000 2330.270 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.930 0.000 2348.210 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2365.870 0.000 2366.150 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2383.810 0.000 2384.090 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2401.750 0.000 2402.030 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.670 0.000 2425.950 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.610 0.000 2443.890 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.550 0.000 2461.830 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.490 0.000 2479.770 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2497.430 0.000 2497.710 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2515.370 0.000 2515.650 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.310 0.000 2533.590 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2551.250 0.000 2551.530 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2569.190 0.000 2569.470 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2587.130 0.000 2587.410 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2605.070 0.000 2605.350 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2623.010 0.000 2623.290 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2640.950 0.000 2641.230 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2658.890 0.000 2659.170 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.830 0.000 2677.110 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2694.770 0.000 2695.050 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2712.710 0.000 2712.990 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2730.650 0.000 2730.930 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.590 0.000 2748.870 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2766.530 0.000 2766.810 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 0.000 829.290 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2784.470 0.000 2784.750 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2802.410 0.000 2802.690 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2820.350 0.000 2820.630 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2838.290 0.000 2838.570 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2856.230 0.000 2856.510 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2874.170 0.000 2874.450 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.110 0.000 2892.390 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.050 0.000 2910.330 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 0.000 865.170 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.770 0.000 901.050 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 0.000 918.990 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.650 0.000 936.930 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.590 0.000 954.870 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.470 0.000 990.750 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 0.000 1062.510 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.170 0.000 1080.450 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.050 0.000 1116.330 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.990 0.000 1134.270 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 0.000 1206.030 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1223.690 0.000 1223.970 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.630 0.000 1241.910 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.570 0.000 1259.850 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.510 0.000 1277.790 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.450 0.000 1295.730 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.390 0.000 1313.670 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.330 0.000 1331.610 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 0.000 1349.550 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 0.000 1367.490 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.030 0.000 1421.310 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.970 0.000 1439.250 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 0.000 1475.130 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 0.000 1493.070 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.730 0.000 1511.010 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 0.000 703.710 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.670 0.000 1528.950 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.610 0.000 1546.890 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.550 0.000 1564.830 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.490 0.000 1582.770 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1618.370 0.000 1618.650 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.310 0.000 1636.590 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.250 0.000 1654.530 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 0.000 1690.410 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.070 0.000 1708.350 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.950 0.000 1744.230 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.890 0.000 1762.170 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 0.000 1780.110 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1797.770 0.000 1798.050 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.710 0.000 1815.990 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.650 0.000 1833.930 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 0.000 1851.870 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.530 0.000 1869.810 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 0.000 1887.750 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.410 0.000 1905.690 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.350 0.000 1923.630 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.290 0.000 1941.570 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.170 0.000 1977.450 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.110 0.000 1995.390 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.050 0.000 2013.330 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.990 0.000 2031.270 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.930 0.000 2049.210 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.870 0.000 2067.150 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.810 0.000 2085.090 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 0.000 2103.030 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2120.690 0.000 2120.970 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.630 0.000 2138.910 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.570 0.000 2156.850 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.510 0.000 2174.790 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2192.450 0.000 2192.730 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.390 0.000 2210.670 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.330 0.000 2228.610 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 0.000 775.470 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.270 0.000 2246.550 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.210 0.000 2264.490 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.150 0.000 2282.430 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2300.090 0.000 2300.370 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.030 0.000 2318.310 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2335.970 0.000 2336.250 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 0.000 2354.190 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2371.850 0.000 2372.130 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.790 0.000 2390.070 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2407.730 0.000 2408.010 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.130 0.000 793.410 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2916.030 0.000 2916.310 4.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 3525.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 -6.220 2931.200 -3.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 3522.800 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.100 -6.220 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.020 -11.020 7.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.020 -11.020 57.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.020 2619.480 57.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.020 -11.020 107.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.020 2619.480 107.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.020 -11.020 157.020 404.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.020 1938.440 157.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.020 2619.480 157.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.020 -11.020 207.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.020 2619.480 207.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 -11.020 257.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 1940.065 257.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 2620.100 257.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.020 -11.020 307.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.020 1995.920 307.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.020 2619.480 307.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.020 -11.020 357.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.020 1979.185 357.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.020 2620.100 357.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 -11.020 407.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 1940.065 407.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 2619.480 407.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.020 -11.020 457.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.020 2619.480 457.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.020 -11.020 507.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.020 1940.065 507.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.020 2619.480 507.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.020 -11.020 557.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.020 1995.920 557.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.020 -11.020 607.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.020 1979.185 607.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.020 -11.020 657.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.020 1940.065 657.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.020 -11.020 707.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 754.020 -11.020 757.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 754.020 1940.065 757.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 804.020 -11.020 807.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 804.020 1995.920 807.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.020 -11.020 857.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.020 1979.185 857.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.020 -11.020 907.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.020 1940.065 907.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.020 -11.020 957.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.020 1940.065 957.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1004.020 -11.020 1007.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1004.020 1995.920 1007.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.020 -11.020 1057.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.020 1979.185 1057.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.020 -11.020 1107.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.020 1979.185 1107.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1154.020 -11.020 1157.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1154.020 1940.065 1157.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1204.020 -11.020 1207.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1204.020 1940.065 1207.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.020 -11.020 1257.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.020 1940.065 1257.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.020 -11.020 1307.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.020 1995.920 1307.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1354.020 -11.020 1357.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1354.020 1995.920 1357.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1404.020 -11.020 1407.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1404.020 1940.065 1407.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.020 -11.020 1457.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.020 1940.065 1457.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.020 -11.020 1507.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.020 1940.065 1507.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.020 -11.020 1557.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.020 1979.185 1557.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.020 -11.020 1607.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.020 1940.065 1607.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.020 -11.020 1657.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.020 1995.920 1657.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.020 -11.020 1707.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.020 1995.920 1707.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.020 -11.020 1757.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.020 1979.185 1757.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.020 -11.020 1807.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.020 1979.185 1807.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.020 -11.020 1857.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.020 1940.065 1857.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.020 -11.020 1907.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.020 1940.065 1907.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.020 -11.020 1957.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.020 1940.065 1957.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.020 -11.020 2007.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.020 1940.065 2007.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.020 -11.020 2057.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.020 1979.185 2057.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.020 -11.020 2107.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.020 1940.065 2107.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.020 -11.020 2157.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.020 1940.065 2157.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2204.020 -11.020 2207.020 339.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2204.020 1995.480 2207.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.020 -11.020 2257.020 405.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.020 1994.385 2257.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.020 -11.020 2307.020 339.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.020 1995.480 2307.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.020 -11.020 2357.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 -11.020 2407.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 859.380 2407.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 1379.480 2407.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 1899.480 2407.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 -11.020 2457.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 859.380 2457.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 1379.480 2457.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 1899.480 2457.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 -11.020 2507.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 859.380 2507.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 1379.480 2507.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 1899.480 2507.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 -11.020 2557.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 860.100 2557.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 1380.100 2557.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 1900.100 2557.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 -11.020 2607.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 860.100 2607.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 1380.100 2607.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 1900.100 2607.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 -11.020 2657.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 860.100 2657.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 1380.100 2657.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 1900.100 2657.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 -11.020 2707.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 860.100 2707.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 1380.100 2707.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 1900.100 2707.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 -11.020 2757.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 859.380 2757.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 1379.480 2757.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 1899.480 2757.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 -11.020 2807.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 859.380 2807.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 1379.480 2807.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 1899.480 2807.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 -11.020 2857.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 859.380 2857.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 1379.480 2857.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 1899.480 2857.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2904.020 -11.020 2907.020 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 9.380 2936.000 12.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 59.380 2936.000 62.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 109.380 2936.000 112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 159.380 2936.000 162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 209.380 2936.000 212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 259.380 2936.000 262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 309.380 2936.000 312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 359.380 2936.000 362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 409.380 2936.000 412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 459.380 2936.000 462.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 509.380 2936.000 512.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 559.380 2936.000 562.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 609.380 2936.000 612.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 659.380 2936.000 662.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 709.380 2936.000 712.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 759.380 2936.000 762.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 809.380 2936.000 812.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 859.380 2936.000 862.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 909.380 2936.000 912.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 959.380 2936.000 962.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1009.380 2936.000 1012.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1059.380 2936.000 1062.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1109.380 2936.000 1112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1159.380 2936.000 1162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1209.380 2936.000 1212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1259.380 2936.000 1262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1309.380 2936.000 1312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1359.380 2936.000 1362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1409.380 2936.000 1412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1459.380 2936.000 1462.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1509.380 2936.000 1512.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1559.380 2936.000 1562.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1609.380 2936.000 1612.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1659.380 2936.000 1662.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1709.380 2936.000 1712.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1759.380 2936.000 1762.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1809.380 2936.000 1812.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1859.380 2936.000 1862.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1909.380 2936.000 1912.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1959.380 2936.000 1962.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2009.380 2936.000 2012.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2059.380 2936.000 2062.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2109.380 2936.000 2112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2159.380 2936.000 2162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2209.380 2936.000 2212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2259.380 2936.000 2262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2309.380 2936.000 2312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2359.380 2936.000 2362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2409.380 2936.000 2412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2459.380 2936.000 2462.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2509.380 2936.000 2512.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2559.380 2936.000 2562.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2609.380 2936.000 2612.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2659.380 2936.000 2662.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2709.380 2936.000 2712.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2759.380 2936.000 2762.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2809.380 2936.000 2812.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2859.380 2936.000 2862.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2909.380 2936.000 2912.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2959.380 2936.000 2962.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3009.380 2936.000 3012.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3059.380 2936.000 3062.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3109.380 2936.000 3112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3159.380 2936.000 3162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3209.380 2936.000 3212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3259.380 2936.000 3262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3309.380 2936.000 3312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3359.380 2936.000 3362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3409.380 2936.000 3412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3459.380 2936.000 3462.380 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 -11.020 2936.000 -7.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3527.600 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2932.900 -11.020 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.720 -11.020 11.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.720 -11.020 61.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.720 2619.480 61.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.720 -11.020 111.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.720 2619.480 111.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 -11.020 161.720 408.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 1931.225 161.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 2619.480 161.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 -11.020 211.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 1940.065 211.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 2620.100 211.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.720 -11.020 261.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.720 1940.065 261.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.720 2620.100 261.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.720 -11.020 311.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.720 1979.185 311.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.720 2620.100 311.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.720 -11.020 361.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.720 1995.920 361.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.720 2620.100 361.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.720 -11.020 411.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.720 1940.065 411.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.720 2619.480 411.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.720 -11.020 461.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.720 1940.065 461.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.720 2619.480 461.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.720 -11.020 511.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.720 1940.065 511.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.720 2619.480 511.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.720 -11.020 561.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.720 1979.185 561.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.720 -11.020 611.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.720 1995.920 611.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.720 -11.020 661.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.720 1940.065 661.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.720 -11.020 711.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.720 1940.065 711.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.720 -11.020 761.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.720 1940.065 761.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.720 -11.020 811.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.720 1979.185 811.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 -11.020 861.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 1995.920 861.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 -11.020 911.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 1940.065 911.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 958.720 -11.020 961.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 958.720 1940.065 961.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.720 -11.020 1011.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.720 1940.065 1011.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.720 -11.020 1061.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.720 1995.920 1061.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.720 -11.020 1111.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.720 1979.185 1111.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.720 -11.020 1161.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.720 1940.065 1161.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.720 -11.020 1211.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.720 1940.065 1211.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.720 -11.020 1261.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.720 1940.065 1261.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.720 -11.020 1311.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.720 1979.185 1311.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.720 -11.020 1361.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.720 1995.920 1361.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.720 -11.020 1411.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.720 1995.920 1411.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.720 -11.020 1461.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.720 1940.065 1461.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.720 -11.020 1511.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.720 1940.065 1511.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.720 -11.020 1561.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.720 1979.185 1561.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.720 -11.020 1611.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.720 1940.065 1611.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.720 -11.020 1661.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.720 1940.065 1661.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1708.720 -11.020 1711.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1708.720 1940.065 1711.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.720 -11.020 1761.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.720 1995.920 1761.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.720 -11.020 1811.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.720 1979.185 1811.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.720 -11.020 1861.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.720 1940.065 1861.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1908.720 -11.020 1911.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.720 -11.020 1961.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.720 1995.920 1961.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.720 -11.020 2011.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.720 1979.185 2011.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.720 -11.020 2061.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.720 1979.185 2061.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.720 -11.020 2111.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.720 1940.065 2111.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.720 -11.020 2161.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.720 1940.065 2161.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.720 -11.020 2211.720 405.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.720 1935.305 2211.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.720 -11.020 2261.720 405.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.720 1994.385 2261.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.720 -11.020 2311.720 339.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.720 1995.480 2311.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.720 -11.020 2361.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 -11.020 2411.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 859.480 2411.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 1379.480 2411.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 1899.480 2411.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 -11.020 2461.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 859.480 2461.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 1379.480 2461.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 1899.480 2461.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 -11.020 2511.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 859.480 2511.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 1379.480 2511.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 1899.480 2511.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 -11.020 2561.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 860.100 2561.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 1380.100 2561.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 1900.100 2561.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 -11.020 2611.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 860.100 2611.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 1380.100 2611.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 1900.100 2611.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 -11.020 2661.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 860.100 2661.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 1380.100 2661.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 1900.100 2661.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 -11.020 2711.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 860.100 2711.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 1380.100 2711.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 1900.100 2711.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 -11.020 2761.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 859.480 2761.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 1379.480 2761.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 1899.480 2761.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 -11.020 2811.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 859.480 2811.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 1379.480 2811.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 1899.480 2811.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 -11.020 2861.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 859.480 2861.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 1379.480 2861.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 1899.480 2861.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2908.720 -11.020 2911.720 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 14.080 2936.000 17.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 64.080 2936.000 67.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 114.080 2936.000 117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 164.080 2936.000 167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 214.080 2936.000 217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 264.080 2936.000 267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 314.080 2936.000 317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 364.080 2936.000 367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 414.080 2936.000 417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 464.080 2936.000 467.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 514.080 2936.000 517.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 564.080 2936.000 567.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 614.080 2936.000 617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 664.080 2936.000 667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 714.080 2936.000 717.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 764.080 2936.000 767.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 814.080 2936.000 817.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 864.080 2936.000 867.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 914.080 2936.000 917.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 964.080 2936.000 967.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1014.080 2936.000 1017.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1064.080 2936.000 1067.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1114.080 2936.000 1117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1164.080 2936.000 1167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1214.080 2936.000 1217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1264.080 2936.000 1267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1314.080 2936.000 1317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1364.080 2936.000 1367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1414.080 2936.000 1417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1464.080 2936.000 1467.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1514.080 2936.000 1517.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1564.080 2936.000 1567.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1614.080 2936.000 1617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1664.080 2936.000 1667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1714.080 2936.000 1717.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1764.080 2936.000 1767.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1814.080 2936.000 1817.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1864.080 2936.000 1867.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1914.080 2936.000 1917.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1964.080 2936.000 1967.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2014.080 2936.000 2017.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2064.080 2936.000 2067.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2114.080 2936.000 2117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2164.080 2936.000 2167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2214.080 2936.000 2217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2264.080 2936.000 2267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2314.080 2936.000 2317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2364.080 2936.000 2367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2414.080 2936.000 2417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2464.080 2936.000 2467.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2514.080 2936.000 2517.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2564.080 2936.000 2567.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2614.080 2936.000 2617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2664.080 2936.000 2667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2714.080 2936.000 2717.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2764.080 2936.000 2767.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2814.080 2936.000 2817.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2864.080 2936.000 2867.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2914.080 2936.000 2917.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2964.080 2936.000 2967.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3014.080 2936.000 3017.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3064.080 2936.000 3067.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3114.080 2936.000 3117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3164.080 2936.000 3167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3214.080 2936.000 3217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3264.080 2936.000 3267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3314.080 2936.000 3317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3364.080 2936.000 3367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3414.080 2936.000 3417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3464.080 2936.000 3467.080 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 422.370 0.000 422.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 547.950 0.000 548.230 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 601.770 0.000 602.050 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 356.590 0.000 356.870 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 410.410 0.000 410.690 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 482.170 0.000 482.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 0.000 560.190 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sta_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END wbs_sta_o
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 2.370 6.500 2917.250 3509.040 ;
      LAYER met2 ;
        RECT 2.400 3515.720 54.090 3516.690 ;
        RECT 54.930 3515.720 162.190 3516.690 ;
        RECT 163.030 3515.720 270.290 3516.690 ;
        RECT 271.130 3515.720 378.390 3516.690 ;
        RECT 379.230 3515.720 486.490 3516.690 ;
        RECT 487.330 3515.720 594.590 3516.690 ;
        RECT 595.430 3515.720 702.690 3516.690 ;
        RECT 703.530 3515.720 810.790 3516.690 ;
        RECT 811.630 3515.720 918.890 3516.690 ;
        RECT 919.730 3515.720 1026.990 3516.690 ;
        RECT 1027.830 3515.720 1135.090 3516.690 ;
        RECT 1135.930 3515.720 1243.190 3516.690 ;
        RECT 1244.030 3515.720 1351.290 3516.690 ;
        RECT 1352.130 3515.720 1459.390 3516.690 ;
        RECT 1460.230 3515.720 1567.490 3516.690 ;
        RECT 1568.330 3515.720 1675.590 3516.690 ;
        RECT 1676.430 3515.720 1783.690 3516.690 ;
        RECT 1784.530 3515.720 1891.790 3516.690 ;
        RECT 1892.630 3515.720 1999.890 3516.690 ;
        RECT 2000.730 3515.720 2107.990 3516.690 ;
        RECT 2108.830 3515.720 2216.090 3516.690 ;
        RECT 2216.930 3515.720 2324.190 3516.690 ;
        RECT 2325.030 3515.720 2432.290 3516.690 ;
        RECT 2433.130 3515.720 2540.390 3516.690 ;
        RECT 2541.230 3515.720 2648.490 3516.690 ;
        RECT 2649.330 3515.720 2756.590 3516.690 ;
        RECT 2757.430 3515.720 2864.690 3516.690 ;
        RECT 2865.530 3515.720 2917.220 3516.690 ;
        RECT 2.400 4.280 2917.220 3515.720 ;
        RECT 2.400 3.670 3.490 4.280 ;
        RECT 4.330 3.670 9.470 4.280 ;
        RECT 10.310 3.670 15.450 4.280 ;
        RECT 16.290 3.670 21.430 4.280 ;
        RECT 22.270 3.670 27.410 4.280 ;
        RECT 28.250 3.670 33.390 4.280 ;
        RECT 34.230 3.670 39.370 4.280 ;
        RECT 40.210 3.670 45.350 4.280 ;
        RECT 46.190 3.670 51.330 4.280 ;
        RECT 52.170 3.670 57.310 4.280 ;
        RECT 58.150 3.670 63.290 4.280 ;
        RECT 64.130 3.670 69.270 4.280 ;
        RECT 70.110 3.670 75.250 4.280 ;
        RECT 76.090 3.670 81.230 4.280 ;
        RECT 82.070 3.670 87.210 4.280 ;
        RECT 88.050 3.670 93.190 4.280 ;
        RECT 94.030 3.670 99.170 4.280 ;
        RECT 100.010 3.670 105.150 4.280 ;
        RECT 105.990 3.670 111.130 4.280 ;
        RECT 111.970 3.670 117.110 4.280 ;
        RECT 117.950 3.670 123.090 4.280 ;
        RECT 123.930 3.670 129.070 4.280 ;
        RECT 129.910 3.670 135.050 4.280 ;
        RECT 135.890 3.670 141.030 4.280 ;
        RECT 141.870 3.670 147.010 4.280 ;
        RECT 147.850 3.670 152.990 4.280 ;
        RECT 153.830 3.670 158.970 4.280 ;
        RECT 159.810 3.670 164.950 4.280 ;
        RECT 165.790 3.670 170.930 4.280 ;
        RECT 171.770 3.670 176.910 4.280 ;
        RECT 177.750 3.670 182.890 4.280 ;
        RECT 183.730 3.670 188.870 4.280 ;
        RECT 189.710 3.670 194.850 4.280 ;
        RECT 195.690 3.670 200.830 4.280 ;
        RECT 201.670 3.670 206.810 4.280 ;
        RECT 207.650 3.670 212.790 4.280 ;
        RECT 213.630 3.670 218.770 4.280 ;
        RECT 219.610 3.670 224.750 4.280 ;
        RECT 225.590 3.670 230.730 4.280 ;
        RECT 231.570 3.670 236.710 4.280 ;
        RECT 237.550 3.670 242.690 4.280 ;
        RECT 243.530 3.670 248.670 4.280 ;
        RECT 249.510 3.670 254.650 4.280 ;
        RECT 255.490 3.670 260.630 4.280 ;
        RECT 261.470 3.670 266.610 4.280 ;
        RECT 267.450 3.670 272.590 4.280 ;
        RECT 273.430 3.670 278.570 4.280 ;
        RECT 279.410 3.670 284.550 4.280 ;
        RECT 285.390 3.670 290.530 4.280 ;
        RECT 291.370 3.670 296.510 4.280 ;
        RECT 297.350 3.670 302.490 4.280 ;
        RECT 303.330 3.670 308.470 4.280 ;
        RECT 309.310 3.670 314.450 4.280 ;
        RECT 315.290 3.670 320.430 4.280 ;
        RECT 321.270 3.670 326.410 4.280 ;
        RECT 327.250 3.670 332.390 4.280 ;
        RECT 333.230 3.670 338.370 4.280 ;
        RECT 339.210 3.670 344.350 4.280 ;
        RECT 345.190 3.670 350.330 4.280 ;
        RECT 351.170 3.670 356.310 4.280 ;
        RECT 357.150 3.670 362.290 4.280 ;
        RECT 363.130 3.670 368.270 4.280 ;
        RECT 369.110 3.670 374.250 4.280 ;
        RECT 375.090 3.670 380.230 4.280 ;
        RECT 381.070 3.670 386.210 4.280 ;
        RECT 387.050 3.670 392.190 4.280 ;
        RECT 393.030 3.670 398.170 4.280 ;
        RECT 399.010 3.670 404.150 4.280 ;
        RECT 404.990 3.670 410.130 4.280 ;
        RECT 410.970 3.670 416.110 4.280 ;
        RECT 416.950 3.670 422.090 4.280 ;
        RECT 422.930 3.670 428.070 4.280 ;
        RECT 428.910 3.670 434.050 4.280 ;
        RECT 434.890 3.670 440.030 4.280 ;
        RECT 440.870 3.670 446.010 4.280 ;
        RECT 446.850 3.670 451.990 4.280 ;
        RECT 452.830 3.670 457.970 4.280 ;
        RECT 458.810 3.670 463.950 4.280 ;
        RECT 464.790 3.670 469.930 4.280 ;
        RECT 470.770 3.670 475.910 4.280 ;
        RECT 476.750 3.670 481.890 4.280 ;
        RECT 482.730 3.670 487.870 4.280 ;
        RECT 488.710 3.670 493.850 4.280 ;
        RECT 494.690 3.670 499.830 4.280 ;
        RECT 500.670 3.670 505.810 4.280 ;
        RECT 506.650 3.670 511.790 4.280 ;
        RECT 512.630 3.670 517.770 4.280 ;
        RECT 518.610 3.670 523.750 4.280 ;
        RECT 524.590 3.670 529.730 4.280 ;
        RECT 530.570 3.670 535.710 4.280 ;
        RECT 536.550 3.670 541.690 4.280 ;
        RECT 542.530 3.670 547.670 4.280 ;
        RECT 548.510 3.670 553.650 4.280 ;
        RECT 554.490 3.670 559.630 4.280 ;
        RECT 560.470 3.670 565.610 4.280 ;
        RECT 566.450 3.670 571.590 4.280 ;
        RECT 572.430 3.670 577.570 4.280 ;
        RECT 578.410 3.670 583.550 4.280 ;
        RECT 584.390 3.670 589.530 4.280 ;
        RECT 590.370 3.670 595.510 4.280 ;
        RECT 596.350 3.670 601.490 4.280 ;
        RECT 602.330 3.670 607.470 4.280 ;
        RECT 608.310 3.670 613.450 4.280 ;
        RECT 614.290 3.670 619.430 4.280 ;
        RECT 620.270 3.670 625.410 4.280 ;
        RECT 626.250 3.670 631.390 4.280 ;
        RECT 632.230 3.670 637.370 4.280 ;
        RECT 638.210 3.670 643.350 4.280 ;
        RECT 644.190 3.670 649.330 4.280 ;
        RECT 650.170 3.670 655.310 4.280 ;
        RECT 656.150 3.670 661.290 4.280 ;
        RECT 662.130 3.670 667.270 4.280 ;
        RECT 668.110 3.670 673.250 4.280 ;
        RECT 674.090 3.670 679.230 4.280 ;
        RECT 680.070 3.670 685.210 4.280 ;
        RECT 686.050 3.670 691.190 4.280 ;
        RECT 692.030 3.670 697.170 4.280 ;
        RECT 698.010 3.670 703.150 4.280 ;
        RECT 703.990 3.670 709.130 4.280 ;
        RECT 709.970 3.670 715.110 4.280 ;
        RECT 715.950 3.670 721.090 4.280 ;
        RECT 721.930 3.670 727.070 4.280 ;
        RECT 727.910 3.670 733.050 4.280 ;
        RECT 733.890 3.670 739.030 4.280 ;
        RECT 739.870 3.670 745.010 4.280 ;
        RECT 745.850 3.670 750.990 4.280 ;
        RECT 751.830 3.670 756.970 4.280 ;
        RECT 757.810 3.670 762.950 4.280 ;
        RECT 763.790 3.670 768.930 4.280 ;
        RECT 769.770 3.670 774.910 4.280 ;
        RECT 775.750 3.670 780.890 4.280 ;
        RECT 781.730 3.670 786.870 4.280 ;
        RECT 787.710 3.670 792.850 4.280 ;
        RECT 793.690 3.670 798.830 4.280 ;
        RECT 799.670 3.670 804.810 4.280 ;
        RECT 805.650 3.670 810.790 4.280 ;
        RECT 811.630 3.670 816.770 4.280 ;
        RECT 817.610 3.670 822.750 4.280 ;
        RECT 823.590 3.670 828.730 4.280 ;
        RECT 829.570 3.670 834.710 4.280 ;
        RECT 835.550 3.670 840.690 4.280 ;
        RECT 841.530 3.670 846.670 4.280 ;
        RECT 847.510 3.670 852.650 4.280 ;
        RECT 853.490 3.670 858.630 4.280 ;
        RECT 859.470 3.670 864.610 4.280 ;
        RECT 865.450 3.670 870.590 4.280 ;
        RECT 871.430 3.670 876.570 4.280 ;
        RECT 877.410 3.670 882.550 4.280 ;
        RECT 883.390 3.670 888.530 4.280 ;
        RECT 889.370 3.670 894.510 4.280 ;
        RECT 895.350 3.670 900.490 4.280 ;
        RECT 901.330 3.670 906.470 4.280 ;
        RECT 907.310 3.670 912.450 4.280 ;
        RECT 913.290 3.670 918.430 4.280 ;
        RECT 919.270 3.670 924.410 4.280 ;
        RECT 925.250 3.670 930.390 4.280 ;
        RECT 931.230 3.670 936.370 4.280 ;
        RECT 937.210 3.670 942.350 4.280 ;
        RECT 943.190 3.670 948.330 4.280 ;
        RECT 949.170 3.670 954.310 4.280 ;
        RECT 955.150 3.670 960.290 4.280 ;
        RECT 961.130 3.670 966.270 4.280 ;
        RECT 967.110 3.670 972.250 4.280 ;
        RECT 973.090 3.670 978.230 4.280 ;
        RECT 979.070 3.670 984.210 4.280 ;
        RECT 985.050 3.670 990.190 4.280 ;
        RECT 991.030 3.670 996.170 4.280 ;
        RECT 997.010 3.670 1002.150 4.280 ;
        RECT 1002.990 3.670 1008.130 4.280 ;
        RECT 1008.970 3.670 1014.110 4.280 ;
        RECT 1014.950 3.670 1020.090 4.280 ;
        RECT 1020.930 3.670 1026.070 4.280 ;
        RECT 1026.910 3.670 1032.050 4.280 ;
        RECT 1032.890 3.670 1038.030 4.280 ;
        RECT 1038.870 3.670 1044.010 4.280 ;
        RECT 1044.850 3.670 1049.990 4.280 ;
        RECT 1050.830 3.670 1055.970 4.280 ;
        RECT 1056.810 3.670 1061.950 4.280 ;
        RECT 1062.790 3.670 1067.930 4.280 ;
        RECT 1068.770 3.670 1073.910 4.280 ;
        RECT 1074.750 3.670 1079.890 4.280 ;
        RECT 1080.730 3.670 1085.870 4.280 ;
        RECT 1086.710 3.670 1091.850 4.280 ;
        RECT 1092.690 3.670 1097.830 4.280 ;
        RECT 1098.670 3.670 1103.810 4.280 ;
        RECT 1104.650 3.670 1109.790 4.280 ;
        RECT 1110.630 3.670 1115.770 4.280 ;
        RECT 1116.610 3.670 1121.750 4.280 ;
        RECT 1122.590 3.670 1127.730 4.280 ;
        RECT 1128.570 3.670 1133.710 4.280 ;
        RECT 1134.550 3.670 1139.690 4.280 ;
        RECT 1140.530 3.670 1145.670 4.280 ;
        RECT 1146.510 3.670 1151.650 4.280 ;
        RECT 1152.490 3.670 1157.630 4.280 ;
        RECT 1158.470 3.670 1163.610 4.280 ;
        RECT 1164.450 3.670 1169.590 4.280 ;
        RECT 1170.430 3.670 1175.570 4.280 ;
        RECT 1176.410 3.670 1181.550 4.280 ;
        RECT 1182.390 3.670 1187.530 4.280 ;
        RECT 1188.370 3.670 1193.510 4.280 ;
        RECT 1194.350 3.670 1199.490 4.280 ;
        RECT 1200.330 3.670 1205.470 4.280 ;
        RECT 1206.310 3.670 1211.450 4.280 ;
        RECT 1212.290 3.670 1217.430 4.280 ;
        RECT 1218.270 3.670 1223.410 4.280 ;
        RECT 1224.250 3.670 1229.390 4.280 ;
        RECT 1230.230 3.670 1235.370 4.280 ;
        RECT 1236.210 3.670 1241.350 4.280 ;
        RECT 1242.190 3.670 1247.330 4.280 ;
        RECT 1248.170 3.670 1253.310 4.280 ;
        RECT 1254.150 3.670 1259.290 4.280 ;
        RECT 1260.130 3.670 1265.270 4.280 ;
        RECT 1266.110 3.670 1271.250 4.280 ;
        RECT 1272.090 3.670 1277.230 4.280 ;
        RECT 1278.070 3.670 1283.210 4.280 ;
        RECT 1284.050 3.670 1289.190 4.280 ;
        RECT 1290.030 3.670 1295.170 4.280 ;
        RECT 1296.010 3.670 1301.150 4.280 ;
        RECT 1301.990 3.670 1307.130 4.280 ;
        RECT 1307.970 3.670 1313.110 4.280 ;
        RECT 1313.950 3.670 1319.090 4.280 ;
        RECT 1319.930 3.670 1325.070 4.280 ;
        RECT 1325.910 3.670 1331.050 4.280 ;
        RECT 1331.890 3.670 1337.030 4.280 ;
        RECT 1337.870 3.670 1343.010 4.280 ;
        RECT 1343.850 3.670 1348.990 4.280 ;
        RECT 1349.830 3.670 1354.970 4.280 ;
        RECT 1355.810 3.670 1360.950 4.280 ;
        RECT 1361.790 3.670 1366.930 4.280 ;
        RECT 1367.770 3.670 1372.910 4.280 ;
        RECT 1373.750 3.670 1378.890 4.280 ;
        RECT 1379.730 3.670 1384.870 4.280 ;
        RECT 1385.710 3.670 1390.850 4.280 ;
        RECT 1391.690 3.670 1396.830 4.280 ;
        RECT 1397.670 3.670 1402.810 4.280 ;
        RECT 1403.650 3.670 1408.790 4.280 ;
        RECT 1409.630 3.670 1414.770 4.280 ;
        RECT 1415.610 3.670 1420.750 4.280 ;
        RECT 1421.590 3.670 1426.730 4.280 ;
        RECT 1427.570 3.670 1432.710 4.280 ;
        RECT 1433.550 3.670 1438.690 4.280 ;
        RECT 1439.530 3.670 1444.670 4.280 ;
        RECT 1445.510 3.670 1450.650 4.280 ;
        RECT 1451.490 3.670 1456.630 4.280 ;
        RECT 1457.470 3.670 1462.610 4.280 ;
        RECT 1463.450 3.670 1468.590 4.280 ;
        RECT 1469.430 3.670 1474.570 4.280 ;
        RECT 1475.410 3.670 1480.550 4.280 ;
        RECT 1481.390 3.670 1486.530 4.280 ;
        RECT 1487.370 3.670 1492.510 4.280 ;
        RECT 1493.350 3.670 1498.490 4.280 ;
        RECT 1499.330 3.670 1504.470 4.280 ;
        RECT 1505.310 3.670 1510.450 4.280 ;
        RECT 1511.290 3.670 1516.430 4.280 ;
        RECT 1517.270 3.670 1522.410 4.280 ;
        RECT 1523.250 3.670 1528.390 4.280 ;
        RECT 1529.230 3.670 1534.370 4.280 ;
        RECT 1535.210 3.670 1540.350 4.280 ;
        RECT 1541.190 3.670 1546.330 4.280 ;
        RECT 1547.170 3.670 1552.310 4.280 ;
        RECT 1553.150 3.670 1558.290 4.280 ;
        RECT 1559.130 3.670 1564.270 4.280 ;
        RECT 1565.110 3.670 1570.250 4.280 ;
        RECT 1571.090 3.670 1576.230 4.280 ;
        RECT 1577.070 3.670 1582.210 4.280 ;
        RECT 1583.050 3.670 1588.190 4.280 ;
        RECT 1589.030 3.670 1594.170 4.280 ;
        RECT 1595.010 3.670 1600.150 4.280 ;
        RECT 1600.990 3.670 1606.130 4.280 ;
        RECT 1606.970 3.670 1612.110 4.280 ;
        RECT 1612.950 3.670 1618.090 4.280 ;
        RECT 1618.930 3.670 1624.070 4.280 ;
        RECT 1624.910 3.670 1630.050 4.280 ;
        RECT 1630.890 3.670 1636.030 4.280 ;
        RECT 1636.870 3.670 1642.010 4.280 ;
        RECT 1642.850 3.670 1647.990 4.280 ;
        RECT 1648.830 3.670 1653.970 4.280 ;
        RECT 1654.810 3.670 1659.950 4.280 ;
        RECT 1660.790 3.670 1665.930 4.280 ;
        RECT 1666.770 3.670 1671.910 4.280 ;
        RECT 1672.750 3.670 1677.890 4.280 ;
        RECT 1678.730 3.670 1683.870 4.280 ;
        RECT 1684.710 3.670 1689.850 4.280 ;
        RECT 1690.690 3.670 1695.830 4.280 ;
        RECT 1696.670 3.670 1701.810 4.280 ;
        RECT 1702.650 3.670 1707.790 4.280 ;
        RECT 1708.630 3.670 1713.770 4.280 ;
        RECT 1714.610 3.670 1719.750 4.280 ;
        RECT 1720.590 3.670 1725.730 4.280 ;
        RECT 1726.570 3.670 1731.710 4.280 ;
        RECT 1732.550 3.670 1737.690 4.280 ;
        RECT 1738.530 3.670 1743.670 4.280 ;
        RECT 1744.510 3.670 1749.650 4.280 ;
        RECT 1750.490 3.670 1755.630 4.280 ;
        RECT 1756.470 3.670 1761.610 4.280 ;
        RECT 1762.450 3.670 1767.590 4.280 ;
        RECT 1768.430 3.670 1773.570 4.280 ;
        RECT 1774.410 3.670 1779.550 4.280 ;
        RECT 1780.390 3.670 1785.530 4.280 ;
        RECT 1786.370 3.670 1791.510 4.280 ;
        RECT 1792.350 3.670 1797.490 4.280 ;
        RECT 1798.330 3.670 1803.470 4.280 ;
        RECT 1804.310 3.670 1809.450 4.280 ;
        RECT 1810.290 3.670 1815.430 4.280 ;
        RECT 1816.270 3.670 1821.410 4.280 ;
        RECT 1822.250 3.670 1827.390 4.280 ;
        RECT 1828.230 3.670 1833.370 4.280 ;
        RECT 1834.210 3.670 1839.350 4.280 ;
        RECT 1840.190 3.670 1845.330 4.280 ;
        RECT 1846.170 3.670 1851.310 4.280 ;
        RECT 1852.150 3.670 1857.290 4.280 ;
        RECT 1858.130 3.670 1863.270 4.280 ;
        RECT 1864.110 3.670 1869.250 4.280 ;
        RECT 1870.090 3.670 1875.230 4.280 ;
        RECT 1876.070 3.670 1881.210 4.280 ;
        RECT 1882.050 3.670 1887.190 4.280 ;
        RECT 1888.030 3.670 1893.170 4.280 ;
        RECT 1894.010 3.670 1899.150 4.280 ;
        RECT 1899.990 3.670 1905.130 4.280 ;
        RECT 1905.970 3.670 1911.110 4.280 ;
        RECT 1911.950 3.670 1917.090 4.280 ;
        RECT 1917.930 3.670 1923.070 4.280 ;
        RECT 1923.910 3.670 1929.050 4.280 ;
        RECT 1929.890 3.670 1935.030 4.280 ;
        RECT 1935.870 3.670 1941.010 4.280 ;
        RECT 1941.850 3.670 1946.990 4.280 ;
        RECT 1947.830 3.670 1952.970 4.280 ;
        RECT 1953.810 3.670 1958.950 4.280 ;
        RECT 1959.790 3.670 1964.930 4.280 ;
        RECT 1965.770 3.670 1970.910 4.280 ;
        RECT 1971.750 3.670 1976.890 4.280 ;
        RECT 1977.730 3.670 1982.870 4.280 ;
        RECT 1983.710 3.670 1988.850 4.280 ;
        RECT 1989.690 3.670 1994.830 4.280 ;
        RECT 1995.670 3.670 2000.810 4.280 ;
        RECT 2001.650 3.670 2006.790 4.280 ;
        RECT 2007.630 3.670 2012.770 4.280 ;
        RECT 2013.610 3.670 2018.750 4.280 ;
        RECT 2019.590 3.670 2024.730 4.280 ;
        RECT 2025.570 3.670 2030.710 4.280 ;
        RECT 2031.550 3.670 2036.690 4.280 ;
        RECT 2037.530 3.670 2042.670 4.280 ;
        RECT 2043.510 3.670 2048.650 4.280 ;
        RECT 2049.490 3.670 2054.630 4.280 ;
        RECT 2055.470 3.670 2060.610 4.280 ;
        RECT 2061.450 3.670 2066.590 4.280 ;
        RECT 2067.430 3.670 2072.570 4.280 ;
        RECT 2073.410 3.670 2078.550 4.280 ;
        RECT 2079.390 3.670 2084.530 4.280 ;
        RECT 2085.370 3.670 2090.510 4.280 ;
        RECT 2091.350 3.670 2096.490 4.280 ;
        RECT 2097.330 3.670 2102.470 4.280 ;
        RECT 2103.310 3.670 2108.450 4.280 ;
        RECT 2109.290 3.670 2114.430 4.280 ;
        RECT 2115.270 3.670 2120.410 4.280 ;
        RECT 2121.250 3.670 2126.390 4.280 ;
        RECT 2127.230 3.670 2132.370 4.280 ;
        RECT 2133.210 3.670 2138.350 4.280 ;
        RECT 2139.190 3.670 2144.330 4.280 ;
        RECT 2145.170 3.670 2150.310 4.280 ;
        RECT 2151.150 3.670 2156.290 4.280 ;
        RECT 2157.130 3.670 2162.270 4.280 ;
        RECT 2163.110 3.670 2168.250 4.280 ;
        RECT 2169.090 3.670 2174.230 4.280 ;
        RECT 2175.070 3.670 2180.210 4.280 ;
        RECT 2181.050 3.670 2186.190 4.280 ;
        RECT 2187.030 3.670 2192.170 4.280 ;
        RECT 2193.010 3.670 2198.150 4.280 ;
        RECT 2198.990 3.670 2204.130 4.280 ;
        RECT 2204.970 3.670 2210.110 4.280 ;
        RECT 2210.950 3.670 2216.090 4.280 ;
        RECT 2216.930 3.670 2222.070 4.280 ;
        RECT 2222.910 3.670 2228.050 4.280 ;
        RECT 2228.890 3.670 2234.030 4.280 ;
        RECT 2234.870 3.670 2240.010 4.280 ;
        RECT 2240.850 3.670 2245.990 4.280 ;
        RECT 2246.830 3.670 2251.970 4.280 ;
        RECT 2252.810 3.670 2257.950 4.280 ;
        RECT 2258.790 3.670 2263.930 4.280 ;
        RECT 2264.770 3.670 2269.910 4.280 ;
        RECT 2270.750 3.670 2275.890 4.280 ;
        RECT 2276.730 3.670 2281.870 4.280 ;
        RECT 2282.710 3.670 2287.850 4.280 ;
        RECT 2288.690 3.670 2293.830 4.280 ;
        RECT 2294.670 3.670 2299.810 4.280 ;
        RECT 2300.650 3.670 2305.790 4.280 ;
        RECT 2306.630 3.670 2311.770 4.280 ;
        RECT 2312.610 3.670 2317.750 4.280 ;
        RECT 2318.590 3.670 2323.730 4.280 ;
        RECT 2324.570 3.670 2329.710 4.280 ;
        RECT 2330.550 3.670 2335.690 4.280 ;
        RECT 2336.530 3.670 2341.670 4.280 ;
        RECT 2342.510 3.670 2347.650 4.280 ;
        RECT 2348.490 3.670 2353.630 4.280 ;
        RECT 2354.470 3.670 2359.610 4.280 ;
        RECT 2360.450 3.670 2365.590 4.280 ;
        RECT 2366.430 3.670 2371.570 4.280 ;
        RECT 2372.410 3.670 2377.550 4.280 ;
        RECT 2378.390 3.670 2383.530 4.280 ;
        RECT 2384.370 3.670 2389.510 4.280 ;
        RECT 2390.350 3.670 2395.490 4.280 ;
        RECT 2396.330 3.670 2401.470 4.280 ;
        RECT 2402.310 3.670 2407.450 4.280 ;
        RECT 2408.290 3.670 2413.430 4.280 ;
        RECT 2414.270 3.670 2419.410 4.280 ;
        RECT 2420.250 3.670 2425.390 4.280 ;
        RECT 2426.230 3.670 2431.370 4.280 ;
        RECT 2432.210 3.670 2437.350 4.280 ;
        RECT 2438.190 3.670 2443.330 4.280 ;
        RECT 2444.170 3.670 2449.310 4.280 ;
        RECT 2450.150 3.670 2455.290 4.280 ;
        RECT 2456.130 3.670 2461.270 4.280 ;
        RECT 2462.110 3.670 2467.250 4.280 ;
        RECT 2468.090 3.670 2473.230 4.280 ;
        RECT 2474.070 3.670 2479.210 4.280 ;
        RECT 2480.050 3.670 2485.190 4.280 ;
        RECT 2486.030 3.670 2491.170 4.280 ;
        RECT 2492.010 3.670 2497.150 4.280 ;
        RECT 2497.990 3.670 2503.130 4.280 ;
        RECT 2503.970 3.670 2509.110 4.280 ;
        RECT 2509.950 3.670 2515.090 4.280 ;
        RECT 2515.930 3.670 2521.070 4.280 ;
        RECT 2521.910 3.670 2527.050 4.280 ;
        RECT 2527.890 3.670 2533.030 4.280 ;
        RECT 2533.870 3.670 2539.010 4.280 ;
        RECT 2539.850 3.670 2544.990 4.280 ;
        RECT 2545.830 3.670 2550.970 4.280 ;
        RECT 2551.810 3.670 2556.950 4.280 ;
        RECT 2557.790 3.670 2562.930 4.280 ;
        RECT 2563.770 3.670 2568.910 4.280 ;
        RECT 2569.750 3.670 2574.890 4.280 ;
        RECT 2575.730 3.670 2580.870 4.280 ;
        RECT 2581.710 3.670 2586.850 4.280 ;
        RECT 2587.690 3.670 2592.830 4.280 ;
        RECT 2593.670 3.670 2598.810 4.280 ;
        RECT 2599.650 3.670 2604.790 4.280 ;
        RECT 2605.630 3.670 2610.770 4.280 ;
        RECT 2611.610 3.670 2616.750 4.280 ;
        RECT 2617.590 3.670 2622.730 4.280 ;
        RECT 2623.570 3.670 2628.710 4.280 ;
        RECT 2629.550 3.670 2634.690 4.280 ;
        RECT 2635.530 3.670 2640.670 4.280 ;
        RECT 2641.510 3.670 2646.650 4.280 ;
        RECT 2647.490 3.670 2652.630 4.280 ;
        RECT 2653.470 3.670 2658.610 4.280 ;
        RECT 2659.450 3.670 2664.590 4.280 ;
        RECT 2665.430 3.670 2670.570 4.280 ;
        RECT 2671.410 3.670 2676.550 4.280 ;
        RECT 2677.390 3.670 2682.530 4.280 ;
        RECT 2683.370 3.670 2688.510 4.280 ;
        RECT 2689.350 3.670 2694.490 4.280 ;
        RECT 2695.330 3.670 2700.470 4.280 ;
        RECT 2701.310 3.670 2706.450 4.280 ;
        RECT 2707.290 3.670 2712.430 4.280 ;
        RECT 2713.270 3.670 2718.410 4.280 ;
        RECT 2719.250 3.670 2724.390 4.280 ;
        RECT 2725.230 3.670 2730.370 4.280 ;
        RECT 2731.210 3.670 2736.350 4.280 ;
        RECT 2737.190 3.670 2742.330 4.280 ;
        RECT 2743.170 3.670 2748.310 4.280 ;
        RECT 2749.150 3.670 2754.290 4.280 ;
        RECT 2755.130 3.670 2760.270 4.280 ;
        RECT 2761.110 3.670 2766.250 4.280 ;
        RECT 2767.090 3.670 2772.230 4.280 ;
        RECT 2773.070 3.670 2778.210 4.280 ;
        RECT 2779.050 3.670 2784.190 4.280 ;
        RECT 2785.030 3.670 2790.170 4.280 ;
        RECT 2791.010 3.670 2796.150 4.280 ;
        RECT 2796.990 3.670 2802.130 4.280 ;
        RECT 2802.970 3.670 2808.110 4.280 ;
        RECT 2808.950 3.670 2814.090 4.280 ;
        RECT 2814.930 3.670 2820.070 4.280 ;
        RECT 2820.910 3.670 2826.050 4.280 ;
        RECT 2826.890 3.670 2832.030 4.280 ;
        RECT 2832.870 3.670 2838.010 4.280 ;
        RECT 2838.850 3.670 2843.990 4.280 ;
        RECT 2844.830 3.670 2849.970 4.280 ;
        RECT 2850.810 3.670 2855.950 4.280 ;
        RECT 2856.790 3.670 2861.930 4.280 ;
        RECT 2862.770 3.670 2867.910 4.280 ;
        RECT 2868.750 3.670 2873.890 4.280 ;
        RECT 2874.730 3.670 2879.870 4.280 ;
        RECT 2880.710 3.670 2885.850 4.280 ;
        RECT 2886.690 3.670 2891.830 4.280 ;
        RECT 2892.670 3.670 2897.810 4.280 ;
        RECT 2898.650 3.670 2903.790 4.280 ;
        RECT 2904.630 3.670 2909.770 4.280 ;
        RECT 2910.610 3.670 2915.750 4.280 ;
        RECT 2916.590 3.670 2917.220 4.280 ;
      LAYER met3 ;
        RECT 2.150 3460.880 2916.000 3508.965 ;
        RECT 4.400 3459.480 2916.000 3460.880 ;
        RECT 2.150 3433.680 2916.000 3459.480 ;
        RECT 2.150 3432.280 2915.600 3433.680 ;
        RECT 2.150 3377.920 2916.000 3432.280 ;
        RECT 4.400 3376.520 2916.000 3377.920 ;
        RECT 2.150 3294.960 2916.000 3376.520 ;
        RECT 4.400 3293.560 2916.000 3294.960 ;
        RECT 2.150 3288.160 2916.000 3293.560 ;
        RECT 2.150 3286.760 2915.600 3288.160 ;
        RECT 2.150 3212.000 2916.000 3286.760 ;
        RECT 4.400 3210.600 2916.000 3212.000 ;
        RECT 2.150 3142.640 2916.000 3210.600 ;
        RECT 2.150 3141.240 2915.600 3142.640 ;
        RECT 2.150 3129.040 2916.000 3141.240 ;
        RECT 4.400 3127.640 2916.000 3129.040 ;
        RECT 2.150 3046.080 2916.000 3127.640 ;
        RECT 4.400 3044.680 2916.000 3046.080 ;
        RECT 2.150 2997.120 2916.000 3044.680 ;
        RECT 2.150 2995.720 2915.600 2997.120 ;
        RECT 2.150 2963.120 2916.000 2995.720 ;
        RECT 4.400 2961.720 2916.000 2963.120 ;
        RECT 2.150 2880.160 2916.000 2961.720 ;
        RECT 4.400 2878.760 2916.000 2880.160 ;
        RECT 2.150 2851.600 2916.000 2878.760 ;
        RECT 2.150 2850.200 2915.600 2851.600 ;
        RECT 2.150 2797.200 2916.000 2850.200 ;
        RECT 4.400 2795.800 2916.000 2797.200 ;
        RECT 2.150 2714.240 2916.000 2795.800 ;
        RECT 4.400 2712.840 2916.000 2714.240 ;
        RECT 2.150 2706.080 2916.000 2712.840 ;
        RECT 2.150 2704.680 2915.600 2706.080 ;
        RECT 2.150 2631.280 2916.000 2704.680 ;
        RECT 4.400 2629.880 2916.000 2631.280 ;
        RECT 2.150 2560.560 2916.000 2629.880 ;
        RECT 2.150 2559.160 2915.600 2560.560 ;
        RECT 2.150 2548.320 2916.000 2559.160 ;
        RECT 4.400 2546.920 2916.000 2548.320 ;
        RECT 2.150 2465.360 2916.000 2546.920 ;
        RECT 4.400 2463.960 2916.000 2465.360 ;
        RECT 2.150 2415.040 2916.000 2463.960 ;
        RECT 2.150 2413.640 2915.600 2415.040 ;
        RECT 2.150 2382.400 2916.000 2413.640 ;
        RECT 4.400 2381.000 2916.000 2382.400 ;
        RECT 2.150 2299.440 2916.000 2381.000 ;
        RECT 4.400 2298.040 2916.000 2299.440 ;
        RECT 2.150 2269.520 2916.000 2298.040 ;
        RECT 2.150 2268.120 2915.600 2269.520 ;
        RECT 2.150 2216.480 2916.000 2268.120 ;
        RECT 4.400 2215.080 2916.000 2216.480 ;
        RECT 2.150 2133.520 2916.000 2215.080 ;
        RECT 4.400 2132.120 2916.000 2133.520 ;
        RECT 2.150 2124.000 2916.000 2132.120 ;
        RECT 2.150 2122.600 2915.600 2124.000 ;
        RECT 2.150 2050.560 2916.000 2122.600 ;
        RECT 4.400 2049.160 2916.000 2050.560 ;
        RECT 2.150 1978.480 2916.000 2049.160 ;
        RECT 2.150 1977.080 2915.600 1978.480 ;
        RECT 2.150 1967.600 2916.000 1977.080 ;
        RECT 4.400 1966.200 2916.000 1967.600 ;
        RECT 2.150 1884.640 2916.000 1966.200 ;
        RECT 4.400 1883.240 2916.000 1884.640 ;
        RECT 2.150 1832.960 2916.000 1883.240 ;
        RECT 2.150 1831.560 2915.600 1832.960 ;
        RECT 2.150 1801.680 2916.000 1831.560 ;
        RECT 4.400 1800.280 2916.000 1801.680 ;
        RECT 2.150 1718.720 2916.000 1800.280 ;
        RECT 4.400 1717.320 2916.000 1718.720 ;
        RECT 2.150 1687.440 2916.000 1717.320 ;
        RECT 2.150 1686.040 2915.600 1687.440 ;
        RECT 2.150 1635.760 2916.000 1686.040 ;
        RECT 4.400 1634.360 2916.000 1635.760 ;
        RECT 2.150 1552.800 2916.000 1634.360 ;
        RECT 4.400 1551.400 2916.000 1552.800 ;
        RECT 2.150 1541.920 2916.000 1551.400 ;
        RECT 2.150 1540.520 2915.600 1541.920 ;
        RECT 2.150 1469.840 2916.000 1540.520 ;
        RECT 4.400 1468.440 2916.000 1469.840 ;
        RECT 2.150 1396.400 2916.000 1468.440 ;
        RECT 2.150 1395.000 2915.600 1396.400 ;
        RECT 2.150 1386.880 2916.000 1395.000 ;
        RECT 4.400 1385.480 2916.000 1386.880 ;
        RECT 2.150 1303.920 2916.000 1385.480 ;
        RECT 4.400 1302.520 2916.000 1303.920 ;
        RECT 2.150 1250.880 2916.000 1302.520 ;
        RECT 2.150 1249.480 2915.600 1250.880 ;
        RECT 2.150 1220.960 2916.000 1249.480 ;
        RECT 4.400 1219.560 2916.000 1220.960 ;
        RECT 2.150 1138.000 2916.000 1219.560 ;
        RECT 4.400 1136.600 2916.000 1138.000 ;
        RECT 2.150 1105.360 2916.000 1136.600 ;
        RECT 2.150 1103.960 2915.600 1105.360 ;
        RECT 2.150 1055.040 2916.000 1103.960 ;
        RECT 4.400 1053.640 2916.000 1055.040 ;
        RECT 2.150 972.080 2916.000 1053.640 ;
        RECT 4.400 970.680 2916.000 972.080 ;
        RECT 2.150 959.840 2916.000 970.680 ;
        RECT 2.150 958.440 2915.600 959.840 ;
        RECT 2.150 889.120 2916.000 958.440 ;
        RECT 4.400 887.720 2916.000 889.120 ;
        RECT 2.150 814.320 2916.000 887.720 ;
        RECT 2.150 812.920 2915.600 814.320 ;
        RECT 2.150 806.160 2916.000 812.920 ;
        RECT 4.400 804.760 2916.000 806.160 ;
        RECT 2.150 723.200 2916.000 804.760 ;
        RECT 4.400 721.800 2916.000 723.200 ;
        RECT 2.150 668.800 2916.000 721.800 ;
        RECT 2.150 667.400 2915.600 668.800 ;
        RECT 2.150 640.240 2916.000 667.400 ;
        RECT 4.400 638.840 2916.000 640.240 ;
        RECT 2.150 557.280 2916.000 638.840 ;
        RECT 4.400 555.880 2916.000 557.280 ;
        RECT 2.150 523.280 2916.000 555.880 ;
        RECT 2.150 521.880 2915.600 523.280 ;
        RECT 2.150 474.320 2916.000 521.880 ;
        RECT 4.400 472.920 2916.000 474.320 ;
        RECT 2.150 391.360 2916.000 472.920 ;
        RECT 4.400 389.960 2916.000 391.360 ;
        RECT 2.150 377.760 2916.000 389.960 ;
        RECT 2.150 376.360 2915.600 377.760 ;
        RECT 2.150 308.400 2916.000 376.360 ;
        RECT 4.400 307.000 2916.000 308.400 ;
        RECT 2.150 232.240 2916.000 307.000 ;
        RECT 2.150 230.840 2915.600 232.240 ;
        RECT 2.150 225.440 2916.000 230.840 ;
        RECT 4.400 224.040 2916.000 225.440 ;
        RECT 2.150 142.480 2916.000 224.040 ;
        RECT 4.400 141.080 2916.000 142.480 ;
        RECT 2.150 86.720 2916.000 141.080 ;
        RECT 2.150 85.320 2915.600 86.720 ;
        RECT 2.150 59.520 2916.000 85.320 ;
        RECT 4.400 58.120 2916.000 59.520 ;
        RECT 2.150 9.695 2916.000 58.120 ;
      LAYER met4 ;
        RECT 15.015 2619.080 53.620 3127.825 ;
        RECT 57.420 2619.080 58.320 3127.825 ;
        RECT 62.120 2619.080 103.620 3127.825 ;
        RECT 107.420 2619.080 108.320 3127.825 ;
        RECT 112.120 2619.080 153.620 3127.825 ;
        RECT 157.420 2619.080 158.320 3127.825 ;
        RECT 162.120 2619.080 203.620 3127.825 ;
        RECT 207.420 2619.700 208.320 3127.825 ;
        RECT 212.120 2619.700 253.620 3127.825 ;
        RECT 257.420 2619.700 258.320 3127.825 ;
        RECT 262.120 2619.700 303.620 3127.825 ;
        RECT 207.420 2619.080 303.620 2619.700 ;
        RECT 307.420 2619.700 308.320 3127.825 ;
        RECT 312.120 2619.700 353.620 3127.825 ;
        RECT 357.420 2619.700 358.320 3127.825 ;
        RECT 362.120 2619.700 403.620 3127.825 ;
        RECT 307.420 2619.080 403.620 2619.700 ;
        RECT 407.420 2619.080 408.320 3127.825 ;
        RECT 412.120 2619.080 453.620 3127.825 ;
        RECT 457.420 2619.080 458.320 3127.825 ;
        RECT 462.120 2619.080 503.620 3127.825 ;
        RECT 507.420 2619.080 508.320 3127.825 ;
        RECT 512.120 2619.080 553.620 3127.825 ;
        RECT 15.015 2202.420 553.620 2619.080 ;
        RECT 15.015 9.695 53.620 2202.420 ;
        RECT 57.420 9.695 58.320 2202.420 ;
        RECT 62.120 9.695 103.620 2202.420 ;
        RECT 107.420 9.695 108.320 2202.420 ;
        RECT 112.120 2201.800 158.320 2202.420 ;
        RECT 112.120 1938.040 153.620 2201.800 ;
        RECT 157.420 1938.040 158.320 2201.800 ;
        RECT 112.120 1930.825 158.320 1938.040 ;
        RECT 162.120 2201.800 353.620 2202.420 ;
        RECT 162.120 1930.825 203.620 2201.800 ;
        RECT 112.120 408.815 203.620 1930.825 ;
        RECT 112.120 405.000 158.320 408.815 ;
        RECT 112.120 9.695 153.620 405.000 ;
        RECT 157.420 9.695 158.320 405.000 ;
        RECT 162.120 9.695 203.620 408.815 ;
        RECT 207.420 1939.665 208.320 2201.800 ;
        RECT 212.120 1939.665 253.620 2201.800 ;
        RECT 257.420 1939.665 258.320 2201.800 ;
        RECT 262.120 1995.520 303.620 2201.800 ;
        RECT 307.420 1995.520 308.320 2201.800 ;
        RECT 262.120 1978.785 308.320 1995.520 ;
        RECT 312.120 1978.785 353.620 2201.800 ;
        RECT 357.420 2201.800 403.620 2202.420 ;
        RECT 357.420 1995.520 358.320 2201.800 ;
        RECT 362.120 1995.520 403.620 2201.800 ;
        RECT 357.420 1978.785 403.620 1995.520 ;
        RECT 262.120 1939.665 403.620 1978.785 ;
        RECT 407.420 1939.665 408.320 2202.420 ;
        RECT 412.120 1939.665 453.620 2202.420 ;
        RECT 207.420 401.335 453.620 1939.665 ;
        RECT 207.420 9.695 208.320 401.335 ;
        RECT 212.120 9.695 253.620 401.335 ;
        RECT 257.420 9.695 258.320 401.335 ;
        RECT 262.120 345.440 308.320 401.335 ;
        RECT 262.120 9.695 303.620 345.440 ;
        RECT 307.420 9.695 308.320 345.440 ;
        RECT 312.120 9.695 353.620 401.335 ;
        RECT 357.420 354.015 453.620 401.335 ;
        RECT 357.420 345.440 403.620 354.015 ;
        RECT 357.420 9.695 358.320 345.440 ;
        RECT 362.120 9.695 403.620 345.440 ;
        RECT 407.420 9.695 408.320 354.015 ;
        RECT 412.120 9.695 453.620 354.015 ;
        RECT 457.420 1939.665 458.320 2202.420 ;
        RECT 462.120 1939.665 503.620 2202.420 ;
        RECT 507.420 1939.665 508.320 2202.420 ;
        RECT 512.120 1995.520 553.620 2202.420 ;
        RECT 557.420 1995.520 558.320 3127.825 ;
        RECT 512.120 1978.785 558.320 1995.520 ;
        RECT 562.120 1978.785 603.620 3127.825 ;
        RECT 607.420 1995.520 608.320 3127.825 ;
        RECT 612.120 1995.520 653.620 3127.825 ;
        RECT 607.420 1978.785 653.620 1995.520 ;
        RECT 512.120 1939.665 653.620 1978.785 ;
        RECT 657.420 1939.665 658.320 3127.825 ;
        RECT 662.120 1939.665 703.620 3127.825 ;
        RECT 457.420 401.335 703.620 1939.665 ;
        RECT 457.420 9.695 458.320 401.335 ;
        RECT 462.120 9.695 503.620 401.335 ;
        RECT 507.420 9.695 508.320 401.335 ;
        RECT 512.120 345.440 558.320 401.335 ;
        RECT 512.120 9.695 553.620 345.440 ;
        RECT 557.420 9.695 558.320 345.440 ;
        RECT 562.120 9.695 603.620 401.335 ;
        RECT 607.420 354.015 703.620 401.335 ;
        RECT 607.420 345.440 653.620 354.015 ;
        RECT 607.420 9.695 608.320 345.440 ;
        RECT 612.120 9.695 653.620 345.440 ;
        RECT 657.420 9.695 658.320 354.015 ;
        RECT 662.120 9.695 703.620 354.015 ;
        RECT 707.420 1939.665 708.320 3127.825 ;
        RECT 712.120 1939.665 753.620 3127.825 ;
        RECT 757.420 1939.665 758.320 3127.825 ;
        RECT 762.120 1995.520 803.620 3127.825 ;
        RECT 807.420 1995.520 808.320 3127.825 ;
        RECT 762.120 1978.785 808.320 1995.520 ;
        RECT 812.120 1978.785 853.620 3127.825 ;
        RECT 857.420 1995.520 858.320 3127.825 ;
        RECT 862.120 1995.520 903.620 3127.825 ;
        RECT 857.420 1978.785 903.620 1995.520 ;
        RECT 762.120 1939.665 903.620 1978.785 ;
        RECT 907.420 1939.665 908.320 3127.825 ;
        RECT 912.120 1939.665 953.620 3127.825 ;
        RECT 957.420 1939.665 958.320 3127.825 ;
        RECT 962.120 1995.520 1003.620 3127.825 ;
        RECT 1007.420 1995.520 1008.320 3127.825 ;
        RECT 962.120 1939.665 1008.320 1995.520 ;
        RECT 1012.120 1978.785 1053.620 3127.825 ;
        RECT 1057.420 1995.520 1058.320 3127.825 ;
        RECT 1062.120 1995.520 1103.620 3127.825 ;
        RECT 1057.420 1978.785 1103.620 1995.520 ;
        RECT 1107.420 1978.785 1108.320 3127.825 ;
        RECT 1112.120 1978.785 1153.620 3127.825 ;
        RECT 1012.120 1939.665 1153.620 1978.785 ;
        RECT 1157.420 1939.665 1158.320 3127.825 ;
        RECT 1162.120 1939.665 1203.620 3127.825 ;
        RECT 1207.420 1939.665 1208.320 3127.825 ;
        RECT 1212.120 1939.665 1253.620 3127.825 ;
        RECT 1257.420 1939.665 1258.320 3127.825 ;
        RECT 1262.120 1995.520 1303.620 3127.825 ;
        RECT 1307.420 1995.520 1308.320 3127.825 ;
        RECT 1262.120 1978.785 1308.320 1995.520 ;
        RECT 1312.120 1995.520 1353.620 3127.825 ;
        RECT 1357.420 1995.520 1358.320 3127.825 ;
        RECT 1362.120 1995.520 1403.620 3127.825 ;
        RECT 1312.120 1978.785 1403.620 1995.520 ;
        RECT 1262.120 1939.665 1403.620 1978.785 ;
        RECT 1407.420 1995.520 1408.320 3127.825 ;
        RECT 1412.120 1995.520 1453.620 3127.825 ;
        RECT 1407.420 1939.665 1453.620 1995.520 ;
        RECT 1457.420 1939.665 1458.320 3127.825 ;
        RECT 1462.120 1939.665 1503.620 3127.825 ;
        RECT 1507.420 1939.665 1508.320 3127.825 ;
        RECT 1512.120 1978.785 1553.620 3127.825 ;
        RECT 1557.420 1978.785 1558.320 3127.825 ;
        RECT 1562.120 1978.785 1603.620 3127.825 ;
        RECT 1512.120 1939.665 1603.620 1978.785 ;
        RECT 1607.420 1939.665 1608.320 3127.825 ;
        RECT 1612.120 1995.520 1653.620 3127.825 ;
        RECT 1657.420 1995.520 1658.320 3127.825 ;
        RECT 1612.120 1939.665 1658.320 1995.520 ;
        RECT 1662.120 1995.520 1703.620 3127.825 ;
        RECT 1707.420 1995.520 1708.320 3127.825 ;
        RECT 1662.120 1939.665 1708.320 1995.520 ;
        RECT 1712.120 1978.785 1753.620 3127.825 ;
        RECT 1757.420 1995.520 1758.320 3127.825 ;
        RECT 1762.120 1995.520 1803.620 3127.825 ;
        RECT 1757.420 1978.785 1803.620 1995.520 ;
        RECT 1807.420 1978.785 1808.320 3127.825 ;
        RECT 1812.120 1978.785 1853.620 3127.825 ;
        RECT 1712.120 1939.665 1853.620 1978.785 ;
        RECT 1857.420 1939.665 1858.320 3127.825 ;
        RECT 1862.120 1939.665 1903.620 3127.825 ;
        RECT 1907.420 1939.665 1908.320 3127.825 ;
        RECT 707.420 401.335 1908.320 1939.665 ;
        RECT 707.420 9.695 708.320 401.335 ;
        RECT 712.120 9.695 753.620 401.335 ;
        RECT 757.420 9.695 758.320 401.335 ;
        RECT 762.120 345.440 808.320 401.335 ;
        RECT 762.120 9.695 803.620 345.440 ;
        RECT 807.420 9.695 808.320 345.440 ;
        RECT 812.120 9.695 853.620 401.335 ;
        RECT 857.420 354.015 953.620 401.335 ;
        RECT 857.420 345.440 903.620 354.015 ;
        RECT 857.420 9.695 858.320 345.440 ;
        RECT 862.120 9.695 903.620 345.440 ;
        RECT 907.420 9.695 908.320 354.015 ;
        RECT 912.120 9.695 953.620 354.015 ;
        RECT 957.420 9.695 958.320 401.335 ;
        RECT 962.120 345.440 1008.320 401.335 ;
        RECT 962.120 9.695 1003.620 345.440 ;
        RECT 1007.420 9.695 1008.320 345.440 ;
        RECT 1012.120 9.695 1053.620 401.335 ;
        RECT 1057.420 345.440 1103.620 401.335 ;
        RECT 1057.420 9.695 1058.320 345.440 ;
        RECT 1062.120 9.695 1103.620 345.440 ;
        RECT 1107.420 9.695 1108.320 401.335 ;
        RECT 1112.120 9.695 1153.620 401.335 ;
        RECT 1157.420 9.695 1158.320 401.335 ;
        RECT 1162.120 9.695 1203.620 401.335 ;
        RECT 1207.420 9.695 1208.320 401.335 ;
        RECT 1212.120 9.695 1253.620 401.335 ;
        RECT 1257.420 9.695 1258.320 401.335 ;
        RECT 1262.120 345.440 1308.320 401.335 ;
        RECT 1262.120 9.695 1303.620 345.440 ;
        RECT 1307.420 9.695 1308.320 345.440 ;
        RECT 1312.120 345.440 1403.620 401.335 ;
        RECT 1312.120 9.695 1353.620 345.440 ;
        RECT 1357.420 9.695 1358.320 345.440 ;
        RECT 1362.120 9.695 1403.620 345.440 ;
        RECT 1407.420 345.440 1453.620 401.335 ;
        RECT 1407.420 9.695 1408.320 345.440 ;
        RECT 1412.120 9.695 1453.620 345.440 ;
        RECT 1457.420 9.695 1458.320 401.335 ;
        RECT 1462.120 9.695 1503.620 401.335 ;
        RECT 1507.420 9.695 1508.320 401.335 ;
        RECT 1512.120 9.695 1553.620 401.335 ;
        RECT 1557.420 9.695 1558.320 401.335 ;
        RECT 1562.120 354.015 1658.320 401.335 ;
        RECT 1562.120 9.695 1603.620 354.015 ;
        RECT 1607.420 9.695 1608.320 354.015 ;
        RECT 1612.120 345.440 1658.320 354.015 ;
        RECT 1612.120 9.695 1653.620 345.440 ;
        RECT 1657.420 9.695 1658.320 345.440 ;
        RECT 1662.120 345.440 1708.320 401.335 ;
        RECT 1662.120 9.695 1703.620 345.440 ;
        RECT 1707.420 9.695 1708.320 345.440 ;
        RECT 1712.120 9.695 1753.620 401.335 ;
        RECT 1757.420 345.440 1803.620 401.335 ;
        RECT 1757.420 9.695 1758.320 345.440 ;
        RECT 1762.120 9.695 1803.620 345.440 ;
        RECT 1807.420 9.695 1808.320 401.335 ;
        RECT 1812.120 354.015 1903.620 401.335 ;
        RECT 1812.120 9.695 1853.620 354.015 ;
        RECT 1857.420 9.695 1858.320 354.015 ;
        RECT 1862.120 9.695 1903.620 354.015 ;
        RECT 1907.420 9.695 1908.320 401.335 ;
        RECT 1912.120 1939.665 1953.620 3127.825 ;
        RECT 1957.420 1995.520 1958.320 3127.825 ;
        RECT 1962.120 1995.520 2003.620 3127.825 ;
        RECT 1957.420 1939.665 2003.620 1995.520 ;
        RECT 2007.420 1978.785 2008.320 3127.825 ;
        RECT 2012.120 1978.785 2053.620 3127.825 ;
        RECT 2057.420 1978.785 2058.320 3127.825 ;
        RECT 2062.120 1978.785 2103.620 3127.825 ;
        RECT 2007.420 1939.665 2103.620 1978.785 ;
        RECT 2107.420 1939.665 2108.320 3127.825 ;
        RECT 2112.120 1939.665 2153.620 3127.825 ;
        RECT 2157.420 1939.665 2158.320 3127.825 ;
        RECT 2162.120 1995.080 2203.620 3127.825 ;
        RECT 2207.420 1995.080 2208.320 3127.825 ;
        RECT 2162.120 1939.665 2208.320 1995.080 ;
        RECT 1912.120 1934.905 2208.320 1939.665 ;
        RECT 2212.120 1993.985 2253.620 3127.825 ;
        RECT 2257.420 1993.985 2258.320 3127.825 ;
        RECT 2262.120 1995.080 2303.620 3127.825 ;
        RECT 2307.420 1995.080 2308.320 3127.825 ;
        RECT 2312.120 1995.080 2353.620 3127.825 ;
        RECT 2262.120 1993.985 2353.620 1995.080 ;
        RECT 2212.120 1934.905 2353.620 1993.985 ;
        RECT 1912.120 405.415 2353.620 1934.905 ;
        RECT 1912.120 401.335 2208.320 405.415 ;
        RECT 1912.120 9.695 1953.620 401.335 ;
        RECT 1957.420 345.440 2003.620 401.335 ;
        RECT 1957.420 9.695 1958.320 345.440 ;
        RECT 1962.120 9.695 2003.620 345.440 ;
        RECT 2007.420 9.695 2008.320 401.335 ;
        RECT 2012.120 9.695 2053.620 401.335 ;
        RECT 2057.420 9.695 2058.320 401.335 ;
        RECT 2062.120 354.015 2153.620 401.335 ;
        RECT 2062.120 9.695 2103.620 354.015 ;
        RECT 2107.420 9.695 2108.320 354.015 ;
        RECT 2112.120 9.695 2153.620 354.015 ;
        RECT 2157.420 9.695 2158.320 401.335 ;
        RECT 2162.120 340.000 2208.320 401.335 ;
        RECT 2162.120 9.695 2203.620 340.000 ;
        RECT 2207.420 9.695 2208.320 340.000 ;
        RECT 2212.120 9.695 2253.620 405.415 ;
        RECT 2257.420 9.695 2258.320 405.415 ;
        RECT 2262.120 340.000 2353.620 405.415 ;
        RECT 2262.120 9.695 2303.620 340.000 ;
        RECT 2307.420 9.695 2308.320 340.000 ;
        RECT 2312.120 9.695 2353.620 340.000 ;
        RECT 2357.420 9.695 2358.320 3127.825 ;
        RECT 2362.120 1899.080 2403.620 3127.825 ;
        RECT 2407.420 1899.080 2408.320 3127.825 ;
        RECT 2412.120 1899.080 2453.620 3127.825 ;
        RECT 2457.420 1899.080 2458.320 3127.825 ;
        RECT 2462.120 1899.080 2503.620 3127.825 ;
        RECT 2507.420 1899.080 2508.320 3127.825 ;
        RECT 2512.120 1899.700 2553.620 3127.825 ;
        RECT 2557.420 1899.700 2558.320 3127.825 ;
        RECT 2562.120 1899.700 2603.620 3127.825 ;
        RECT 2607.420 1899.700 2608.320 3127.825 ;
        RECT 2612.120 1899.700 2653.620 3127.825 ;
        RECT 2657.420 1899.700 2658.320 3127.825 ;
        RECT 2662.120 1899.700 2703.620 3127.825 ;
        RECT 2707.420 1899.700 2708.320 3127.825 ;
        RECT 2712.120 1899.700 2753.620 3127.825 ;
        RECT 2512.120 1899.080 2753.620 1899.700 ;
        RECT 2757.420 1899.080 2758.320 3127.825 ;
        RECT 2762.120 1899.080 2803.620 3127.825 ;
        RECT 2807.420 1899.080 2808.320 3127.825 ;
        RECT 2812.120 1899.080 2853.620 3127.825 ;
        RECT 2857.420 1899.080 2858.320 3127.825 ;
        RECT 2862.120 1899.080 2873.160 3127.825 ;
        RECT 2362.120 1482.420 2873.160 1899.080 ;
        RECT 2362.120 1379.080 2403.620 1482.420 ;
        RECT 2407.420 1379.080 2408.320 1482.420 ;
        RECT 2412.120 1379.080 2453.620 1482.420 ;
        RECT 2457.420 1379.080 2458.320 1482.420 ;
        RECT 2462.120 1481.800 2753.620 1482.420 ;
        RECT 2462.120 1379.080 2503.620 1481.800 ;
        RECT 2507.420 1379.080 2508.320 1481.800 ;
        RECT 2512.120 1379.700 2553.620 1481.800 ;
        RECT 2557.420 1379.700 2558.320 1481.800 ;
        RECT 2562.120 1379.700 2603.620 1481.800 ;
        RECT 2607.420 1379.700 2608.320 1481.800 ;
        RECT 2612.120 1379.700 2653.620 1481.800 ;
        RECT 2657.420 1379.700 2658.320 1481.800 ;
        RECT 2662.120 1379.700 2703.620 1481.800 ;
        RECT 2707.420 1379.700 2708.320 1481.800 ;
        RECT 2712.120 1379.700 2753.620 1481.800 ;
        RECT 2512.120 1379.080 2753.620 1379.700 ;
        RECT 2757.420 1379.080 2758.320 1482.420 ;
        RECT 2762.120 1481.800 2853.620 1482.420 ;
        RECT 2762.120 1379.080 2803.620 1481.800 ;
        RECT 2807.420 1379.080 2808.320 1481.800 ;
        RECT 2812.120 1379.080 2853.620 1481.800 ;
        RECT 2857.420 1379.080 2858.320 1482.420 ;
        RECT 2862.120 1379.080 2873.160 1482.420 ;
        RECT 2362.120 962.420 2873.160 1379.080 ;
        RECT 2362.120 858.980 2403.620 962.420 ;
        RECT 2407.420 859.080 2408.320 962.420 ;
        RECT 2412.120 859.080 2453.620 962.420 ;
        RECT 2407.420 858.980 2453.620 859.080 ;
        RECT 2457.420 859.080 2458.320 962.420 ;
        RECT 2462.120 961.800 2753.620 962.420 ;
        RECT 2462.120 859.080 2503.620 961.800 ;
        RECT 2457.420 858.980 2503.620 859.080 ;
        RECT 2507.420 859.080 2508.320 961.800 ;
        RECT 2512.120 859.700 2553.620 961.800 ;
        RECT 2557.420 859.700 2558.320 961.800 ;
        RECT 2562.120 859.700 2603.620 961.800 ;
        RECT 2607.420 859.700 2608.320 961.800 ;
        RECT 2612.120 859.700 2653.620 961.800 ;
        RECT 2657.420 859.700 2658.320 961.800 ;
        RECT 2662.120 859.700 2703.620 961.800 ;
        RECT 2707.420 859.700 2708.320 961.800 ;
        RECT 2712.120 859.700 2753.620 961.800 ;
        RECT 2512.120 859.080 2753.620 859.700 ;
        RECT 2507.420 858.980 2753.620 859.080 ;
        RECT 2757.420 859.080 2758.320 962.420 ;
        RECT 2762.120 961.800 2853.620 962.420 ;
        RECT 2762.120 859.080 2803.620 961.800 ;
        RECT 2757.420 858.980 2803.620 859.080 ;
        RECT 2807.420 859.080 2808.320 961.800 ;
        RECT 2812.120 859.080 2853.620 961.800 ;
        RECT 2807.420 858.980 2853.620 859.080 ;
        RECT 2857.420 859.080 2858.320 962.420 ;
        RECT 2862.120 859.080 2873.160 962.420 ;
        RECT 2857.420 858.980 2873.160 859.080 ;
        RECT 2362.120 442.420 2873.160 858.980 ;
        RECT 2362.120 9.695 2403.620 442.420 ;
        RECT 2407.420 9.695 2408.320 442.420 ;
        RECT 2412.120 9.695 2453.620 442.420 ;
        RECT 2457.420 9.695 2458.320 442.420 ;
        RECT 2462.120 441.800 2753.620 442.420 ;
        RECT 2462.120 9.695 2503.620 441.800 ;
        RECT 2507.420 9.695 2508.320 441.800 ;
        RECT 2512.120 9.695 2553.620 441.800 ;
        RECT 2557.420 9.695 2558.320 441.800 ;
        RECT 2562.120 9.695 2603.620 441.800 ;
        RECT 2607.420 9.695 2608.320 441.800 ;
        RECT 2612.120 9.695 2653.620 441.800 ;
        RECT 2657.420 9.695 2658.320 441.800 ;
        RECT 2662.120 9.695 2703.620 441.800 ;
        RECT 2707.420 9.695 2708.320 441.800 ;
        RECT 2712.120 9.695 2753.620 441.800 ;
        RECT 2757.420 9.695 2758.320 442.420 ;
        RECT 2762.120 441.800 2853.620 442.420 ;
        RECT 2762.120 9.695 2803.620 441.800 ;
        RECT 2807.420 9.695 2808.320 441.800 ;
        RECT 2812.120 9.695 2853.620 441.800 ;
        RECT 2857.420 9.695 2858.320 442.420 ;
        RECT 2862.120 9.695 2873.160 442.420 ;
      LAYER met5 ;
        RECT 48.420 2518.680 2850.500 2535.500 ;
        RECT 48.420 2468.680 2850.500 2507.780 ;
        RECT 48.420 2418.680 2850.500 2457.780 ;
        RECT 48.420 2368.680 2850.500 2407.780 ;
        RECT 48.420 2318.680 2850.500 2357.780 ;
        RECT 48.420 2268.680 2850.500 2307.780 ;
        RECT 48.420 2218.680 2850.500 2257.780 ;
        RECT 48.420 2168.680 2850.500 2207.780 ;
        RECT 48.420 2118.680 2850.500 2157.780 ;
        RECT 48.420 2068.680 2850.500 2107.780 ;
        RECT 48.420 2018.680 2850.500 2057.780 ;
        RECT 48.420 1968.680 2850.500 2007.780 ;
        RECT 48.420 1918.680 2850.500 1957.780 ;
        RECT 48.420 1868.680 2850.500 1907.780 ;
        RECT 48.420 1818.680 2850.500 1857.780 ;
        RECT 48.420 1768.680 2850.500 1807.780 ;
        RECT 48.420 1718.680 2850.500 1757.780 ;
        RECT 48.420 1668.680 2850.500 1707.780 ;
        RECT 48.420 1618.680 2850.500 1657.780 ;
        RECT 48.420 1568.680 2850.500 1607.780 ;
        RECT 48.420 1518.680 2850.500 1557.780 ;
        RECT 48.420 1468.680 2850.500 1507.780 ;
        RECT 48.420 1418.680 2850.500 1457.780 ;
        RECT 48.420 1368.680 2850.500 1407.780 ;
        RECT 48.420 1318.680 2850.500 1357.780 ;
        RECT 48.420 1268.680 2850.500 1307.780 ;
        RECT 48.420 1218.680 2850.500 1257.780 ;
        RECT 48.420 1168.680 2850.500 1207.780 ;
        RECT 48.420 1118.680 2850.500 1157.780 ;
        RECT 48.420 1068.680 2850.500 1107.780 ;
        RECT 48.420 1018.680 2850.500 1057.780 ;
        RECT 48.420 968.680 2850.500 1007.780 ;
        RECT 48.420 918.680 2850.500 957.780 ;
        RECT 48.420 868.680 2850.500 907.780 ;
        RECT 48.420 818.680 2850.500 857.780 ;
        RECT 48.420 768.680 2850.500 807.780 ;
        RECT 48.420 718.680 2850.500 757.780 ;
        RECT 48.420 668.680 2850.500 707.780 ;
        RECT 48.420 618.680 2850.500 657.780 ;
        RECT 48.420 568.680 2850.500 607.780 ;
        RECT 48.420 518.680 2850.500 557.780 ;
        RECT 48.420 468.680 2850.500 507.780 ;
        RECT 48.420 418.680 2850.500 457.780 ;
        RECT 48.420 388.500 2850.500 407.780 ;
  END
END summer_school_top_wrapper
END LIBRARY

