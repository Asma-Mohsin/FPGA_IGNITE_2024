VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BlockRAM_1KB
  CLASS BLOCK ;
  FOREIGN BlockRAM_1KB ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 455.230 ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 1.000 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 1.000 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 1.000 398.440 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 1.000 395.040 ;
    END
  END C3
  PIN C4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 1.000 ;
    END
  END C4
  PIN C5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 1.000 391.640 ;
    END
  END C5
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 1.000 418.840 ;
    END
  END clk
  PIN rd_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 447.670 454.230 447.950 455.230 ;
    END
  END rd_addr[0]
  PIN rd_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 599.000 119.040 600.000 119.640 ;
    END
  END rd_addr[1]
  PIN rd_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 599.000 108.840 600.000 109.440 ;
    END
  END rd_addr[2]
  PIN rd_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 599.000 102.040 600.000 102.640 ;
    END
  END rd_addr[3]
  PIN rd_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 1.000 ;
    END
  END rd_addr[4]
  PIN rd_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 1.000 ;
    END
  END rd_addr[5]
  PIN rd_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 463.770 0.000 464.050 1.000 ;
    END
  END rd_addr[6]
  PIN rd_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 1.000 ;
    END
  END rd_addr[7]
  PIN rd_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 1.000 354.240 ;
    END
  END rd_data[0]
  PIN rd_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 1.000 337.240 ;
    END
  END rd_data[10]
  PIN rd_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 1.000 344.040 ;
    END
  END rd_data[11]
  PIN rd_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 483.090 454.230 483.370 455.230 ;
    END
  END rd_data[12]
  PIN rd_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 599.000 414.840 600.000 415.440 ;
    END
  END rd_data[13]
  PIN rd_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 599.000 428.440 600.000 429.040 ;
    END
  END rd_data[14]
  PIN rd_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 454.230 96.970 455.230 ;
    END
  END rd_data[15]
  PIN rd_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 1.000 347.440 ;
    END
  END rd_data[16]
  PIN rd_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 1.000 439.240 ;
    END
  END rd_data[17]
  PIN rd_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 1.000 408.640 ;
    END
  END rd_data[18]
  PIN rd_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 1.000 364.440 ;
    END
  END rd_data[19]
  PIN rd_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 1.000 381.440 ;
    END
  END rd_data[1]
  PIN rd_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 1.000 422.240 ;
    END
  END rd_data[20]
  PIN rd_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 1.000 401.840 ;
    END
  END rd_data[21]
  PIN rd_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 1.000 432.440 ;
    END
  END rd_data[22]
  PIN rd_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 1.000 415.440 ;
    END
  END rd_data[23]
  PIN rd_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 1.000 384.840 ;
    END
  END rd_data[24]
  PIN rd_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 1.000 435.840 ;
    END
  END rd_data[25]
  PIN rd_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 1.000 412.040 ;
    END
  END rd_data[26]
  PIN rd_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 1.000 388.240 ;
    END
  END rd_data[27]
  PIN rd_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 1.000 429.040 ;
    END
  END rd_data[28]
  PIN rd_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 1.000 374.640 ;
    END
  END rd_data[29]
  PIN rd_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 1.000 357.640 ;
    END
  END rd_data[2]
  PIN rd_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 1.000 405.240 ;
    END
  END rd_data[30]
  PIN rd_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 1.000 425.640 ;
    END
  END rd_data[31]
  PIN rd_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 1.000 371.240 ;
    END
  END rd_data[3]
  PIN rd_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 1.000 361.040 ;
    END
  END rd_data[4]
  PIN rd_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 1.000 340.640 ;
    END
  END rd_data[5]
  PIN rd_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 1.000 378.040 ;
    END
  END rd_data[6]
  PIN rd_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 1.000 367.840 ;
    END
  END rd_data[7]
  PIN rd_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 1.000 327.040 ;
    END
  END rd_data[8]
  PIN rd_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 1.000 350.840 ;
    END
  END rd_data[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 25.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 594.560 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 594.560 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 594.560 334.690 ;
    END
    PORT
      LAYER met4 ;
        RECT 564.540 21.520 566.140 443.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.040 14.500 594.560 16.100 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 25.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 25.320 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 594.560 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 594.560 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 594.560 337.990 ;
    END
    PORT
      LAYER met4 ;
        RECT 568.220 21.520 569.820 443.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 21.040 17.900 594.560 19.500 ;
    END
  END vssd1
  PIN wr_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 1.000 ;
    END
  END wr_addr[0]
  PIN wr_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 1.000 163.840 ;
    END
  END wr_addr[1]
  PIN wr_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 1.000 174.040 ;
    END
  END wr_addr[2]
  PIN wr_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 1.000 177.440 ;
    END
  END wr_addr[3]
  PIN wr_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 1.000 184.240 ;
    END
  END wr_addr[4]
  PIN wr_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 1.000 191.040 ;
    END
  END wr_addr[5]
  PIN wr_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 1.000 201.240 ;
    END
  END wr_addr[6]
  PIN wr_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 1.000 204.640 ;
    END
  END wr_addr[7]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 1.000 ;
    END
  END wr_data[0]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 1.000 ;
    END
  END wr_data[10]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 1.000 ;
    END
  END wr_data[11]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 1.000 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 1.000 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 1.000 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 1.000 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 1.000 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 1.000 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 1.000 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 1.000 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 1.000 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 1.000 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 1.000 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 1.000 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 1.000 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 1.000 160.440 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 1.000 170.640 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 1.000 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 1.000 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 1.000 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 1.000 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 1.000 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 1.000 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 1.000 ;
    END
  END wr_data[31]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 1.000 ;
    END
  END wr_data[3]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 1.000 ;
    END
  END wr_data[4]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 1.000 ;
    END
  END wr_data[5]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 1.000 ;
    END
  END wr_data[6]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 1.000 ;
    END
  END wr_data[7]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 1.000 ;
    END
  END wr_data[8]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 1.000 ;
    END
  END wr_data[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 443.445 ;
      LAYER met1 ;
        RECT 3.750 10.640 594.320 454.880 ;
      LAYER met2 ;
        RECT 3.770 453.950 96.410 454.910 ;
        RECT 97.250 453.950 447.390 454.910 ;
        RECT 448.230 453.950 482.810 454.910 ;
        RECT 483.650 453.950 592.850 454.910 ;
        RECT 3.770 1.280 592.850 453.950 ;
        RECT 3.770 0.270 109.290 1.280 ;
        RECT 110.130 0.270 112.510 1.280 ;
        RECT 113.350 0.270 128.610 1.280 ;
        RECT 129.450 0.270 157.590 1.280 ;
        RECT 158.430 0.270 164.030 1.280 ;
        RECT 164.870 0.270 167.250 1.280 ;
        RECT 168.090 0.270 170.470 1.280 ;
        RECT 171.310 0.270 173.690 1.280 ;
        RECT 174.530 0.270 176.910 1.280 ;
        RECT 177.750 0.270 180.130 1.280 ;
        RECT 180.970 0.270 183.350 1.280 ;
        RECT 184.190 0.270 186.570 1.280 ;
        RECT 187.410 0.270 189.790 1.280 ;
        RECT 190.630 0.270 193.010 1.280 ;
        RECT 193.850 0.270 196.230 1.280 ;
        RECT 197.070 0.270 199.450 1.280 ;
        RECT 200.290 0.270 202.670 1.280 ;
        RECT 203.510 0.270 205.890 1.280 ;
        RECT 206.730 0.270 209.110 1.280 ;
        RECT 209.950 0.270 212.330 1.280 ;
        RECT 213.170 0.270 215.550 1.280 ;
        RECT 216.390 0.270 218.770 1.280 ;
        RECT 219.610 0.270 221.990 1.280 ;
        RECT 222.830 0.270 225.210 1.280 ;
        RECT 226.050 0.270 228.430 1.280 ;
        RECT 229.270 0.270 231.650 1.280 ;
        RECT 232.490 0.270 234.870 1.280 ;
        RECT 235.710 0.270 238.090 1.280 ;
        RECT 238.930 0.270 241.310 1.280 ;
        RECT 242.150 0.270 244.530 1.280 ;
        RECT 245.370 0.270 247.750 1.280 ;
        RECT 248.590 0.270 250.970 1.280 ;
        RECT 251.810 0.270 254.190 1.280 ;
        RECT 255.030 0.270 260.630 1.280 ;
        RECT 261.470 0.270 460.270 1.280 ;
        RECT 461.110 0.270 463.490 1.280 ;
        RECT 464.330 0.270 466.710 1.280 ;
        RECT 467.550 0.270 469.930 1.280 ;
        RECT 470.770 0.270 592.850 1.280 ;
      LAYER met3 ;
        RECT 1.000 439.640 599.000 443.525 ;
        RECT 1.400 438.240 599.000 439.640 ;
        RECT 1.000 436.240 599.000 438.240 ;
        RECT 1.400 434.840 599.000 436.240 ;
        RECT 1.000 432.840 599.000 434.840 ;
        RECT 1.400 431.440 599.000 432.840 ;
        RECT 1.000 429.440 599.000 431.440 ;
        RECT 1.400 428.040 598.600 429.440 ;
        RECT 1.000 426.040 599.000 428.040 ;
        RECT 1.400 424.640 599.000 426.040 ;
        RECT 1.000 422.640 599.000 424.640 ;
        RECT 1.400 421.240 599.000 422.640 ;
        RECT 1.000 419.240 599.000 421.240 ;
        RECT 1.400 417.840 599.000 419.240 ;
        RECT 1.000 415.840 599.000 417.840 ;
        RECT 1.400 414.440 598.600 415.840 ;
        RECT 1.000 412.440 599.000 414.440 ;
        RECT 1.400 411.040 599.000 412.440 ;
        RECT 1.000 409.040 599.000 411.040 ;
        RECT 1.400 407.640 599.000 409.040 ;
        RECT 1.000 405.640 599.000 407.640 ;
        RECT 1.400 404.240 599.000 405.640 ;
        RECT 1.000 402.240 599.000 404.240 ;
        RECT 1.400 400.840 599.000 402.240 ;
        RECT 1.000 398.840 599.000 400.840 ;
        RECT 1.400 397.440 599.000 398.840 ;
        RECT 1.000 395.440 599.000 397.440 ;
        RECT 1.400 394.040 599.000 395.440 ;
        RECT 1.000 392.040 599.000 394.040 ;
        RECT 1.400 390.640 599.000 392.040 ;
        RECT 1.000 388.640 599.000 390.640 ;
        RECT 1.400 387.240 599.000 388.640 ;
        RECT 1.000 385.240 599.000 387.240 ;
        RECT 1.400 383.840 599.000 385.240 ;
        RECT 1.000 381.840 599.000 383.840 ;
        RECT 1.400 380.440 599.000 381.840 ;
        RECT 1.000 378.440 599.000 380.440 ;
        RECT 1.400 377.040 599.000 378.440 ;
        RECT 1.000 375.040 599.000 377.040 ;
        RECT 1.400 373.640 599.000 375.040 ;
        RECT 1.000 371.640 599.000 373.640 ;
        RECT 1.400 370.240 599.000 371.640 ;
        RECT 1.000 368.240 599.000 370.240 ;
        RECT 1.400 366.840 599.000 368.240 ;
        RECT 1.000 364.840 599.000 366.840 ;
        RECT 1.400 363.440 599.000 364.840 ;
        RECT 1.000 361.440 599.000 363.440 ;
        RECT 1.400 360.040 599.000 361.440 ;
        RECT 1.000 358.040 599.000 360.040 ;
        RECT 1.400 356.640 599.000 358.040 ;
        RECT 1.000 354.640 599.000 356.640 ;
        RECT 1.400 353.240 599.000 354.640 ;
        RECT 1.000 351.240 599.000 353.240 ;
        RECT 1.400 349.840 599.000 351.240 ;
        RECT 1.000 347.840 599.000 349.840 ;
        RECT 1.400 346.440 599.000 347.840 ;
        RECT 1.000 344.440 599.000 346.440 ;
        RECT 1.400 343.040 599.000 344.440 ;
        RECT 1.000 341.040 599.000 343.040 ;
        RECT 1.400 339.640 599.000 341.040 ;
        RECT 1.000 337.640 599.000 339.640 ;
        RECT 1.400 336.240 599.000 337.640 ;
        RECT 1.000 327.440 599.000 336.240 ;
        RECT 1.400 326.040 599.000 327.440 ;
        RECT 1.000 205.040 599.000 326.040 ;
        RECT 1.400 203.640 599.000 205.040 ;
        RECT 1.000 201.640 599.000 203.640 ;
        RECT 1.400 200.240 599.000 201.640 ;
        RECT 1.000 191.440 599.000 200.240 ;
        RECT 1.400 190.040 599.000 191.440 ;
        RECT 1.000 184.640 599.000 190.040 ;
        RECT 1.400 183.240 599.000 184.640 ;
        RECT 1.000 177.840 599.000 183.240 ;
        RECT 1.400 176.440 599.000 177.840 ;
        RECT 1.000 174.440 599.000 176.440 ;
        RECT 1.400 173.040 599.000 174.440 ;
        RECT 1.000 171.040 599.000 173.040 ;
        RECT 1.400 169.640 599.000 171.040 ;
        RECT 1.000 164.240 599.000 169.640 ;
        RECT 1.400 162.840 599.000 164.240 ;
        RECT 1.000 160.840 599.000 162.840 ;
        RECT 1.400 159.440 599.000 160.840 ;
        RECT 1.000 120.040 599.000 159.440 ;
        RECT 1.000 118.640 598.600 120.040 ;
        RECT 1.000 109.840 599.000 118.640 ;
        RECT 1.000 108.440 598.600 109.840 ;
        RECT 1.000 103.040 599.000 108.440 ;
        RECT 1.000 101.640 598.600 103.040 ;
        RECT 1.000 10.715 599.000 101.640 ;
      LAYER met4 ;
        RECT 18.695 20.575 20.640 442.505 ;
        RECT 23.040 20.575 23.940 442.505 ;
        RECT 26.340 25.720 529.160 442.505 ;
        RECT 26.340 24.885 177.540 25.720 ;
        RECT 26.340 20.575 174.240 24.885 ;
        RECT 176.640 20.575 177.540 24.885 ;
        RECT 179.940 24.885 481.440 25.720 ;
        RECT 179.940 20.575 327.840 24.885 ;
        RECT 330.240 24.800 481.440 24.885 ;
        RECT 330.240 20.575 331.140 24.800 ;
        RECT 333.540 20.575 481.440 24.800 ;
        RECT 483.840 20.575 484.740 25.720 ;
        RECT 487.140 20.575 529.160 25.720 ;
  END
END BlockRAM_1KB
END LIBRARY

