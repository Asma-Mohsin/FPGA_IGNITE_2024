VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_IO
  CLASS BLOCK ;
  FOREIGN RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 223.115 ;
  PIN Config_accessC_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 45.600 130.000 46.200 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 48.320 130.000 48.920 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 51.040 130.000 51.640 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 53.760 130.000 54.360 ;
    END
  END Config_accessC_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.800 84.960 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 0.800 86.320 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 0.800 88.360 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 0.800 89.720 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 0.800 105.360 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 0.800 107.400 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 0.800 108.760 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 0.800 110.800 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 0.800 112.840 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 0.800 114.200 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 0.800 116.240 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 0.800 117.600 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 0.800 91.760 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 0.800 93.120 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 0.800 95.160 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 0.800 96.520 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 0.800 98.560 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 0.800 100.600 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 0.800 101.960 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.800 104.000 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.800 147.520 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 0.800 164.520 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 0.800 166.560 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 0.800 148.880 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 0.800 150.920 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 0.800 152.280 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 0.800 154.320 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 0.800 156.360 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 0.800 157.720 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 0.800 159.760 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 0.800 161.120 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 0.800 163.160 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 0.800 119.640 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 0.800 136.640 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 0.800 138.680 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 0.800 140.720 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 0.800 142.080 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 0.800 144.120 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 0.800 145.480 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 0.800 121.000 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 0.800 123.040 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 0.800 124.400 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 0.800 126.440 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.800 128.480 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 0.800 129.840 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 0.800 131.880 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 0.800 133.240 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 0.800 135.280 ;
    END
  END EE4END[9]
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 78.920 130.000 79.520 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 81.640 130.000 82.240 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 85.040 130.000 85.640 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 87.760 130.000 88.360 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 68.040 130.000 68.640 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 70.760 130.000 71.360 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 73.480 130.000 74.080 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 76.200 130.000 76.800 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 57.160 130.000 57.760 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 59.880 130.000 60.480 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 62.600 130.000 63.200 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 65.320 130.000 65.920 ;
    END
  END FAB2RAM_C_O3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 123.800 130.000 124.400 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 126.520 130.000 127.120 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 129.240 130.000 129.840 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 131.960 130.000 132.560 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 112.920 130.000 113.520 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 115.640 130.000 116.240 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 118.360 130.000 118.960 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 121.080 130.000 121.680 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 101.360 130.000 101.960 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 104.080 130.000 104.680 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 106.800 130.000 107.400 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 109.520 130.000 110.120 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 90.480 130.000 91.080 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 93.200 130.000 93.800 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 95.920 130.000 96.520 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 98.640 130.000 99.240 ;
    END
  END FAB2RAM_D3_O3
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 0.800 168.600 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 0.800 185.600 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 0.800 187.640 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 0.800 189.000 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 0.800 191.040 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 0.800 192.400 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 0.800 194.440 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.800 196.480 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 0.800 197.840 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 0.800 199.880 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 0.800 201.240 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 0.800 169.960 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 0.800 203.280 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 0.800 204.640 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 0.800 206.680 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 0.800 208.040 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 0.800 210.080 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 0.800 212.120 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 0.800 213.480 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 0.800 215.520 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 0.800 216.880 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 0.800 218.920 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.800 172.000 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 0.800 220.280 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 0.800 222.320 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 0.800 173.360 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 0.800 175.400 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 0.800 176.760 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 0.800 178.800 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 0.800 180.160 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 0.800 182.200 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 0.800 184.240 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 134.680 130.000 135.280 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 162.560 130.000 163.160 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 165.280 130.000 165.880 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 168.680 130.000 169.280 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 171.400 130.000 172.000 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 174.120 130.000 174.720 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 176.840 130.000 177.440 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 179.560 130.000 180.160 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 182.280 130.000 182.880 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 185.000 130.000 185.600 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 187.720 130.000 188.320 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 137.400 130.000 138.000 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 190.440 130.000 191.040 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 193.160 130.000 193.760 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 196.560 130.000 197.160 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 199.280 130.000 199.880 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 202.000 130.000 202.600 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 204.720 130.000 205.320 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 207.440 130.000 208.040 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 210.160 130.000 210.760 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 212.880 130.000 213.480 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 215.600 130.000 216.200 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 140.800 130.000 141.400 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 218.320 130.000 218.920 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 221.040 130.000 221.640 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 143.520 130.000 144.120 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 146.240 130.000 146.840 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 148.960 130.000 149.560 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 151.680 130.000 152.280 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 154.400 130.000 155.000 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 157.120 130.000 157.720 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 159.840 130.000 160.440 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 222.315 102.950 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 222.315 116.750 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 222.315 118.130 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 222.315 119.510 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 222.315 120.890 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 222.315 122.270 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 222.315 123.650 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 222.315 125.030 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 222.315 126.410 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 222.315 127.790 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 222.315 129.170 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 222.315 104.330 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 222.315 105.710 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 222.315 107.090 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 222.315 108.470 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 222.315 109.850 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 222.315 111.230 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 222.315 112.610 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 222.315 113.990 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 222.315 115.370 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 222.315 0.830 223.115 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 222.315 2.210 223.115 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 222.315 3.590 223.115 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 222.315 4.970 223.115 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 0.800 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 0.800 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 0.800 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 0.800 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 222.315 6.350 223.115 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 222.315 7.730 223.115 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 222.315 9.110 223.115 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 222.315 10.490 223.115 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 222.315 11.870 223.115 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 222.315 13.250 223.115 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 222.315 14.630 223.115 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 222.315 16.010 223.115 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 222.315 17.390 223.115 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 222.315 18.770 223.115 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 222.315 20.150 223.115 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 222.315 21.530 223.115 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 222.315 22.910 223.115 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 222.315 24.290 223.115 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 222.315 25.670 223.115 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 222.315 27.050 223.115 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 0.800 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 0.800 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 0.800 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 0.800 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 0.800 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 0.800 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 0.800 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 0.800 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 0.800 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 0.800 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 0.800 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 0.800 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 0.800 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 0.800 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 0.800 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 0.800 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 222.315 28.430 223.115 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 222.315 42.690 223.115 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 222.315 44.070 223.115 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 222.315 45.450 223.115 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 222.315 46.830 223.115 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 222.315 48.210 223.115 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 222.315 49.590 223.115 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 222.315 29.810 223.115 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 222.315 31.190 223.115 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 222.315 32.570 223.115 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 222.315 34.410 223.115 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 222.315 35.790 223.115 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 222.315 37.170 223.115 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 222.315 38.550 223.115 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 222.315 39.930 223.115 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 222.315 41.310 223.115 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 0.800 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 0.800 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.800 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 0.800 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 0.800 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 0.800 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 0.800 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 0.800 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 0.800 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 0.800 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 0.800 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 0.800 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 0.800 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 0.800 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.800 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 0.800 ;
    END
  END N4END[9]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 34.720 130.000 35.320 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 37.440 130.000 38.040 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 40.160 130.000 40.760 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 42.880 130.000 43.480 ;
    END
  END RAM2FAB_D0_I3
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 23.160 130.000 23.760 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 25.880 130.000 26.480 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 29.280 130.000 29.880 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 32.000 130.000 32.600 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 12.280 130.000 12.880 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 15.000 130.000 15.600 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 17.720 130.000 18.320 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 20.440 130.000 21.040 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 1.400 130.000 2.000 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 4.120 130.000 4.720 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 6.840 130.000 7.440 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.200 9.560 130.000 10.160 ;
    END
  END RAM2FAB_D3_I3
  PIN S1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 0.800 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 0.800 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 0.800 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 0.800 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 222.315 50.970 223.115 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 222.315 52.350 223.115 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 222.315 53.730 223.115 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 222.315 55.110 223.115 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 0.800 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 0.800 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 0.800 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 0.800 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 0.800 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 0.800 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 0.800 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 0.800 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 0.800 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 0.800 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.800 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 0.800 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 0.800 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 0.800 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 0.800 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 0.800 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 222.315 56.490 223.115 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 222.315 57.870 223.115 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 222.315 59.250 223.115 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 222.315 60.630 223.115 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 222.315 62.010 223.115 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 222.315 63.390 223.115 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 222.315 64.770 223.115 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 222.315 66.610 223.115 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 222.315 67.990 223.115 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 222.315 69.370 223.115 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 222.315 70.750 223.115 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 222.315 72.130 223.115 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 222.315 73.510 223.115 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 222.315 74.890 223.115 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 222.315 76.270 223.115 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 222.315 77.650 223.115 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 0.800 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 0.800 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 0.800 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 0.800 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 0.800 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 0.800 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 0.800 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 0.800 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 0.800 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 0.800 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 0.800 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 0.800 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 0.800 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 0.800 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 0.800 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 0.800 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 222.315 79.030 223.115 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 222.315 92.830 223.115 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 222.315 94.210 223.115 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 222.315 95.590 223.115 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 222.315 96.970 223.115 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 222.315 98.810 223.115 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 222.315 100.190 223.115 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 222.315 80.410 223.115 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 222.315 81.790 223.115 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 222.315 83.170 223.115 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 222.315 84.550 223.115 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 222.315 85.930 223.115 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 222.315 87.310 223.115 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 222.315 88.690 223.115 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 222.315 90.070 223.115 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 222.315 91.450 223.115 ;
    END
  END S4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 222.315 101.570 223.115 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 44.370 5.200 45.970 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.025 5.200 85.625 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.545 5.200 26.145 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.195 5.200 65.795 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.850 5.200 105.450 217.840 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 0.800 1.320 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 0.800 2.680 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 0.800 4.720 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 0.800 6.080 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 0.800 8.120 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 0.800 9.480 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 0.800 11.520 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 0.800 12.880 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 0.800 14.920 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 0.800 16.960 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 0.800 18.320 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 0.800 20.360 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 0.800 21.720 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 0.800 23.760 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 0.800 25.120 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 0.800 27.160 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 0.800 29.200 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 0.800 30.560 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 0.800 32.600 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 0.800 33.960 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 0.800 63.880 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 0.800 80.880 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 0.800 82.920 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 0.800 65.240 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 0.800 67.280 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 0.800 68.640 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 0.800 70.680 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 0.800 72.720 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 0.800 74.080 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 0.800 76.120 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 0.800 77.480 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 0.800 79.520 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.800 36.000 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 0.800 53.000 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 0.800 55.040 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 0.800 57.080 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 0.800 58.440 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.800 60.480 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 0.800 61.840 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 0.800 37.360 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 0.800 39.400 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 0.800 40.760 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 0.800 42.800 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 0.800 44.840 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 0.800 46.200 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 0.800 48.240 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 0.800 49.600 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 0.800 51.640 ;
    END
  END WW4BEG[9]
  OBS
      LAYER li1 ;
        RECT 4.285 207.995 130.000 221.595 ;
        RECT 4.285 160.565 130.035 207.995 ;
        RECT 4.285 158.355 130.000 160.565 ;
        RECT 4.285 133.025 130.035 158.355 ;
        RECT 4.285 110.415 130.000 133.025 ;
        RECT 4.285 70.465 130.035 110.415 ;
        RECT 4.285 0.765 130.000 70.465 ;
      LAYER met1 ;
        RECT 0.530 159.020 130.000 221.640 ;
        RECT 0.530 158.200 130.020 159.020 ;
        RECT 0.530 0.040 130.000 158.200 ;
      LAYER met2 ;
        RECT 1.110 222.035 1.650 222.315 ;
        RECT 2.490 222.035 3.030 222.315 ;
        RECT 3.870 222.035 4.410 222.315 ;
        RECT 5.250 222.035 5.790 222.315 ;
        RECT 6.630 222.035 7.170 222.315 ;
        RECT 8.010 222.035 8.550 222.315 ;
        RECT 9.390 222.035 9.930 222.315 ;
        RECT 10.770 222.035 11.310 222.315 ;
        RECT 12.150 222.035 12.690 222.315 ;
        RECT 13.530 222.035 14.070 222.315 ;
        RECT 14.910 222.035 15.450 222.315 ;
        RECT 16.290 222.035 16.830 222.315 ;
        RECT 17.670 222.035 18.210 222.315 ;
        RECT 19.050 222.035 19.590 222.315 ;
        RECT 20.430 222.035 20.970 222.315 ;
        RECT 21.810 222.035 22.350 222.315 ;
        RECT 23.190 222.035 23.730 222.315 ;
        RECT 24.570 222.035 25.110 222.315 ;
        RECT 25.950 222.035 26.490 222.315 ;
        RECT 27.330 222.035 27.870 222.315 ;
        RECT 28.710 222.035 29.250 222.315 ;
        RECT 30.090 222.035 30.630 222.315 ;
        RECT 31.470 222.035 32.010 222.315 ;
        RECT 32.850 222.035 33.850 222.315 ;
        RECT 34.690 222.035 35.230 222.315 ;
        RECT 36.070 222.035 36.610 222.315 ;
        RECT 37.450 222.035 37.990 222.315 ;
        RECT 38.830 222.035 39.370 222.315 ;
        RECT 40.210 222.035 40.750 222.315 ;
        RECT 41.590 222.035 42.130 222.315 ;
        RECT 42.970 222.035 43.510 222.315 ;
        RECT 44.350 222.035 44.890 222.315 ;
        RECT 45.730 222.035 46.270 222.315 ;
        RECT 47.110 222.035 47.650 222.315 ;
        RECT 48.490 222.035 49.030 222.315 ;
        RECT 49.870 222.035 50.410 222.315 ;
        RECT 51.250 222.035 51.790 222.315 ;
        RECT 52.630 222.035 53.170 222.315 ;
        RECT 54.010 222.035 54.550 222.315 ;
        RECT 55.390 222.035 55.930 222.315 ;
        RECT 56.770 222.035 57.310 222.315 ;
        RECT 58.150 222.035 58.690 222.315 ;
        RECT 59.530 222.035 60.070 222.315 ;
        RECT 60.910 222.035 61.450 222.315 ;
        RECT 62.290 222.035 62.830 222.315 ;
        RECT 63.670 222.035 64.210 222.315 ;
        RECT 65.050 222.035 66.050 222.315 ;
        RECT 66.890 222.035 67.430 222.315 ;
        RECT 68.270 222.035 68.810 222.315 ;
        RECT 69.650 222.035 70.190 222.315 ;
        RECT 71.030 222.035 71.570 222.315 ;
        RECT 72.410 222.035 72.950 222.315 ;
        RECT 73.790 222.035 74.330 222.315 ;
        RECT 75.170 222.035 75.710 222.315 ;
        RECT 76.550 222.035 77.090 222.315 ;
        RECT 77.930 222.035 78.470 222.315 ;
        RECT 79.310 222.035 79.850 222.315 ;
        RECT 80.690 222.035 81.230 222.315 ;
        RECT 82.070 222.035 82.610 222.315 ;
        RECT 83.450 222.035 83.990 222.315 ;
        RECT 84.830 222.035 85.370 222.315 ;
        RECT 86.210 222.035 86.750 222.315 ;
        RECT 87.590 222.035 88.130 222.315 ;
        RECT 88.970 222.035 89.510 222.315 ;
        RECT 90.350 222.035 90.890 222.315 ;
        RECT 91.730 222.035 92.270 222.315 ;
        RECT 93.110 222.035 93.650 222.315 ;
        RECT 94.490 222.035 95.030 222.315 ;
        RECT 95.870 222.035 96.410 222.315 ;
        RECT 97.250 222.035 98.250 222.315 ;
        RECT 99.090 222.035 99.630 222.315 ;
        RECT 100.470 222.035 101.010 222.315 ;
        RECT 101.850 222.035 102.390 222.315 ;
        RECT 103.230 222.035 103.770 222.315 ;
        RECT 104.610 222.035 105.150 222.315 ;
        RECT 105.990 222.035 106.530 222.315 ;
        RECT 107.370 222.035 107.910 222.315 ;
        RECT 108.750 222.035 109.290 222.315 ;
        RECT 110.130 222.035 110.670 222.315 ;
        RECT 111.510 222.035 112.050 222.315 ;
        RECT 112.890 222.035 113.430 222.315 ;
        RECT 114.270 222.035 114.810 222.315 ;
        RECT 115.650 222.035 116.190 222.315 ;
        RECT 117.030 222.035 117.570 222.315 ;
        RECT 118.410 222.035 118.950 222.315 ;
        RECT 119.790 222.035 120.330 222.315 ;
        RECT 121.170 222.035 121.710 222.315 ;
        RECT 122.550 222.035 123.090 222.315 ;
        RECT 123.930 222.035 124.470 222.315 ;
        RECT 125.310 222.035 125.850 222.315 ;
        RECT 126.690 222.035 127.230 222.315 ;
        RECT 128.070 222.035 128.610 222.315 ;
        RECT 129.450 222.035 130.000 222.315 ;
        RECT 0.560 87.960 130.000 222.035 ;
        RECT 0.560 44.300 130.020 87.960 ;
        RECT 0.560 1.080 130.000 44.300 ;
        RECT 1.110 0.010 1.650 1.080 ;
        RECT 2.490 0.010 3.030 1.080 ;
        RECT 3.870 0.010 4.410 1.080 ;
        RECT 5.250 0.010 5.790 1.080 ;
        RECT 6.630 0.010 7.170 1.080 ;
        RECT 8.010 0.010 8.550 1.080 ;
        RECT 9.390 0.010 9.930 1.080 ;
        RECT 10.770 0.010 11.310 1.080 ;
        RECT 12.150 0.010 12.690 1.080 ;
        RECT 13.530 0.010 14.070 1.080 ;
        RECT 14.910 0.010 15.450 1.080 ;
        RECT 16.290 0.010 16.830 1.080 ;
        RECT 17.670 0.010 18.210 1.080 ;
        RECT 19.050 0.010 19.590 1.080 ;
        RECT 20.430 0.010 20.970 1.080 ;
        RECT 21.810 0.010 22.350 1.080 ;
        RECT 23.190 0.010 23.730 1.080 ;
        RECT 24.570 0.010 25.110 1.080 ;
        RECT 25.950 0.010 26.490 1.080 ;
        RECT 27.330 0.010 27.870 1.080 ;
        RECT 28.710 0.010 29.250 1.080 ;
        RECT 30.090 0.010 30.630 1.080 ;
        RECT 31.470 0.010 32.010 1.080 ;
        RECT 32.850 0.010 33.850 1.080 ;
        RECT 34.690 0.010 35.230 1.080 ;
        RECT 36.070 0.010 36.610 1.080 ;
        RECT 37.450 0.010 37.990 1.080 ;
        RECT 38.830 0.010 39.370 1.080 ;
        RECT 40.210 0.010 40.750 1.080 ;
        RECT 41.590 0.010 42.130 1.080 ;
        RECT 42.970 0.010 43.510 1.080 ;
        RECT 44.350 0.010 44.890 1.080 ;
        RECT 45.730 0.010 46.270 1.080 ;
        RECT 47.110 0.010 47.650 1.080 ;
        RECT 48.490 0.010 49.030 1.080 ;
        RECT 49.870 0.010 50.410 1.080 ;
        RECT 51.250 0.010 51.790 1.080 ;
        RECT 52.630 0.010 53.170 1.080 ;
        RECT 54.010 0.010 54.550 1.080 ;
        RECT 55.390 0.010 55.930 1.080 ;
        RECT 56.770 0.010 57.310 1.080 ;
        RECT 58.150 0.010 58.690 1.080 ;
        RECT 59.530 0.010 60.070 1.080 ;
        RECT 60.910 0.010 61.450 1.080 ;
        RECT 62.290 0.010 62.830 1.080 ;
        RECT 63.670 0.010 64.210 1.080 ;
        RECT 65.050 0.010 66.050 1.080 ;
        RECT 66.890 0.010 67.430 1.080 ;
        RECT 68.270 0.010 68.810 1.080 ;
        RECT 69.650 0.010 70.190 1.080 ;
        RECT 71.030 0.010 71.570 1.080 ;
        RECT 72.410 0.010 72.950 1.080 ;
        RECT 73.790 0.010 74.330 1.080 ;
        RECT 75.170 0.010 75.710 1.080 ;
        RECT 76.550 0.010 77.090 1.080 ;
        RECT 77.930 0.010 78.470 1.080 ;
        RECT 79.310 0.010 79.850 1.080 ;
        RECT 80.690 0.010 81.230 1.080 ;
        RECT 82.070 0.010 82.610 1.080 ;
        RECT 83.450 0.010 83.990 1.080 ;
        RECT 84.830 0.010 85.370 1.080 ;
        RECT 86.210 0.010 86.750 1.080 ;
        RECT 87.590 0.010 88.130 1.080 ;
        RECT 88.970 0.010 89.510 1.080 ;
        RECT 90.350 0.010 90.890 1.080 ;
        RECT 91.730 0.010 92.270 1.080 ;
        RECT 93.110 0.010 93.650 1.080 ;
        RECT 94.490 0.010 95.030 1.080 ;
        RECT 95.870 0.010 96.410 1.080 ;
        RECT 97.250 0.010 98.250 1.080 ;
        RECT 99.090 0.010 99.630 1.080 ;
        RECT 100.470 0.010 101.010 1.080 ;
        RECT 101.850 0.010 102.390 1.080 ;
        RECT 103.230 0.010 103.770 1.080 ;
        RECT 104.610 0.010 105.150 1.080 ;
        RECT 105.990 0.010 106.530 1.080 ;
        RECT 107.370 0.010 107.910 1.080 ;
        RECT 108.750 0.010 109.290 1.080 ;
        RECT 110.130 0.010 110.670 1.080 ;
        RECT 111.510 0.010 112.050 1.080 ;
        RECT 112.890 0.010 113.430 1.080 ;
        RECT 114.270 0.010 114.810 1.080 ;
        RECT 115.650 0.010 116.190 1.080 ;
        RECT 117.030 0.010 117.570 1.080 ;
        RECT 118.410 0.010 118.950 1.080 ;
        RECT 119.790 0.010 120.330 1.080 ;
        RECT 121.170 0.010 121.710 1.080 ;
        RECT 122.550 0.010 123.090 1.080 ;
        RECT 123.930 0.010 124.470 1.080 ;
        RECT 125.310 0.010 125.850 1.080 ;
        RECT 126.690 0.010 127.230 1.080 ;
        RECT 128.070 0.010 128.610 1.080 ;
        RECT 129.450 0.010 130.000 1.080 ;
      LAYER met3 ;
        RECT 1.200 222.040 129.655 222.185 ;
        RECT 1.200 221.320 128.800 222.040 ;
        RECT 0.800 220.680 128.800 221.320 ;
        RECT 1.200 220.640 128.800 220.680 ;
        RECT 1.200 219.320 129.655 220.640 ;
        RECT 1.200 217.920 128.800 219.320 ;
        RECT 0.800 217.280 129.655 217.920 ;
        RECT 1.200 216.600 129.655 217.280 ;
        RECT 1.200 215.200 128.800 216.600 ;
        RECT 1.200 214.520 129.655 215.200 ;
        RECT 0.800 213.880 129.655 214.520 ;
        RECT 1.200 212.480 128.800 213.880 ;
        RECT 1.200 211.160 129.655 212.480 ;
        RECT 1.200 211.120 128.800 211.160 ;
        RECT 0.800 210.480 128.800 211.120 ;
        RECT 1.200 209.760 128.800 210.480 ;
        RECT 1.200 209.080 129.655 209.760 ;
        RECT 0.800 208.440 129.655 209.080 ;
        RECT 1.200 207.040 128.800 208.440 ;
        RECT 1.200 205.720 129.655 207.040 ;
        RECT 1.200 205.680 128.800 205.720 ;
        RECT 0.800 205.040 128.800 205.680 ;
        RECT 1.200 204.320 128.800 205.040 ;
        RECT 1.200 203.000 129.655 204.320 ;
        RECT 1.200 202.280 128.800 203.000 ;
        RECT 0.800 201.640 128.800 202.280 ;
        RECT 1.200 201.600 128.800 201.640 ;
        RECT 1.200 200.280 129.655 201.600 ;
        RECT 1.200 198.880 128.800 200.280 ;
        RECT 0.800 198.240 129.655 198.880 ;
        RECT 1.200 197.560 129.655 198.240 ;
        RECT 1.200 196.160 128.800 197.560 ;
        RECT 1.200 195.480 129.655 196.160 ;
        RECT 0.800 194.840 129.655 195.480 ;
        RECT 1.200 194.160 129.655 194.840 ;
        RECT 1.200 193.440 128.800 194.160 ;
        RECT 0.800 192.800 128.800 193.440 ;
        RECT 1.200 192.760 128.800 192.800 ;
        RECT 1.200 191.440 129.655 192.760 ;
        RECT 1.200 190.040 128.800 191.440 ;
        RECT 0.800 189.400 129.655 190.040 ;
        RECT 1.200 188.720 129.655 189.400 ;
        RECT 1.200 187.320 128.800 188.720 ;
        RECT 1.200 186.640 129.655 187.320 ;
        RECT 0.800 186.000 129.655 186.640 ;
        RECT 1.200 184.600 128.800 186.000 ;
        RECT 1.200 183.280 129.655 184.600 ;
        RECT 1.200 183.240 128.800 183.280 ;
        RECT 0.800 182.600 128.800 183.240 ;
        RECT 1.200 181.880 128.800 182.600 ;
        RECT 1.200 181.200 129.655 181.880 ;
        RECT 0.800 180.560 129.655 181.200 ;
        RECT 1.200 179.160 128.800 180.560 ;
        RECT 1.200 177.840 129.655 179.160 ;
        RECT 1.200 177.800 128.800 177.840 ;
        RECT 0.800 177.160 128.800 177.800 ;
        RECT 1.200 176.440 128.800 177.160 ;
        RECT 1.200 175.120 129.655 176.440 ;
        RECT 1.200 174.400 128.800 175.120 ;
        RECT 0.800 173.760 128.800 174.400 ;
        RECT 1.200 173.720 128.800 173.760 ;
        RECT 1.200 172.400 129.655 173.720 ;
        RECT 1.200 171.000 128.800 172.400 ;
        RECT 0.800 170.360 129.655 171.000 ;
        RECT 1.200 169.680 129.655 170.360 ;
        RECT 1.200 168.280 128.800 169.680 ;
        RECT 1.200 167.600 129.655 168.280 ;
        RECT 0.800 166.960 129.655 167.600 ;
        RECT 1.200 166.280 129.655 166.960 ;
        RECT 1.200 165.560 128.800 166.280 ;
        RECT 0.800 164.920 128.800 165.560 ;
        RECT 1.200 164.880 128.800 164.920 ;
        RECT 1.200 163.560 129.655 164.880 ;
        RECT 1.200 162.160 128.800 163.560 ;
        RECT 0.800 161.520 129.655 162.160 ;
        RECT 1.200 160.840 129.655 161.520 ;
        RECT 1.200 159.440 128.800 160.840 ;
        RECT 1.200 158.760 129.655 159.440 ;
        RECT 0.800 158.120 129.655 158.760 ;
        RECT 1.200 156.720 128.800 158.120 ;
        RECT 1.200 155.400 129.655 156.720 ;
        RECT 1.200 155.360 128.800 155.400 ;
        RECT 0.800 154.720 128.800 155.360 ;
        RECT 1.200 154.000 128.800 154.720 ;
        RECT 1.200 153.320 129.655 154.000 ;
        RECT 0.800 152.680 129.655 153.320 ;
        RECT 1.200 151.280 128.800 152.680 ;
        RECT 1.200 149.960 129.655 151.280 ;
        RECT 1.200 149.920 128.800 149.960 ;
        RECT 0.800 149.280 128.800 149.920 ;
        RECT 1.200 148.560 128.800 149.280 ;
        RECT 1.200 147.240 129.655 148.560 ;
        RECT 1.200 146.520 128.800 147.240 ;
        RECT 0.800 145.880 128.800 146.520 ;
        RECT 1.200 145.840 128.800 145.880 ;
        RECT 1.200 144.520 129.655 145.840 ;
        RECT 1.200 143.120 128.800 144.520 ;
        RECT 0.800 142.480 129.655 143.120 ;
        RECT 1.200 141.800 129.655 142.480 ;
        RECT 1.200 140.400 128.800 141.800 ;
        RECT 1.200 139.720 129.655 140.400 ;
        RECT 0.800 139.080 129.655 139.720 ;
        RECT 1.200 138.400 129.655 139.080 ;
        RECT 1.200 137.680 128.800 138.400 ;
        RECT 0.800 137.040 128.800 137.680 ;
        RECT 1.200 137.000 128.800 137.040 ;
        RECT 1.200 135.680 129.655 137.000 ;
        RECT 1.200 134.280 128.800 135.680 ;
        RECT 0.800 133.640 129.655 134.280 ;
        RECT 1.200 132.960 129.655 133.640 ;
        RECT 1.200 131.560 128.800 132.960 ;
        RECT 1.200 130.880 129.655 131.560 ;
        RECT 0.800 130.240 129.655 130.880 ;
        RECT 1.200 128.840 128.800 130.240 ;
        RECT 1.200 127.520 129.655 128.840 ;
        RECT 1.200 127.480 128.800 127.520 ;
        RECT 0.800 126.840 128.800 127.480 ;
        RECT 1.200 126.120 128.800 126.840 ;
        RECT 1.200 125.440 129.655 126.120 ;
        RECT 0.800 124.800 129.655 125.440 ;
        RECT 1.200 123.400 128.800 124.800 ;
        RECT 1.200 122.080 129.655 123.400 ;
        RECT 1.200 122.040 128.800 122.080 ;
        RECT 0.800 121.400 128.800 122.040 ;
        RECT 1.200 120.680 128.800 121.400 ;
        RECT 1.200 119.360 129.655 120.680 ;
        RECT 1.200 118.640 128.800 119.360 ;
        RECT 0.800 118.000 128.800 118.640 ;
        RECT 1.200 117.960 128.800 118.000 ;
        RECT 1.200 116.640 129.655 117.960 ;
        RECT 1.200 115.240 128.800 116.640 ;
        RECT 0.800 114.600 129.655 115.240 ;
        RECT 1.200 113.920 129.655 114.600 ;
        RECT 1.200 112.520 128.800 113.920 ;
        RECT 1.200 111.840 129.655 112.520 ;
        RECT 0.800 111.200 129.655 111.840 ;
        RECT 1.200 110.520 129.655 111.200 ;
        RECT 1.200 109.800 128.800 110.520 ;
        RECT 0.800 109.160 128.800 109.800 ;
        RECT 1.200 109.120 128.800 109.160 ;
        RECT 1.200 107.800 129.655 109.120 ;
        RECT 1.200 106.400 128.800 107.800 ;
        RECT 0.800 105.760 129.655 106.400 ;
        RECT 1.200 105.080 129.655 105.760 ;
        RECT 1.200 103.680 128.800 105.080 ;
        RECT 1.200 103.000 129.655 103.680 ;
        RECT 0.800 102.360 129.655 103.000 ;
        RECT 1.200 100.960 128.800 102.360 ;
        RECT 1.200 99.640 129.655 100.960 ;
        RECT 1.200 99.600 128.800 99.640 ;
        RECT 0.800 98.960 128.800 99.600 ;
        RECT 1.200 98.240 128.800 98.960 ;
        RECT 1.200 97.560 129.655 98.240 ;
        RECT 0.800 96.920 129.655 97.560 ;
        RECT 1.200 95.520 128.800 96.920 ;
        RECT 1.200 94.200 129.655 95.520 ;
        RECT 1.200 94.160 128.800 94.200 ;
        RECT 0.800 93.520 128.800 94.160 ;
        RECT 1.200 92.800 128.800 93.520 ;
        RECT 1.200 91.480 129.655 92.800 ;
        RECT 1.200 90.760 128.800 91.480 ;
        RECT 0.800 90.120 128.800 90.760 ;
        RECT 1.200 90.080 128.800 90.120 ;
        RECT 1.200 88.760 129.655 90.080 ;
        RECT 1.200 87.360 128.800 88.760 ;
        RECT 0.800 86.720 129.655 87.360 ;
        RECT 1.200 86.040 129.655 86.720 ;
        RECT 1.200 84.640 128.800 86.040 ;
        RECT 1.200 83.960 129.655 84.640 ;
        RECT 0.800 83.320 129.655 83.960 ;
        RECT 1.200 82.640 129.655 83.320 ;
        RECT 1.200 81.920 128.800 82.640 ;
        RECT 0.800 81.280 128.800 81.920 ;
        RECT 1.200 81.240 128.800 81.280 ;
        RECT 1.200 79.920 129.655 81.240 ;
        RECT 1.200 78.520 128.800 79.920 ;
        RECT 0.800 77.880 129.655 78.520 ;
        RECT 1.200 77.200 129.655 77.880 ;
        RECT 1.200 75.800 128.800 77.200 ;
        RECT 1.200 75.120 129.655 75.800 ;
        RECT 0.800 74.480 129.655 75.120 ;
        RECT 1.200 73.080 128.800 74.480 ;
        RECT 1.200 71.760 129.655 73.080 ;
        RECT 1.200 71.720 128.800 71.760 ;
        RECT 0.800 71.080 128.800 71.720 ;
        RECT 1.200 70.360 128.800 71.080 ;
        RECT 1.200 69.680 129.655 70.360 ;
        RECT 0.800 69.040 129.655 69.680 ;
        RECT 1.200 67.640 128.800 69.040 ;
        RECT 1.200 66.320 129.655 67.640 ;
        RECT 1.200 66.280 128.800 66.320 ;
        RECT 0.800 65.640 128.800 66.280 ;
        RECT 1.200 64.920 128.800 65.640 ;
        RECT 1.200 63.600 129.655 64.920 ;
        RECT 1.200 62.880 128.800 63.600 ;
        RECT 0.800 62.240 128.800 62.880 ;
        RECT 1.200 62.200 128.800 62.240 ;
        RECT 1.200 60.880 129.655 62.200 ;
        RECT 1.200 59.480 128.800 60.880 ;
        RECT 0.800 58.840 129.655 59.480 ;
        RECT 1.200 58.160 129.655 58.840 ;
        RECT 1.200 56.760 128.800 58.160 ;
        RECT 1.200 56.080 129.655 56.760 ;
        RECT 0.800 55.440 129.655 56.080 ;
        RECT 1.200 54.760 129.655 55.440 ;
        RECT 1.200 54.040 128.800 54.760 ;
        RECT 0.800 53.400 128.800 54.040 ;
        RECT 1.200 53.360 128.800 53.400 ;
        RECT 1.200 52.040 129.655 53.360 ;
        RECT 1.200 50.640 128.800 52.040 ;
        RECT 0.800 50.000 129.655 50.640 ;
        RECT 1.200 49.320 129.655 50.000 ;
        RECT 1.200 47.920 128.800 49.320 ;
        RECT 1.200 47.240 129.655 47.920 ;
        RECT 0.800 46.600 129.655 47.240 ;
        RECT 1.200 45.200 128.800 46.600 ;
        RECT 1.200 43.880 129.655 45.200 ;
        RECT 1.200 43.840 128.800 43.880 ;
        RECT 0.800 43.200 128.800 43.840 ;
        RECT 1.200 42.480 128.800 43.200 ;
        RECT 1.200 41.800 129.655 42.480 ;
        RECT 0.800 41.160 129.655 41.800 ;
        RECT 1.200 39.760 128.800 41.160 ;
        RECT 1.200 38.440 129.655 39.760 ;
        RECT 1.200 38.400 128.800 38.440 ;
        RECT 0.800 37.760 128.800 38.400 ;
        RECT 1.200 37.040 128.800 37.760 ;
        RECT 1.200 35.720 129.655 37.040 ;
        RECT 1.200 35.000 128.800 35.720 ;
        RECT 0.800 34.360 128.800 35.000 ;
        RECT 1.200 34.320 128.800 34.360 ;
        RECT 1.200 33.000 129.655 34.320 ;
        RECT 1.200 31.600 128.800 33.000 ;
        RECT 0.800 30.960 129.655 31.600 ;
        RECT 1.200 30.280 129.655 30.960 ;
        RECT 1.200 28.880 128.800 30.280 ;
        RECT 1.200 28.200 129.655 28.880 ;
        RECT 0.800 27.560 129.655 28.200 ;
        RECT 1.200 26.880 129.655 27.560 ;
        RECT 1.200 26.160 128.800 26.880 ;
        RECT 0.800 25.520 128.800 26.160 ;
        RECT 1.200 25.480 128.800 25.520 ;
        RECT 1.200 24.160 129.655 25.480 ;
        RECT 1.200 22.760 128.800 24.160 ;
        RECT 0.800 22.120 129.655 22.760 ;
        RECT 1.200 21.440 129.655 22.120 ;
        RECT 1.200 20.040 128.800 21.440 ;
        RECT 1.200 19.360 129.655 20.040 ;
        RECT 0.800 18.720 129.655 19.360 ;
        RECT 1.200 17.320 128.800 18.720 ;
        RECT 1.200 16.000 129.655 17.320 ;
        RECT 1.200 15.960 128.800 16.000 ;
        RECT 0.800 15.320 128.800 15.960 ;
        RECT 1.200 14.600 128.800 15.320 ;
        RECT 1.200 13.920 129.655 14.600 ;
        RECT 0.800 13.280 129.655 13.920 ;
        RECT 1.200 11.880 128.800 13.280 ;
        RECT 1.200 10.560 129.655 11.880 ;
        RECT 1.200 10.520 128.800 10.560 ;
        RECT 0.800 9.880 128.800 10.520 ;
        RECT 1.200 9.160 128.800 9.880 ;
        RECT 1.200 7.840 129.655 9.160 ;
        RECT 1.200 7.120 128.800 7.840 ;
        RECT 0.800 6.480 128.800 7.120 ;
        RECT 1.200 6.440 128.800 6.480 ;
        RECT 1.200 5.120 129.655 6.440 ;
        RECT 1.200 3.720 128.800 5.120 ;
        RECT 0.800 3.080 129.655 3.720 ;
        RECT 1.200 2.400 129.655 3.080 ;
        RECT 1.200 1.000 128.800 2.400 ;
        RECT 1.200 0.855 129.655 1.000 ;
      LAYER met4 ;
        RECT 4.895 218.240 114.705 220.145 ;
        RECT 4.895 4.800 24.145 218.240 ;
        RECT 26.545 4.800 43.970 218.240 ;
        RECT 46.370 4.800 63.795 218.240 ;
        RECT 66.195 4.800 83.625 218.240 ;
        RECT 86.025 4.800 103.450 218.240 ;
        RECT 105.850 4.800 114.705 218.240 ;
        RECT 4.895 3.575 114.705 4.800 ;
  END
END RAM_IO
END LIBRARY

