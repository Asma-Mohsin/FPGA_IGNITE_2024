VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM_IO
  CLASS BLOCK ;
  FOREIGN RAM_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 181.000 BY 231.000 ;
  PIN Config_accessC_bit0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 217.750 181.000 218.130 ;
    END
  END Config_accessC_bit0
  PIN Config_accessC_bit1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 220.470 181.000 220.850 ;
    END
  END Config_accessC_bit1
  PIN Config_accessC_bit2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 223.190 181.000 223.570 ;
    END
  END Config_accessC_bit2
  PIN Config_accessC_bit3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 225.910 181.000 226.290 ;
    END
  END Config_accessC_bit3
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.550 0.700 3.930 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.590 0.700 5.970 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.950 0.700 7.330 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.990 0.700 9.370 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.630 0.700 25.010 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.990 0.700 26.370 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.030 0.700 28.410 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.390 0.700 29.770 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.430 0.700 31.810 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.470 0.700 33.850 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.830 0.700 35.210 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.870 0.700 37.250 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.350 0.700 10.730 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.390 0.700 12.770 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.750 0.700 14.130 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.790 0.700 16.170 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.150 0.700 17.530 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.190 0.700 19.570 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.230 0.700 21.610 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.590 0.700 22.970 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.110 0.700 66.490 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.790 0.700 84.170 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.150 0.700 85.530 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.150 0.700 68.530 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.510 0.700 69.890 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.550 0.700 71.930 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.910 0.700 73.290 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.950 0.700 75.330 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.310 0.700 76.690 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.350 0.700 78.730 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.390 0.700 80.770 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.750 0.700 82.130 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.230 0.700 38.610 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.910 0.700 56.290 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.270 0.700 57.650 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.310 0.700 59.690 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.670 0.700 61.050 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.710 0.700 63.090 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.750 0.700 65.130 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.270 0.700 40.650 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.630 0.700 42.010 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.670 0.700 44.050 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.030 0.700 45.410 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.070 0.700 47.450 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.110 0.700 49.490 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.470 0.700 50.850 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.510 0.700 52.890 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.870 0.700 54.250 ;
    END
  END EE4END[9]
  PIN FAB2RAM_A0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 183.750 181.000 184.130 ;
    END
  END FAB2RAM_A0_O0
  PIN FAB2RAM_A0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 186.470 181.000 186.850 ;
    END
  END FAB2RAM_A0_O1
  PIN FAB2RAM_A0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 189.190 181.000 189.570 ;
    END
  END FAB2RAM_A0_O2
  PIN FAB2RAM_A0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 191.910 181.000 192.290 ;
    END
  END FAB2RAM_A0_O3
  PIN FAB2RAM_A1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 195.310 181.000 195.690 ;
    END
  END FAB2RAM_A1_O0
  PIN FAB2RAM_A1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 198.030 181.000 198.410 ;
    END
  END FAB2RAM_A1_O1
  PIN FAB2RAM_A1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 200.750 181.000 201.130 ;
    END
  END FAB2RAM_A1_O2
  PIN FAB2RAM_A1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 203.470 181.000 203.850 ;
    END
  END FAB2RAM_A1_O3
  PIN FAB2RAM_C_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 206.190 181.000 206.570 ;
    END
  END FAB2RAM_C_O0
  PIN FAB2RAM_C_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 208.910 181.000 209.290 ;
    END
  END FAB2RAM_C_O1
  PIN FAB2RAM_C_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 211.630 181.000 212.010 ;
    END
  END FAB2RAM_C_O2
  PIN FAB2RAM_C_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 214.350 181.000 214.730 ;
    END
  END FAB2RAM_C_O3
  PIN FAB2RAM_D0_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 138.870 181.000 139.250 ;
    END
  END FAB2RAM_D0_O0
  PIN FAB2RAM_D0_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 141.590 181.000 141.970 ;
    END
  END FAB2RAM_D0_O1
  PIN FAB2RAM_D0_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 144.310 181.000 144.690 ;
    END
  END FAB2RAM_D0_O2
  PIN FAB2RAM_D0_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 147.710 181.000 148.090 ;
    END
  END FAB2RAM_D0_O3
  PIN FAB2RAM_D1_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 150.430 181.000 150.810 ;
    END
  END FAB2RAM_D1_O0
  PIN FAB2RAM_D1_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 153.150 181.000 153.530 ;
    END
  END FAB2RAM_D1_O1
  PIN FAB2RAM_D1_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 155.870 181.000 156.250 ;
    END
  END FAB2RAM_D1_O2
  PIN FAB2RAM_D1_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 158.590 181.000 158.970 ;
    END
  END FAB2RAM_D1_O3
  PIN FAB2RAM_D2_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 161.310 181.000 161.690 ;
    END
  END FAB2RAM_D2_O0
  PIN FAB2RAM_D2_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 164.030 181.000 164.410 ;
    END
  END FAB2RAM_D2_O1
  PIN FAB2RAM_D2_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 166.750 181.000 167.130 ;
    END
  END FAB2RAM_D2_O2
  PIN FAB2RAM_D2_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 170.150 181.000 170.530 ;
    END
  END FAB2RAM_D2_O3
  PIN FAB2RAM_D3_O0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 172.870 181.000 173.250 ;
    END
  END FAB2RAM_D3_O0
  PIN FAB2RAM_D3_O1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 175.590 181.000 175.970 ;
    END
  END FAB2RAM_D3_O1
  PIN FAB2RAM_D3_O2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 178.310 181.000 178.690 ;
    END
  END FAB2RAM_D3_O2
  PIN FAB2RAM_D3_O3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 181.030 181.000 181.410 ;
    END
  END FAB2RAM_D3_O3
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.830 0.700 171.210 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.830 0.700 188.210 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.870 0.700 190.250 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.230 0.700 191.610 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.270 0.700 193.650 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.630 0.700 195.010 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.670 0.700 197.050 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.710 0.700 199.090 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.070 0.700 200.450 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.110 0.700 202.490 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.470 0.700 203.850 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.190 0.700 172.570 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.510 0.700 205.890 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.870 0.700 207.250 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.910 0.700 209.290 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.950 0.700 211.330 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.310 0.700 212.690 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.350 0.700 214.730 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.710 0.700 216.090 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.750 0.700 218.130 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.110 0.700 219.490 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.150 0.700 221.530 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.230 0.700 174.610 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.510 0.700 222.890 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.550 0.700 224.930 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.590 0.700 175.970 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.630 0.700 178.010 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.990 0.700 179.370 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.030 0.700 181.410 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.070 0.700 183.450 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.430 0.700 184.810 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.470 0.700 186.850 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 4.910 181.000 5.290 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 32.790 181.000 33.170 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 35.510 181.000 35.890 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 38.230 181.000 38.610 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 40.950 181.000 41.330 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 43.670 181.000 44.050 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 46.390 181.000 46.770 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 49.110 181.000 49.490 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 52.510 181.000 52.890 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 55.230 181.000 55.610 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 57.950 181.000 58.330 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 7.630 181.000 8.010 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 60.670 181.000 61.050 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 63.390 181.000 63.770 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 66.110 181.000 66.490 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 68.830 181.000 69.210 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 71.550 181.000 71.930 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 74.950 181.000 75.330 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 77.670 181.000 78.050 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 80.390 181.000 80.770 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 83.110 181.000 83.490 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 85.830 181.000 86.210 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 10.350 181.000 10.730 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 88.550 181.000 88.930 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 91.270 181.000 91.650 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 13.070 181.000 13.450 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 15.790 181.000 16.170 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 18.510 181.000 18.890 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 21.230 181.000 21.610 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 23.950 181.000 24.330 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 27.350 181.000 27.730 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 30.070 181.000 30.450 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 138.960 0.000 139.340 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 157.820 0.000 158.200 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 159.660 0.000 160.040 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 161.500 0.000 161.880 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 163.340 0.000 163.720 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 165.180 0.000 165.560 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 167.480 0.000 167.860 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.320 0.000 169.700 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 171.160 0.000 171.540 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.000 0.000 173.380 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 174.840 0.000 175.220 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 140.800 0.000 141.180 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 142.640 0.000 143.020 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.480 0.000 144.860 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 146.780 0.000 147.160 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 148.620 0.000 149.000 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 150.460 0.000 150.840 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 152.300 0.000 152.680 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 154.140 0.000 154.520 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 155.980 0.000 156.360 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.960 230.300 139.340 231.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 157.820 230.300 158.200 231.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 159.660 230.300 160.040 231.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.500 230.300 161.880 231.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 163.340 230.300 163.720 231.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.180 230.300 165.560 231.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.480 230.300 167.860 231.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 169.320 230.300 169.700 231.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 171.160 230.300 171.540 231.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.000 230.300 173.380 231.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 174.840 230.300 175.220 231.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.800 230.300 141.180 231.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.640 230.300 143.020 231.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.480 230.300 144.860 231.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.780 230.300 147.160 231.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.620 230.300 149.000 231.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.460 230.300 150.840 231.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.300 230.300 152.680 231.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.140 230.300 154.520 231.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.980 230.300 156.360 231.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 3.720 230.300 4.100 231.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 5.560 230.300 5.940 231.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 7.400 230.300 7.780 231.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.240 230.300 9.620 231.000 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 3.720 0.000 4.100 0.700 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 5.560 0.000 5.940 0.700 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 7.400 0.000 7.780 0.700 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 9.240 0.000 9.620 0.700 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 11.080 230.300 11.460 231.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 12.920 230.300 13.300 231.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 14.760 230.300 15.140 231.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.060 230.300 17.440 231.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 18.900 230.300 19.280 231.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 20.740 230.300 21.120 231.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.580 230.300 22.960 231.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.420 230.300 24.800 231.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 26.260 230.300 26.640 231.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 28.100 230.300 28.480 231.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.940 230.300 30.320 231.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 31.780 230.300 32.160 231.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.620 230.300 34.000 231.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.460 230.300 35.840 231.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 37.760 230.300 38.140 231.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 39.600 230.300 39.980 231.000 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 26.260 0.000 26.640 0.700 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 28.100 0.000 28.480 0.700 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.940 0.000 30.320 0.700 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 31.780 0.000 32.160 0.700 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 33.620 0.000 34.000 0.700 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.460 0.000 35.840 0.700 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 37.760 0.000 38.140 0.700 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 39.600 0.000 39.980 0.700 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 11.080 0.000 11.460 0.700 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.920 0.000 13.300 0.700 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 14.760 0.000 15.140 0.700 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 17.060 0.000 17.440 0.700 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 18.900 0.000 19.280 0.700 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 20.740 0.000 21.120 0.700 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 22.580 0.000 22.960 0.700 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 24.420 0.000 24.800 0.700 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.440 230.300 41.820 231.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 60.300 230.300 60.680 231.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 62.140 230.300 62.520 231.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 63.980 230.300 64.360 231.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.820 230.300 66.200 231.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.660 230.300 68.040 231.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.500 230.300 69.880 231.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 43.280 230.300 43.660 231.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.120 230.300 45.500 231.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.960 230.300 47.340 231.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.800 230.300 49.180 231.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 50.640 230.300 51.020 231.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.480 230.300 52.860 231.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.320 230.300 54.700 231.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 56.160 230.300 56.540 231.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 230.300 58.380 231.000 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.440 0.000 41.820 0.700 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 60.300 0.000 60.680 0.700 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 62.140 0.000 62.520 0.700 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 63.980 0.000 64.360 0.700 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 65.820 0.000 66.200 0.700 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.660 0.000 68.040 0.700 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 69.500 0.000 69.880 0.700 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 43.280 0.000 43.660 0.700 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 45.120 0.000 45.500 0.700 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 46.960 0.000 47.340 0.700 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.800 0.000 49.180 0.700 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 50.640 0.000 51.020 0.700 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 52.480 0.000 52.860 0.700 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.320 0.000 54.700 0.700 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.160 0.000 56.540 0.700 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 58.000 0.000 58.380 0.700 ;
    END
  END N4END[9]
  PIN RAM2FAB_D0_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 93.990 181.000 94.370 ;
    END
  END RAM2FAB_D0_I0
  PIN RAM2FAB_D0_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 96.710 181.000 97.090 ;
    END
  END RAM2FAB_D0_I1
  PIN RAM2FAB_D0_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 100.110 181.000 100.490 ;
    END
  END RAM2FAB_D0_I2
  PIN RAM2FAB_D0_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 102.830 181.000 103.210 ;
    END
  END RAM2FAB_D0_I3
  PIN RAM2FAB_D1_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 105.550 181.000 105.930 ;
    END
  END RAM2FAB_D1_I0
  PIN RAM2FAB_D1_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 108.270 181.000 108.650 ;
    END
  END RAM2FAB_D1_I1
  PIN RAM2FAB_D1_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 110.990 181.000 111.370 ;
    END
  END RAM2FAB_D1_I2
  PIN RAM2FAB_D1_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 113.710 181.000 114.090 ;
    END
  END RAM2FAB_D1_I3
  PIN RAM2FAB_D2_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 180.300 116.430 181.000 116.810 ;
    END
  END RAM2FAB_D2_I0
  PIN RAM2FAB_D2_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 119.150 181.000 119.530 ;
    END
  END RAM2FAB_D2_I1
  PIN RAM2FAB_D2_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 122.550 181.000 122.930 ;
    END
  END RAM2FAB_D2_I2
  PIN RAM2FAB_D2_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 125.270 181.000 125.650 ;
    END
  END RAM2FAB_D2_I3
  PIN RAM2FAB_D3_I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 127.990 181.000 128.370 ;
    END
  END RAM2FAB_D3_I0
  PIN RAM2FAB_D3_I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 130.710 181.000 131.090 ;
    END
  END RAM2FAB_D3_I1
  PIN RAM2FAB_D3_I2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 180.300 133.430 181.000 133.810 ;
    END
  END RAM2FAB_D3_I2
  PIN RAM2FAB_D3_I3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 180.300 136.150 181.000 136.530 ;
    END
  END RAM2FAB_D3_I3
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 71.340 0.000 71.720 0.700 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.180 0.000 73.560 0.700 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 75.020 0.000 75.400 0.700 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 76.860 0.000 77.240 0.700 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 71.340 230.300 71.720 231.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 73.180 230.300 73.560 231.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 75.020 230.300 75.400 231.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 76.860 230.300 77.240 231.000 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.700 0.000 79.080 0.700 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 81.000 0.000 81.380 0.700 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.840 0.000 83.220 0.700 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 84.680 0.000 85.060 0.700 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 0.000 86.900 0.700 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 88.360 0.000 88.740 0.700 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.200 0.000 90.580 0.700 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.040 0.000 92.420 0.700 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.880 0.000 94.260 0.700 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 95.720 0.000 96.100 0.700 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 97.560 0.000 97.940 0.700 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.400 0.000 99.780 0.700 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.240 0.000 101.620 0.700 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.540 0.000 103.920 0.700 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.380 0.000 105.760 0.700 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.220 0.000 107.600 0.700 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 93.880 230.300 94.260 231.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 95.720 230.300 96.100 231.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 97.560 230.300 97.940 231.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.400 230.300 99.780 231.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 101.240 230.300 101.620 231.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 103.540 230.300 103.920 231.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 105.380 230.300 105.760 231.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 107.220 230.300 107.600 231.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 78.700 230.300 79.080 231.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 81.000 230.300 81.380 231.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.840 230.300 83.220 231.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 84.680 230.300 85.060 231.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 230.300 86.900 231.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 88.360 230.300 88.740 231.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 90.200 230.300 90.580 231.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 92.040 230.300 92.420 231.000 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.060 0.000 109.440 0.700 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.920 0.000 128.300 0.700 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 129.760 0.000 130.140 0.700 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 131.600 0.000 131.980 0.700 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 133.440 0.000 133.820 0.700 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.280 0.000 135.660 0.700 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 137.120 0.000 137.500 0.700 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.900 0.000 111.280 0.700 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.740 0.000 113.120 0.700 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.580 0.000 114.960 0.700 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.420 0.000 116.800 0.700 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.260 0.000 118.640 0.700 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 120.100 0.000 120.480 0.700 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.940 0.000 122.320 0.700 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.240 0.000 124.620 0.700 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 126.080 0.000 126.460 0.700 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.060 230.300 109.440 231.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.920 230.300 128.300 231.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 129.760 230.300 130.140 231.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 131.600 230.300 131.980 231.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 133.440 230.300 133.820 231.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 135.280 230.300 135.660 231.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 137.120 230.300 137.500 231.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.900 230.300 111.280 231.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 112.740 230.300 113.120 231.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 114.580 230.300 114.960 231.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 116.420 230.300 116.800 231.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 118.260 230.300 118.640 231.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 120.100 230.300 120.480 231.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 121.940 230.300 122.320 231.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.240 230.300 124.620 231.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 126.080 230.300 126.460 231.000 ;
    END
  END S4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 176.680 0.000 177.060 0.700 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 176.680 230.300 177.060 231.000 ;
    END
  END UserCLKo
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.190 0.700 87.570 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.550 0.700 88.930 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.590 0.700 90.970 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.630 0.700 93.010 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.990 0.700 94.370 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.030 0.700 96.410 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.390 0.700 97.770 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.430 0.700 99.810 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.790 0.700 101.170 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.830 0.700 103.210 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.190 0.700 104.570 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.230 0.700 106.610 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.270 0.700 108.650 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.630 0.700 110.010 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.670 0.700 112.050 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.030 0.700 113.410 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.070 0.700 115.450 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.430 0.700 116.810 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.470 0.700 118.850 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.830 0.700 120.210 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.750 0.700 150.130 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.430 0.700 167.810 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.790 0.700 169.170 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.790 0.700 152.170 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.150 0.700 153.530 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.190 0.700 155.570 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.550 0.700 156.930 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.590 0.700 158.970 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.950 0.700 160.330 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.990 0.700 162.370 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.350 0.700 163.730 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.390 0.700 165.770 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.870 0.700 122.250 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.550 0.700 139.930 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.910 0.700 141.290 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.950 0.700 143.330 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.310 0.700 144.690 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.350 0.700 146.730 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.710 0.700 148.090 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.910 0.700 124.290 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.270 0.700 125.650 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.310 0.700 127.690 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.670 0.700 129.050 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.710 0.700 131.090 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.070 0.700 132.450 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.110 0.700 134.490 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.470 0.700 135.850 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.510 0.700 137.890 ;
    END
  END WW4BEG[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -12.040 -11.660 -8.940 242.860 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 -11.660 192.820 -8.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 239.760 192.820 242.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.720 -11.660 192.820 242.860 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.580 -16.460 22.180 247.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 -16.460 175.780 247.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 21.290 197.620 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 174.470 197.620 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.840 -16.460 -13.740 247.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 -16.460 197.620 -13.360 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 244.560 197.620 247.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 194.520 -16.460 197.620 247.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.880 -16.460 25.480 247.660 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 24.590 197.620 26.190 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 177.770 197.620 179.370 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 4.870 5.355 175.910 225.950 ;
      LAYER li1 ;
        RECT 5.060 5.355 175.720 225.845 ;
      LAYER met1 ;
        RECT 1.450 1.740 180.250 229.800 ;
      LAYER met2 ;
        RECT 1.470 230.020 3.440 230.300 ;
        RECT 4.380 230.020 5.280 230.300 ;
        RECT 6.220 230.020 7.120 230.300 ;
        RECT 8.060 230.020 8.960 230.300 ;
        RECT 9.900 230.020 10.800 230.300 ;
        RECT 11.740 230.020 12.640 230.300 ;
        RECT 13.580 230.020 14.480 230.300 ;
        RECT 15.420 230.020 16.780 230.300 ;
        RECT 17.720 230.020 18.620 230.300 ;
        RECT 19.560 230.020 20.460 230.300 ;
        RECT 21.400 230.020 22.300 230.300 ;
        RECT 23.240 230.020 24.140 230.300 ;
        RECT 25.080 230.020 25.980 230.300 ;
        RECT 26.920 230.020 27.820 230.300 ;
        RECT 28.760 230.020 29.660 230.300 ;
        RECT 30.600 230.020 31.500 230.300 ;
        RECT 32.440 230.020 33.340 230.300 ;
        RECT 34.280 230.020 35.180 230.300 ;
        RECT 36.120 230.020 37.480 230.300 ;
        RECT 38.420 230.020 39.320 230.300 ;
        RECT 40.260 230.020 41.160 230.300 ;
        RECT 42.100 230.020 43.000 230.300 ;
        RECT 43.940 230.020 44.840 230.300 ;
        RECT 45.780 230.020 46.680 230.300 ;
        RECT 47.620 230.020 48.520 230.300 ;
        RECT 49.460 230.020 50.360 230.300 ;
        RECT 51.300 230.020 52.200 230.300 ;
        RECT 53.140 230.020 54.040 230.300 ;
        RECT 54.980 230.020 55.880 230.300 ;
        RECT 56.820 230.020 57.720 230.300 ;
        RECT 58.660 230.020 60.020 230.300 ;
        RECT 60.960 230.020 61.860 230.300 ;
        RECT 62.800 230.020 63.700 230.300 ;
        RECT 64.640 230.020 65.540 230.300 ;
        RECT 66.480 230.020 67.380 230.300 ;
        RECT 68.320 230.020 69.220 230.300 ;
        RECT 70.160 230.020 71.060 230.300 ;
        RECT 72.000 230.020 72.900 230.300 ;
        RECT 73.840 230.020 74.740 230.300 ;
        RECT 75.680 230.020 76.580 230.300 ;
        RECT 77.520 230.020 78.420 230.300 ;
        RECT 79.360 230.020 80.720 230.300 ;
        RECT 81.660 230.020 82.560 230.300 ;
        RECT 83.500 230.020 84.400 230.300 ;
        RECT 85.340 230.020 86.240 230.300 ;
        RECT 87.180 230.020 88.080 230.300 ;
        RECT 89.020 230.020 89.920 230.300 ;
        RECT 90.860 230.020 91.760 230.300 ;
        RECT 92.700 230.020 93.600 230.300 ;
        RECT 94.540 230.020 95.440 230.300 ;
        RECT 96.380 230.020 97.280 230.300 ;
        RECT 98.220 230.020 99.120 230.300 ;
        RECT 100.060 230.020 100.960 230.300 ;
        RECT 101.900 230.020 103.260 230.300 ;
        RECT 104.200 230.020 105.100 230.300 ;
        RECT 106.040 230.020 106.940 230.300 ;
        RECT 107.880 230.020 108.780 230.300 ;
        RECT 109.720 230.020 110.620 230.300 ;
        RECT 111.560 230.020 112.460 230.300 ;
        RECT 113.400 230.020 114.300 230.300 ;
        RECT 115.240 230.020 116.140 230.300 ;
        RECT 117.080 230.020 117.980 230.300 ;
        RECT 118.920 230.020 119.820 230.300 ;
        RECT 120.760 230.020 121.660 230.300 ;
        RECT 122.600 230.020 123.960 230.300 ;
        RECT 124.900 230.020 125.800 230.300 ;
        RECT 126.740 230.020 127.640 230.300 ;
        RECT 128.580 230.020 129.480 230.300 ;
        RECT 130.420 230.020 131.320 230.300 ;
        RECT 132.260 230.020 133.160 230.300 ;
        RECT 134.100 230.020 135.000 230.300 ;
        RECT 135.940 230.020 136.840 230.300 ;
        RECT 137.780 230.020 138.680 230.300 ;
        RECT 139.620 230.020 140.520 230.300 ;
        RECT 141.460 230.020 142.360 230.300 ;
        RECT 143.300 230.020 144.200 230.300 ;
        RECT 145.140 230.020 146.500 230.300 ;
        RECT 147.440 230.020 148.340 230.300 ;
        RECT 149.280 230.020 150.180 230.300 ;
        RECT 151.120 230.020 152.020 230.300 ;
        RECT 152.960 230.020 153.860 230.300 ;
        RECT 154.800 230.020 155.700 230.300 ;
        RECT 156.640 230.020 157.540 230.300 ;
        RECT 158.480 230.020 159.380 230.300 ;
        RECT 160.320 230.020 161.220 230.300 ;
        RECT 162.160 230.020 163.060 230.300 ;
        RECT 164.000 230.020 164.900 230.300 ;
        RECT 165.840 230.020 167.200 230.300 ;
        RECT 168.140 230.020 169.040 230.300 ;
        RECT 169.980 230.020 170.880 230.300 ;
        RECT 171.820 230.020 172.720 230.300 ;
        RECT 173.660 230.020 174.560 230.300 ;
        RECT 175.500 230.020 176.400 230.300 ;
        RECT 177.340 230.020 180.220 230.300 ;
        RECT 1.470 0.980 180.220 230.020 ;
        RECT 1.470 0.270 3.440 0.980 ;
        RECT 4.380 0.270 5.280 0.980 ;
        RECT 6.220 0.270 7.120 0.980 ;
        RECT 8.060 0.270 8.960 0.980 ;
        RECT 9.900 0.270 10.800 0.980 ;
        RECT 11.740 0.270 12.640 0.980 ;
        RECT 13.580 0.270 14.480 0.980 ;
        RECT 15.420 0.270 16.780 0.980 ;
        RECT 17.720 0.270 18.620 0.980 ;
        RECT 19.560 0.270 20.460 0.980 ;
        RECT 21.400 0.270 22.300 0.980 ;
        RECT 23.240 0.270 24.140 0.980 ;
        RECT 25.080 0.270 25.980 0.980 ;
        RECT 26.920 0.270 27.820 0.980 ;
        RECT 28.760 0.270 29.660 0.980 ;
        RECT 30.600 0.270 31.500 0.980 ;
        RECT 32.440 0.270 33.340 0.980 ;
        RECT 34.280 0.270 35.180 0.980 ;
        RECT 36.120 0.270 37.480 0.980 ;
        RECT 38.420 0.270 39.320 0.980 ;
        RECT 40.260 0.270 41.160 0.980 ;
        RECT 42.100 0.270 43.000 0.980 ;
        RECT 43.940 0.270 44.840 0.980 ;
        RECT 45.780 0.270 46.680 0.980 ;
        RECT 47.620 0.270 48.520 0.980 ;
        RECT 49.460 0.270 50.360 0.980 ;
        RECT 51.300 0.270 52.200 0.980 ;
        RECT 53.140 0.270 54.040 0.980 ;
        RECT 54.980 0.270 55.880 0.980 ;
        RECT 56.820 0.270 57.720 0.980 ;
        RECT 58.660 0.270 60.020 0.980 ;
        RECT 60.960 0.270 61.860 0.980 ;
        RECT 62.800 0.270 63.700 0.980 ;
        RECT 64.640 0.270 65.540 0.980 ;
        RECT 66.480 0.270 67.380 0.980 ;
        RECT 68.320 0.270 69.220 0.980 ;
        RECT 70.160 0.270 71.060 0.980 ;
        RECT 72.000 0.270 72.900 0.980 ;
        RECT 73.840 0.270 74.740 0.980 ;
        RECT 75.680 0.270 76.580 0.980 ;
        RECT 77.520 0.270 78.420 0.980 ;
        RECT 79.360 0.270 80.720 0.980 ;
        RECT 81.660 0.270 82.560 0.980 ;
        RECT 83.500 0.270 84.400 0.980 ;
        RECT 85.340 0.270 86.240 0.980 ;
        RECT 87.180 0.270 88.080 0.980 ;
        RECT 89.020 0.270 89.920 0.980 ;
        RECT 90.860 0.270 91.760 0.980 ;
        RECT 92.700 0.270 93.600 0.980 ;
        RECT 94.540 0.270 95.440 0.980 ;
        RECT 96.380 0.270 97.280 0.980 ;
        RECT 98.220 0.270 99.120 0.980 ;
        RECT 100.060 0.270 100.960 0.980 ;
        RECT 101.900 0.270 103.260 0.980 ;
        RECT 104.200 0.270 105.100 0.980 ;
        RECT 106.040 0.270 106.940 0.980 ;
        RECT 107.880 0.270 108.780 0.980 ;
        RECT 109.720 0.270 110.620 0.980 ;
        RECT 111.560 0.270 112.460 0.980 ;
        RECT 113.400 0.270 114.300 0.980 ;
        RECT 115.240 0.270 116.140 0.980 ;
        RECT 117.080 0.270 117.980 0.980 ;
        RECT 118.920 0.270 119.820 0.980 ;
        RECT 120.760 0.270 121.660 0.980 ;
        RECT 122.600 0.270 123.960 0.980 ;
        RECT 124.900 0.270 125.800 0.980 ;
        RECT 126.740 0.270 127.640 0.980 ;
        RECT 128.580 0.270 129.480 0.980 ;
        RECT 130.420 0.270 131.320 0.980 ;
        RECT 132.260 0.270 133.160 0.980 ;
        RECT 134.100 0.270 135.000 0.980 ;
        RECT 135.940 0.270 136.840 0.980 ;
        RECT 137.780 0.270 138.680 0.980 ;
        RECT 139.620 0.270 140.520 0.980 ;
        RECT 141.460 0.270 142.360 0.980 ;
        RECT 143.300 0.270 144.200 0.980 ;
        RECT 145.140 0.270 146.500 0.980 ;
        RECT 147.440 0.270 148.340 0.980 ;
        RECT 149.280 0.270 150.180 0.980 ;
        RECT 151.120 0.270 152.020 0.980 ;
        RECT 152.960 0.270 153.860 0.980 ;
        RECT 154.800 0.270 155.700 0.980 ;
        RECT 156.640 0.270 157.540 0.980 ;
        RECT 158.480 0.270 159.380 0.980 ;
        RECT 160.320 0.270 161.220 0.980 ;
        RECT 162.160 0.270 163.060 0.980 ;
        RECT 164.000 0.270 164.900 0.980 ;
        RECT 165.840 0.270 167.200 0.980 ;
        RECT 168.140 0.270 169.040 0.980 ;
        RECT 169.980 0.270 170.880 0.980 ;
        RECT 171.820 0.270 172.720 0.980 ;
        RECT 173.660 0.270 174.560 0.980 ;
        RECT 175.500 0.270 176.400 0.980 ;
        RECT 177.340 0.270 180.220 0.980 ;
      LAYER met3 ;
        RECT 0.700 225.510 179.900 226.250 ;
        RECT 0.700 225.330 180.300 225.510 ;
        RECT 1.100 224.150 180.300 225.330 ;
        RECT 0.700 223.970 180.300 224.150 ;
        RECT 0.700 223.290 179.900 223.970 ;
        RECT 1.100 222.790 179.900 223.290 ;
        RECT 1.100 222.110 180.300 222.790 ;
        RECT 0.700 221.930 180.300 222.110 ;
        RECT 1.100 221.250 180.300 221.930 ;
        RECT 1.100 220.750 179.900 221.250 ;
        RECT 0.700 220.070 179.900 220.750 ;
        RECT 0.700 219.890 180.300 220.070 ;
        RECT 1.100 218.710 180.300 219.890 ;
        RECT 0.700 218.530 180.300 218.710 ;
        RECT 1.100 217.350 179.900 218.530 ;
        RECT 0.700 216.490 180.300 217.350 ;
        RECT 1.100 215.310 180.300 216.490 ;
        RECT 0.700 215.130 180.300 215.310 ;
        RECT 1.100 213.950 179.900 215.130 ;
        RECT 0.700 213.090 180.300 213.950 ;
        RECT 1.100 212.410 180.300 213.090 ;
        RECT 1.100 211.910 179.900 212.410 ;
        RECT 0.700 211.730 179.900 211.910 ;
        RECT 1.100 211.230 179.900 211.730 ;
        RECT 1.100 210.550 180.300 211.230 ;
        RECT 0.700 209.690 180.300 210.550 ;
        RECT 1.100 208.510 179.900 209.690 ;
        RECT 0.700 207.650 180.300 208.510 ;
        RECT 1.100 206.970 180.300 207.650 ;
        RECT 1.100 206.470 179.900 206.970 ;
        RECT 0.700 206.290 179.900 206.470 ;
        RECT 1.100 205.790 179.900 206.290 ;
        RECT 1.100 205.110 180.300 205.790 ;
        RECT 0.700 204.250 180.300 205.110 ;
        RECT 1.100 203.070 179.900 204.250 ;
        RECT 0.700 202.890 180.300 203.070 ;
        RECT 1.100 201.710 180.300 202.890 ;
        RECT 0.700 201.530 180.300 201.710 ;
        RECT 0.700 200.850 179.900 201.530 ;
        RECT 1.100 200.350 179.900 200.850 ;
        RECT 1.100 199.670 180.300 200.350 ;
        RECT 0.700 199.490 180.300 199.670 ;
        RECT 1.100 198.810 180.300 199.490 ;
        RECT 1.100 198.310 179.900 198.810 ;
        RECT 0.700 197.630 179.900 198.310 ;
        RECT 0.700 197.450 180.300 197.630 ;
        RECT 1.100 196.270 180.300 197.450 ;
        RECT 0.700 196.090 180.300 196.270 ;
        RECT 0.700 195.410 179.900 196.090 ;
        RECT 1.100 194.910 179.900 195.410 ;
        RECT 1.100 194.230 180.300 194.910 ;
        RECT 0.700 194.050 180.300 194.230 ;
        RECT 1.100 192.870 180.300 194.050 ;
        RECT 0.700 192.690 180.300 192.870 ;
        RECT 0.700 192.010 179.900 192.690 ;
        RECT 1.100 191.510 179.900 192.010 ;
        RECT 1.100 190.830 180.300 191.510 ;
        RECT 0.700 190.650 180.300 190.830 ;
        RECT 1.100 189.970 180.300 190.650 ;
        RECT 1.100 189.470 179.900 189.970 ;
        RECT 0.700 188.790 179.900 189.470 ;
        RECT 0.700 188.610 180.300 188.790 ;
        RECT 1.100 187.430 180.300 188.610 ;
        RECT 0.700 187.250 180.300 187.430 ;
        RECT 1.100 186.070 179.900 187.250 ;
        RECT 0.700 185.210 180.300 186.070 ;
        RECT 1.100 184.530 180.300 185.210 ;
        RECT 1.100 184.030 179.900 184.530 ;
        RECT 0.700 183.850 179.900 184.030 ;
        RECT 1.100 183.350 179.900 183.850 ;
        RECT 1.100 182.670 180.300 183.350 ;
        RECT 0.700 181.810 180.300 182.670 ;
        RECT 1.100 180.630 179.900 181.810 ;
        RECT 0.700 179.770 180.300 180.630 ;
        RECT 1.100 179.090 180.300 179.770 ;
        RECT 1.100 178.590 179.900 179.090 ;
        RECT 0.700 178.410 179.900 178.590 ;
        RECT 1.100 177.910 179.900 178.410 ;
        RECT 1.100 177.230 180.300 177.910 ;
        RECT 0.700 176.370 180.300 177.230 ;
        RECT 1.100 175.190 179.900 176.370 ;
        RECT 0.700 175.010 180.300 175.190 ;
        RECT 1.100 173.830 180.300 175.010 ;
        RECT 0.700 173.650 180.300 173.830 ;
        RECT 0.700 172.970 179.900 173.650 ;
        RECT 1.100 172.470 179.900 172.970 ;
        RECT 1.100 171.790 180.300 172.470 ;
        RECT 0.700 171.610 180.300 171.790 ;
        RECT 1.100 170.930 180.300 171.610 ;
        RECT 1.100 170.430 179.900 170.930 ;
        RECT 0.700 169.750 179.900 170.430 ;
        RECT 0.700 169.570 180.300 169.750 ;
        RECT 1.100 168.390 180.300 169.570 ;
        RECT 0.700 168.210 180.300 168.390 ;
        RECT 1.100 167.530 180.300 168.210 ;
        RECT 1.100 167.030 179.900 167.530 ;
        RECT 0.700 166.350 179.900 167.030 ;
        RECT 0.700 166.170 180.300 166.350 ;
        RECT 1.100 164.990 180.300 166.170 ;
        RECT 0.700 164.810 180.300 164.990 ;
        RECT 0.700 164.130 179.900 164.810 ;
        RECT 1.100 163.630 179.900 164.130 ;
        RECT 1.100 162.950 180.300 163.630 ;
        RECT 0.700 162.770 180.300 162.950 ;
        RECT 1.100 162.090 180.300 162.770 ;
        RECT 1.100 161.590 179.900 162.090 ;
        RECT 0.700 160.910 179.900 161.590 ;
        RECT 0.700 160.730 180.300 160.910 ;
        RECT 1.100 159.550 180.300 160.730 ;
        RECT 0.700 159.370 180.300 159.550 ;
        RECT 1.100 158.190 179.900 159.370 ;
        RECT 0.700 157.330 180.300 158.190 ;
        RECT 1.100 156.650 180.300 157.330 ;
        RECT 1.100 156.150 179.900 156.650 ;
        RECT 0.700 155.970 179.900 156.150 ;
        RECT 1.100 155.470 179.900 155.970 ;
        RECT 1.100 154.790 180.300 155.470 ;
        RECT 0.700 153.930 180.300 154.790 ;
        RECT 1.100 152.750 179.900 153.930 ;
        RECT 0.700 152.570 180.300 152.750 ;
        RECT 1.100 151.390 180.300 152.570 ;
        RECT 0.700 151.210 180.300 151.390 ;
        RECT 0.700 150.530 179.900 151.210 ;
        RECT 1.100 150.030 179.900 150.530 ;
        RECT 1.100 149.350 180.300 150.030 ;
        RECT 0.700 148.490 180.300 149.350 ;
        RECT 1.100 147.310 179.900 148.490 ;
        RECT 0.700 147.130 180.300 147.310 ;
        RECT 1.100 145.950 180.300 147.130 ;
        RECT 0.700 145.090 180.300 145.950 ;
        RECT 1.100 143.910 179.900 145.090 ;
        RECT 0.700 143.730 180.300 143.910 ;
        RECT 1.100 142.550 180.300 143.730 ;
        RECT 0.700 142.370 180.300 142.550 ;
        RECT 0.700 141.690 179.900 142.370 ;
        RECT 1.100 141.190 179.900 141.690 ;
        RECT 1.100 140.510 180.300 141.190 ;
        RECT 0.700 140.330 180.300 140.510 ;
        RECT 1.100 139.650 180.300 140.330 ;
        RECT 1.100 139.150 179.900 139.650 ;
        RECT 0.700 138.470 179.900 139.150 ;
        RECT 0.700 138.290 180.300 138.470 ;
        RECT 1.100 137.110 180.300 138.290 ;
        RECT 0.700 136.930 180.300 137.110 ;
        RECT 0.700 136.250 179.900 136.930 ;
        RECT 1.100 135.750 179.900 136.250 ;
        RECT 1.100 135.070 180.300 135.750 ;
        RECT 0.700 134.890 180.300 135.070 ;
        RECT 1.100 134.210 180.300 134.890 ;
        RECT 1.100 133.710 179.900 134.210 ;
        RECT 0.700 133.030 179.900 133.710 ;
        RECT 0.700 132.850 180.300 133.030 ;
        RECT 1.100 131.670 180.300 132.850 ;
        RECT 0.700 131.490 180.300 131.670 ;
        RECT 1.100 130.310 179.900 131.490 ;
        RECT 0.700 129.450 180.300 130.310 ;
        RECT 1.100 128.770 180.300 129.450 ;
        RECT 1.100 128.270 179.900 128.770 ;
        RECT 0.700 128.090 179.900 128.270 ;
        RECT 1.100 127.590 179.900 128.090 ;
        RECT 1.100 126.910 180.300 127.590 ;
        RECT 0.700 126.050 180.300 126.910 ;
        RECT 1.100 124.870 179.900 126.050 ;
        RECT 0.700 124.690 180.300 124.870 ;
        RECT 1.100 123.510 180.300 124.690 ;
        RECT 0.700 123.330 180.300 123.510 ;
        RECT 0.700 122.650 179.900 123.330 ;
        RECT 1.100 122.150 179.900 122.650 ;
        RECT 1.100 121.470 180.300 122.150 ;
        RECT 0.700 120.610 180.300 121.470 ;
        RECT 1.100 119.930 180.300 120.610 ;
        RECT 1.100 119.430 179.900 119.930 ;
        RECT 0.700 119.250 179.900 119.430 ;
        RECT 1.100 118.750 179.900 119.250 ;
        RECT 1.100 118.070 180.300 118.750 ;
        RECT 0.700 117.210 180.300 118.070 ;
        RECT 1.100 116.030 179.900 117.210 ;
        RECT 0.700 115.850 180.300 116.030 ;
        RECT 1.100 114.670 180.300 115.850 ;
        RECT 0.700 114.490 180.300 114.670 ;
        RECT 0.700 113.810 179.900 114.490 ;
        RECT 1.100 113.310 179.900 113.810 ;
        RECT 1.100 112.630 180.300 113.310 ;
        RECT 0.700 112.450 180.300 112.630 ;
        RECT 1.100 111.770 180.300 112.450 ;
        RECT 1.100 111.270 179.900 111.770 ;
        RECT 0.700 110.590 179.900 111.270 ;
        RECT 0.700 110.410 180.300 110.590 ;
        RECT 1.100 109.230 180.300 110.410 ;
        RECT 0.700 109.050 180.300 109.230 ;
        RECT 1.100 107.870 179.900 109.050 ;
        RECT 0.700 107.010 180.300 107.870 ;
        RECT 1.100 106.330 180.300 107.010 ;
        RECT 1.100 105.830 179.900 106.330 ;
        RECT 0.700 105.150 179.900 105.830 ;
        RECT 0.700 104.970 180.300 105.150 ;
        RECT 1.100 103.790 180.300 104.970 ;
        RECT 0.700 103.610 180.300 103.790 ;
        RECT 1.100 102.430 179.900 103.610 ;
        RECT 0.700 101.570 180.300 102.430 ;
        RECT 1.100 100.890 180.300 101.570 ;
        RECT 1.100 100.390 179.900 100.890 ;
        RECT 0.700 100.210 179.900 100.390 ;
        RECT 1.100 99.710 179.900 100.210 ;
        RECT 1.100 99.030 180.300 99.710 ;
        RECT 0.700 98.170 180.300 99.030 ;
        RECT 1.100 97.490 180.300 98.170 ;
        RECT 1.100 96.990 179.900 97.490 ;
        RECT 0.700 96.810 179.900 96.990 ;
        RECT 1.100 96.310 179.900 96.810 ;
        RECT 1.100 95.630 180.300 96.310 ;
        RECT 0.700 94.770 180.300 95.630 ;
        RECT 1.100 93.590 179.900 94.770 ;
        RECT 0.700 93.410 180.300 93.590 ;
        RECT 1.100 92.230 180.300 93.410 ;
        RECT 0.700 92.050 180.300 92.230 ;
        RECT 0.700 91.370 179.900 92.050 ;
        RECT 1.100 90.870 179.900 91.370 ;
        RECT 1.100 90.190 180.300 90.870 ;
        RECT 0.700 89.330 180.300 90.190 ;
        RECT 1.100 88.150 179.900 89.330 ;
        RECT 0.700 87.970 180.300 88.150 ;
        RECT 1.100 86.790 180.300 87.970 ;
        RECT 0.700 86.610 180.300 86.790 ;
        RECT 0.700 85.930 179.900 86.610 ;
        RECT 1.100 85.430 179.900 85.930 ;
        RECT 1.100 84.750 180.300 85.430 ;
        RECT 0.700 84.570 180.300 84.750 ;
        RECT 1.100 83.890 180.300 84.570 ;
        RECT 1.100 83.390 179.900 83.890 ;
        RECT 0.700 82.710 179.900 83.390 ;
        RECT 0.700 82.530 180.300 82.710 ;
        RECT 1.100 81.350 180.300 82.530 ;
        RECT 0.700 81.170 180.300 81.350 ;
        RECT 1.100 79.990 179.900 81.170 ;
        RECT 0.700 79.130 180.300 79.990 ;
        RECT 1.100 78.450 180.300 79.130 ;
        RECT 1.100 77.950 179.900 78.450 ;
        RECT 0.700 77.270 179.900 77.950 ;
        RECT 0.700 77.090 180.300 77.270 ;
        RECT 1.100 75.910 180.300 77.090 ;
        RECT 0.700 75.730 180.300 75.910 ;
        RECT 1.100 74.550 179.900 75.730 ;
        RECT 0.700 73.690 180.300 74.550 ;
        RECT 1.100 72.510 180.300 73.690 ;
        RECT 0.700 72.330 180.300 72.510 ;
        RECT 1.100 71.150 179.900 72.330 ;
        RECT 0.700 70.290 180.300 71.150 ;
        RECT 1.100 69.610 180.300 70.290 ;
        RECT 1.100 69.110 179.900 69.610 ;
        RECT 0.700 68.930 179.900 69.110 ;
        RECT 1.100 68.430 179.900 68.930 ;
        RECT 1.100 67.750 180.300 68.430 ;
        RECT 0.700 66.890 180.300 67.750 ;
        RECT 1.100 65.710 179.900 66.890 ;
        RECT 0.700 65.530 180.300 65.710 ;
        RECT 1.100 64.350 180.300 65.530 ;
        RECT 0.700 64.170 180.300 64.350 ;
        RECT 0.700 63.490 179.900 64.170 ;
        RECT 1.100 62.990 179.900 63.490 ;
        RECT 1.100 62.310 180.300 62.990 ;
        RECT 0.700 61.450 180.300 62.310 ;
        RECT 1.100 60.270 179.900 61.450 ;
        RECT 0.700 60.090 180.300 60.270 ;
        RECT 1.100 58.910 180.300 60.090 ;
        RECT 0.700 58.730 180.300 58.910 ;
        RECT 0.700 58.050 179.900 58.730 ;
        RECT 1.100 57.550 179.900 58.050 ;
        RECT 1.100 56.870 180.300 57.550 ;
        RECT 0.700 56.690 180.300 56.870 ;
        RECT 1.100 56.010 180.300 56.690 ;
        RECT 1.100 55.510 179.900 56.010 ;
        RECT 0.700 54.830 179.900 55.510 ;
        RECT 0.700 54.650 180.300 54.830 ;
        RECT 1.100 53.470 180.300 54.650 ;
        RECT 0.700 53.290 180.300 53.470 ;
        RECT 1.100 52.110 179.900 53.290 ;
        RECT 0.700 51.250 180.300 52.110 ;
        RECT 1.100 50.070 180.300 51.250 ;
        RECT 0.700 49.890 180.300 50.070 ;
        RECT 1.100 48.710 179.900 49.890 ;
        RECT 0.700 47.850 180.300 48.710 ;
        RECT 1.100 47.170 180.300 47.850 ;
        RECT 1.100 46.670 179.900 47.170 ;
        RECT 0.700 45.990 179.900 46.670 ;
        RECT 0.700 45.810 180.300 45.990 ;
        RECT 1.100 44.630 180.300 45.810 ;
        RECT 0.700 44.450 180.300 44.630 ;
        RECT 1.100 43.270 179.900 44.450 ;
        RECT 0.700 42.410 180.300 43.270 ;
        RECT 1.100 41.730 180.300 42.410 ;
        RECT 1.100 41.230 179.900 41.730 ;
        RECT 0.700 41.050 179.900 41.230 ;
        RECT 1.100 40.550 179.900 41.050 ;
        RECT 1.100 39.870 180.300 40.550 ;
        RECT 0.700 39.010 180.300 39.870 ;
        RECT 1.100 37.830 179.900 39.010 ;
        RECT 0.700 37.650 180.300 37.830 ;
        RECT 1.100 36.470 180.300 37.650 ;
        RECT 0.700 36.290 180.300 36.470 ;
        RECT 0.700 35.610 179.900 36.290 ;
        RECT 1.100 35.110 179.900 35.610 ;
        RECT 1.100 34.430 180.300 35.110 ;
        RECT 0.700 34.250 180.300 34.430 ;
        RECT 1.100 33.570 180.300 34.250 ;
        RECT 1.100 33.070 179.900 33.570 ;
        RECT 0.700 32.390 179.900 33.070 ;
        RECT 0.700 32.210 180.300 32.390 ;
        RECT 1.100 31.030 180.300 32.210 ;
        RECT 0.700 30.850 180.300 31.030 ;
        RECT 0.700 30.170 179.900 30.850 ;
        RECT 1.100 29.670 179.900 30.170 ;
        RECT 1.100 28.990 180.300 29.670 ;
        RECT 0.700 28.810 180.300 28.990 ;
        RECT 1.100 28.130 180.300 28.810 ;
        RECT 1.100 27.630 179.900 28.130 ;
        RECT 0.700 26.950 179.900 27.630 ;
        RECT 0.700 26.770 180.300 26.950 ;
        RECT 1.100 25.590 180.300 26.770 ;
        RECT 0.700 25.410 180.300 25.590 ;
        RECT 1.100 24.730 180.300 25.410 ;
        RECT 1.100 24.230 179.900 24.730 ;
        RECT 0.700 23.550 179.900 24.230 ;
        RECT 0.700 23.370 180.300 23.550 ;
        RECT 1.100 22.190 180.300 23.370 ;
        RECT 0.700 22.010 180.300 22.190 ;
        RECT 1.100 20.830 179.900 22.010 ;
        RECT 0.700 19.970 180.300 20.830 ;
        RECT 1.100 19.290 180.300 19.970 ;
        RECT 1.100 18.790 179.900 19.290 ;
        RECT 0.700 18.110 179.900 18.790 ;
        RECT 0.700 17.930 180.300 18.110 ;
        RECT 1.100 16.750 180.300 17.930 ;
        RECT 0.700 16.570 180.300 16.750 ;
        RECT 1.100 15.390 179.900 16.570 ;
        RECT 0.700 14.530 180.300 15.390 ;
        RECT 1.100 13.850 180.300 14.530 ;
        RECT 1.100 13.350 179.900 13.850 ;
        RECT 0.700 13.170 179.900 13.350 ;
        RECT 1.100 12.670 179.900 13.170 ;
        RECT 1.100 11.990 180.300 12.670 ;
        RECT 0.700 11.130 180.300 11.990 ;
        RECT 1.100 9.950 179.900 11.130 ;
        RECT 0.700 9.770 180.300 9.950 ;
        RECT 1.100 8.590 180.300 9.770 ;
        RECT 0.700 8.410 180.300 8.590 ;
        RECT 0.700 7.730 179.900 8.410 ;
        RECT 1.100 7.230 179.900 7.730 ;
        RECT 1.100 6.550 180.300 7.230 ;
        RECT 0.700 6.370 180.300 6.550 ;
        RECT 1.100 5.690 180.300 6.370 ;
        RECT 1.100 5.190 179.900 5.690 ;
        RECT 0.700 4.510 179.900 5.190 ;
        RECT 0.700 4.330 180.300 4.510 ;
        RECT 1.100 3.575 180.300 4.330 ;
      LAYER met4 ;
        RECT 8.575 3.575 20.180 224.225 ;
        RECT 22.580 3.575 23.480 224.225 ;
        RECT 25.880 3.575 172.665 224.225 ;
  END
END RAM_IO
END LIBRARY

