magic
tech sky130A
magscale 1 2
timestamp 1732488443
<< viali >>
rect 1869 43401 1903 43435
rect 2789 43401 2823 43435
rect 3157 43401 3191 43435
rect 4629 43401 4663 43435
rect 5549 43401 5583 43435
rect 6101 43401 6135 43435
rect 6377 43401 6411 43435
rect 7021 43401 7055 43435
rect 7389 43401 7423 43435
rect 7757 43401 7791 43435
rect 8309 43401 8343 43435
rect 8677 43401 8711 43435
rect 9229 43401 9263 43435
rect 9781 43401 9815 43435
rect 10517 43401 10551 43435
rect 12265 43401 12299 43435
rect 20085 43401 20119 43435
rect 21005 43401 21039 43435
rect 22017 43401 22051 43435
rect 22385 43401 22419 43435
rect 22937 43401 22971 43435
rect 23489 43401 23523 43435
rect 6745 43333 6779 43367
rect 8033 43333 8067 43367
rect 12449 43333 12483 43367
rect 12817 43333 12851 43367
rect 14197 43333 14231 43367
rect 14749 43333 14783 43367
rect 15117 43333 15151 43367
rect 16313 43333 16347 43367
rect 16773 43333 16807 43367
rect 1593 43265 1627 43299
rect 1777 43265 1811 43299
rect 2513 43265 2547 43299
rect 3065 43265 3099 43299
rect 3985 43265 4019 43299
rect 4537 43265 4571 43299
rect 5273 43265 5307 43299
rect 5917 43265 5951 43299
rect 6561 43265 6595 43299
rect 7205 43265 7239 43299
rect 7573 43265 7607 43299
rect 8493 43265 8527 43299
rect 9045 43265 9079 43299
rect 9505 43265 9539 43299
rect 9965 43265 9999 43299
rect 10333 43265 10367 43299
rect 10701 43265 10735 43299
rect 11069 43265 11103 43299
rect 11529 43265 11563 43299
rect 12081 43265 12115 43299
rect 13645 43265 13679 43299
rect 15485 43265 15519 43299
rect 15853 43265 15887 43299
rect 16497 43265 16531 43299
rect 17509 43265 17543 43299
rect 17785 43265 17819 43299
rect 18061 43265 18095 43299
rect 18337 43265 18371 43299
rect 18613 43265 18647 43299
rect 18889 43265 18923 43299
rect 19441 43265 19475 43299
rect 19717 43265 19751 43299
rect 19901 43265 19935 43299
rect 20361 43265 20395 43299
rect 20913 43265 20947 43299
rect 21373 43265 21407 43299
rect 21833 43265 21867 43299
rect 22293 43265 22327 43299
rect 22845 43265 22879 43299
rect 23397 43265 23431 43299
rect 23949 43265 23983 43299
rect 3801 43129 3835 43163
rect 14933 43129 14967 43163
rect 17877 43129 17911 43163
rect 19257 43129 19291 43163
rect 20637 43129 20671 43163
rect 21557 43129 21591 43163
rect 1409 43061 1443 43095
rect 4353 43061 4387 43095
rect 10149 43061 10183 43095
rect 10885 43061 10919 43095
rect 11253 43061 11287 43095
rect 11713 43061 11747 43095
rect 12541 43061 12575 43095
rect 12909 43061 12943 43095
rect 13829 43061 13863 43095
rect 14289 43061 14323 43095
rect 15209 43061 15243 43095
rect 15669 43061 15703 43095
rect 16037 43061 16071 43095
rect 16865 43061 16899 43095
rect 17325 43061 17359 43095
rect 17601 43061 17635 43095
rect 18153 43061 18187 43095
rect 18429 43061 18463 43095
rect 18705 43061 18739 43095
rect 19533 43061 19567 43095
rect 24133 43061 24167 43095
rect 2237 42857 2271 42891
rect 3341 42857 3375 42891
rect 4169 42857 4203 42891
rect 6101 42857 6135 42891
rect 6837 42857 6871 42891
rect 7389 42857 7423 42891
rect 10333 42857 10367 42891
rect 10609 42857 10643 42891
rect 16313 42857 16347 42891
rect 18889 42857 18923 42891
rect 8953 42789 8987 42823
rect 18061 42789 18095 42823
rect 1777 42721 1811 42755
rect 2973 42721 3007 42755
rect 5365 42721 5399 42755
rect 8677 42721 8711 42755
rect 9781 42721 9815 42755
rect 23489 42721 23523 42755
rect 2145 42653 2179 42687
rect 4537 42653 4571 42687
rect 5089 42653 5123 42687
rect 5549 42653 5583 42687
rect 7757 42653 7791 42687
rect 9137 42653 9171 42687
rect 9505 42653 9539 42687
rect 10057 42653 10091 42687
rect 10517 42653 10551 42687
rect 10793 42653 10827 42687
rect 11621 42653 11655 42687
rect 11897 42653 11931 42687
rect 12725 42653 12759 42687
rect 13001 42653 13035 42687
rect 14105 42653 14139 42687
rect 14381 42653 14415 42687
rect 14657 42653 14691 42687
rect 15301 42653 15335 42687
rect 15577 42653 15611 42687
rect 16497 42653 16531 42687
rect 16589 42653 16623 42687
rect 17141 42653 17175 42687
rect 17417 42653 17451 42687
rect 17693 42653 17727 42687
rect 17969 42653 18003 42687
rect 18245 42653 18279 42687
rect 18521 42653 18555 42687
rect 18797 42653 18831 42687
rect 19073 42653 19107 42687
rect 19257 42653 19291 42687
rect 21281 42653 21315 42687
rect 21925 42653 21959 42687
rect 22661 42653 22695 42687
rect 23213 42653 23247 42687
rect 24133 42653 24167 42687
rect 1501 42585 1535 42619
rect 2697 42585 2731 42619
rect 3249 42585 3283 42619
rect 4077 42585 4111 42619
rect 6009 42585 6043 42619
rect 6745 42585 6779 42619
rect 7297 42585 7331 42619
rect 8401 42585 8435 42619
rect 21557 42585 21591 42619
rect 22109 42585 22143 42619
rect 22477 42585 22511 42619
rect 23765 42585 23799 42619
rect 4721 42517 4755 42551
rect 5733 42517 5767 42551
rect 7941 42517 7975 42551
rect 10241 42517 10275 42551
rect 11805 42517 11839 42551
rect 12081 42517 12115 42551
rect 12909 42517 12943 42551
rect 13185 42517 13219 42551
rect 14289 42517 14323 42551
rect 14565 42517 14599 42551
rect 14841 42517 14875 42551
rect 15485 42517 15519 42551
rect 15761 42517 15795 42551
rect 16773 42517 16807 42551
rect 16957 42517 16991 42551
rect 17233 42517 17267 42551
rect 17509 42517 17543 42551
rect 17785 42517 17819 42551
rect 18337 42517 18371 42551
rect 18613 42517 18647 42551
rect 20545 42517 20579 42551
rect 21097 42517 21131 42551
rect 22753 42517 22787 42551
rect 1593 42313 1627 42347
rect 2513 42313 2547 42347
rect 3433 42313 3467 42347
rect 3709 42313 3743 42347
rect 4997 42313 5031 42347
rect 5181 42313 5215 42347
rect 6009 42313 6043 42347
rect 8493 42313 8527 42347
rect 9965 42313 9999 42347
rect 19717 42313 19751 42347
rect 19993 42313 20027 42347
rect 20545 42313 20579 42347
rect 20821 42313 20855 42347
rect 21833 42313 21867 42347
rect 22569 42313 22603 42347
rect 23121 42313 23155 42347
rect 23673 42313 23707 42347
rect 1501 42245 1535 42279
rect 2053 42245 2087 42279
rect 16773 42245 16807 42279
rect 17141 42245 17175 42279
rect 17509 42245 17543 42279
rect 17877 42245 17911 42279
rect 18245 42245 18279 42279
rect 18613 42245 18647 42279
rect 18981 42245 19015 42279
rect 19349 42245 19383 42279
rect 2697 42177 2731 42211
rect 2789 42177 2823 42211
rect 3617 42177 3651 42211
rect 3893 42177 3927 42211
rect 3985 42177 4019 42211
rect 4721 42177 4755 42211
rect 4813 42177 4847 42211
rect 5365 42177 5399 42211
rect 5733 42177 5767 42211
rect 6193 42177 6227 42211
rect 6561 42177 6595 42211
rect 6837 42177 6871 42211
rect 7481 42177 7515 42211
rect 7941 42177 7975 42211
rect 8217 42177 8251 42211
rect 8401 42177 8435 42211
rect 9045 42177 9079 42211
rect 9413 42177 9447 42211
rect 9873 42177 9907 42211
rect 10149 42177 10183 42211
rect 16129 42177 16163 42211
rect 19901 42177 19935 42211
rect 20177 42177 20211 42211
rect 20453 42177 20487 42211
rect 20729 42177 20763 42211
rect 21005 42177 21039 42211
rect 21281 42177 21315 42211
rect 21649 42177 21683 42211
rect 22017 42177 22051 42211
rect 22293 42177 22327 42211
rect 22845 42177 22879 42211
rect 23397 42177 23431 42211
rect 24041 42177 24075 42211
rect 7205 42109 7239 42143
rect 2973 42041 3007 42075
rect 4169 42041 4203 42075
rect 6377 42041 6411 42075
rect 6653 42041 6687 42075
rect 9689 42041 9723 42075
rect 16957 42041 16991 42075
rect 17325 42041 17359 42075
rect 17693 42041 17727 42075
rect 18061 42041 18095 42075
rect 19165 42041 19199 42075
rect 19533 42041 19567 42075
rect 2145 41973 2179 42007
rect 4537 41973 4571 42007
rect 7297 41973 7331 42007
rect 7757 41973 7791 42007
rect 8033 41973 8067 42007
rect 8861 41973 8895 42007
rect 16313 41973 16347 42007
rect 18337 41973 18371 42007
rect 18705 41973 18739 42007
rect 20269 41973 20303 42007
rect 24317 41973 24351 42007
rect 1593 41769 1627 41803
rect 2145 41769 2179 41803
rect 2513 41769 2547 41803
rect 3157 41769 3191 41803
rect 3433 41769 3467 41803
rect 4077 41769 4111 41803
rect 4629 41769 4663 41803
rect 5733 41769 5767 41803
rect 7205 41769 7239 41803
rect 7573 41769 7607 41803
rect 8125 41769 8159 41803
rect 8401 41769 8435 41803
rect 8953 41769 8987 41803
rect 18797 41769 18831 41803
rect 19625 41769 19659 41803
rect 20729 41769 20763 41803
rect 23029 41769 23063 41803
rect 24133 41769 24167 41803
rect 3801 41701 3835 41735
rect 4353 41701 4387 41735
rect 4905 41701 4939 41735
rect 5457 41701 5491 41735
rect 6561 41701 6595 41735
rect 6929 41701 6963 41735
rect 10701 41701 10735 41735
rect 17969 41701 18003 41735
rect 19349 41701 19383 41735
rect 20913 41701 20947 41735
rect 23581 41701 23615 41735
rect 22477 41633 22511 41667
rect 2697 41565 2731 41599
rect 3341 41565 3375 41599
rect 3617 41565 3651 41599
rect 3985 41565 4019 41599
rect 4261 41565 4295 41599
rect 4537 41565 4571 41599
rect 4813 41565 4847 41599
rect 5089 41565 5123 41599
rect 5365 41565 5399 41599
rect 5641 41565 5675 41599
rect 5917 41565 5951 41599
rect 6745 41565 6779 41599
rect 7113 41565 7147 41599
rect 7389 41565 7423 41599
rect 7757 41565 7791 41599
rect 8033 41565 8067 41599
rect 8309 41565 8343 41599
rect 8585 41565 8619 41599
rect 9137 41565 9171 41599
rect 9689 41565 9723 41599
rect 9963 41565 9997 41599
rect 18153 41565 18187 41599
rect 18337 41565 18371 41599
rect 18981 41565 19015 41599
rect 19533 41565 19567 41599
rect 19809 41565 19843 41599
rect 20177 41565 20211 41599
rect 20453 41565 20487 41599
rect 20545 41565 20579 41599
rect 21097 41565 21131 41599
rect 21373 41565 21407 41599
rect 21649 41565 21683 41599
rect 21925 41565 21959 41599
rect 1501 41497 1535 41531
rect 2053 41497 2087 41531
rect 22201 41497 22235 41531
rect 22753 41497 22787 41531
rect 23305 41497 23339 41531
rect 23857 41497 23891 41531
rect 2973 41429 3007 41463
rect 5181 41429 5215 41463
rect 6193 41429 6227 41463
rect 7849 41429 7883 41463
rect 18429 41429 18463 41463
rect 19993 41429 20027 41463
rect 20269 41429 20303 41463
rect 21189 41429 21223 41463
rect 21465 41429 21499 41463
rect 21741 41429 21775 41463
rect 2697 41225 2731 41259
rect 7757 41225 7791 41259
rect 19533 41225 19567 41259
rect 19809 41225 19843 41259
rect 20361 41225 20395 41259
rect 20637 41225 20671 41259
rect 20913 41225 20947 41259
rect 21465 41225 21499 41259
rect 21833 41225 21867 41259
rect 22109 41225 22143 41259
rect 23121 41225 23155 41259
rect 24225 41225 24259 41259
rect 23949 41157 23983 41191
rect 1409 41089 1443 41123
rect 2237 41089 2271 41123
rect 2513 41089 2547 41123
rect 3249 41089 3283 41123
rect 3799 41089 3833 41123
rect 4905 41089 4939 41123
rect 5179 41089 5213 41123
rect 7941 41089 7975 41123
rect 8859 41089 8893 41123
rect 10057 41089 10091 41123
rect 10331 41089 10365 41123
rect 19257 41089 19291 41123
rect 19717 41089 19751 41123
rect 19993 41089 20027 41123
rect 20269 41089 20303 41123
rect 20545 41089 20579 41123
rect 20821 41089 20855 41123
rect 21097 41089 21131 41123
rect 21373 41089 21407 41123
rect 21649 41089 21683 41123
rect 22017 41089 22051 41123
rect 22293 41089 22327 41123
rect 22569 41089 22603 41123
rect 22845 41089 22879 41123
rect 23397 41089 23431 41123
rect 3525 41021 3559 41055
rect 8585 41021 8619 41055
rect 3065 40953 3099 40987
rect 6929 40953 6963 40987
rect 20085 40953 20119 40987
rect 4537 40885 4571 40919
rect 5917 40885 5951 40919
rect 7481 40885 7515 40919
rect 9597 40885 9631 40919
rect 11069 40885 11103 40919
rect 19073 40885 19107 40919
rect 21189 40885 21223 40919
rect 22385 40885 22419 40919
rect 23673 40885 23707 40919
rect 3433 40681 3467 40715
rect 20821 40681 20855 40715
rect 21097 40681 21131 40715
rect 22201 40681 22235 40715
rect 22477 40681 22511 40715
rect 22753 40681 22787 40715
rect 23029 40681 23063 40715
rect 23489 40681 23523 40715
rect 4813 40613 4847 40647
rect 10517 40613 10551 40647
rect 19533 40613 19567 40647
rect 20269 40613 20303 40647
rect 2237 40545 2271 40579
rect 3801 40545 3835 40579
rect 5549 40545 5583 40579
rect 10057 40545 10091 40579
rect 11069 40545 11103 40579
rect 11805 40545 11839 40579
rect 3617 40477 3651 40511
rect 4075 40477 4109 40511
rect 5823 40477 5857 40511
rect 6929 40477 6963 40511
rect 7203 40477 7237 40511
rect 9873 40477 9907 40511
rect 10793 40477 10827 40511
rect 10910 40477 10944 40511
rect 12063 40447 12097 40481
rect 13369 40477 13403 40511
rect 19349 40477 19383 40511
rect 19809 40477 19843 40511
rect 20177 40477 20211 40511
rect 20453 40477 20487 40511
rect 20729 40477 20763 40511
rect 21005 40477 21039 40511
rect 21281 40477 21315 40511
rect 21565 40477 21599 40511
rect 21833 40477 21867 40511
rect 22109 40477 22143 40511
rect 22385 40477 22419 40511
rect 22661 40477 22695 40511
rect 22937 40477 22971 40511
rect 23213 40477 23247 40511
rect 23673 40477 23707 40511
rect 1409 40409 1443 40443
rect 2421 40409 2455 40443
rect 3157 40409 3191 40443
rect 23857 40409 23891 40443
rect 24225 40409 24259 40443
rect 6561 40341 6595 40375
rect 7941 40341 7975 40375
rect 11713 40341 11747 40375
rect 12817 40341 12851 40375
rect 19625 40341 19659 40375
rect 19993 40341 20027 40375
rect 20545 40341 20579 40375
rect 21373 40341 21407 40375
rect 21649 40341 21683 40375
rect 21925 40341 21959 40375
rect 4169 40137 4203 40171
rect 7481 40137 7515 40171
rect 8585 40137 8619 40171
rect 20913 40137 20947 40171
rect 21189 40137 21223 40171
rect 21833 40137 21867 40171
rect 1685 40069 1719 40103
rect 3617 40069 3651 40103
rect 7757 40069 7791 40103
rect 7849 40069 7883 40103
rect 8217 40069 8251 40103
rect 9137 40069 9171 40103
rect 9413 40069 9447 40103
rect 9505 40069 9539 40103
rect 9873 40069 9907 40103
rect 10241 40069 10275 40103
rect 19257 40069 19291 40103
rect 1409 40001 1443 40035
rect 2219 40031 2253 40065
rect 3341 40001 3375 40035
rect 4353 40001 4387 40035
rect 4905 40001 4939 40035
rect 5179 40001 5213 40035
rect 11069 40001 11103 40035
rect 12725 40001 12759 40035
rect 19993 40001 20027 40035
rect 20269 40001 20303 40035
rect 20545 40001 20579 40035
rect 20821 40001 20855 40035
rect 21097 40001 21131 40035
rect 21373 40001 21407 40035
rect 21649 40001 21683 40035
rect 22017 40001 22051 40035
rect 22293 40001 22327 40035
rect 22569 40001 22603 40035
rect 22845 40001 22879 40035
rect 23121 40001 23155 40035
rect 23397 40001 23431 40035
rect 23857 40001 23891 40035
rect 24133 40001 24167 40035
rect 1961 39933 1995 39967
rect 11805 39933 11839 39967
rect 11989 39933 12023 39967
rect 12449 39933 12483 39967
rect 12842 39933 12876 39967
rect 13001 39933 13035 39967
rect 8769 39865 8803 39899
rect 19441 39865 19475 39899
rect 19809 39865 19843 39899
rect 20085 39865 20119 39899
rect 20361 39865 20395 39899
rect 20637 39865 20671 39899
rect 22661 39865 22695 39899
rect 23213 39865 23247 39899
rect 2973 39797 3007 39831
rect 4077 39797 4111 39831
rect 4629 39797 4663 39831
rect 5917 39797 5951 39831
rect 10425 39797 10459 39831
rect 13645 39797 13679 39831
rect 21465 39797 21499 39831
rect 22109 39797 22143 39831
rect 22385 39797 22419 39831
rect 22937 39797 22971 39831
rect 23673 39797 23707 39831
rect 24409 39797 24443 39831
rect 3433 39593 3467 39627
rect 8401 39593 8435 39627
rect 10517 39593 10551 39627
rect 13369 39593 13403 39627
rect 20729 39593 20763 39627
rect 21557 39593 21591 39627
rect 21833 39593 21867 39627
rect 22385 39593 22419 39627
rect 6101 39525 6135 39559
rect 22109 39525 22143 39559
rect 5457 39457 5491 39491
rect 6377 39457 6411 39491
rect 7389 39457 7423 39491
rect 12357 39457 12391 39491
rect 2237 39389 2271 39423
rect 3617 39389 3651 39423
rect 4353 39389 4387 39423
rect 5641 39389 5675 39423
rect 6494 39389 6528 39423
rect 6653 39389 6687 39423
rect 7663 39389 7697 39423
rect 9505 39389 9539 39423
rect 9779 39389 9813 39423
rect 12599 39389 12633 39423
rect 20913 39389 20947 39423
rect 21281 39389 21315 39423
rect 21741 39389 21775 39423
rect 22017 39389 22051 39423
rect 22293 39389 22327 39423
rect 22569 39389 22603 39423
rect 23029 39389 23063 39423
rect 23397 39389 23431 39423
rect 23857 39389 23891 39423
rect 23949 39389 23983 39423
rect 1501 39321 1535 39355
rect 1685 39321 1719 39355
rect 2329 39321 2363 39355
rect 2697 39321 2731 39355
rect 4261 39321 4295 39355
rect 4721 39321 4755 39355
rect 1961 39253 1995 39287
rect 3065 39253 3099 39287
rect 3249 39253 3283 39287
rect 3985 39253 4019 39287
rect 5089 39253 5123 39287
rect 5273 39253 5307 39287
rect 7297 39253 7331 39287
rect 21097 39253 21131 39287
rect 22845 39253 22879 39287
rect 23213 39253 23247 39287
rect 23673 39253 23707 39287
rect 24133 39253 24167 39287
rect 20453 39049 20487 39083
rect 20729 39049 20763 39083
rect 23397 39049 23431 39083
rect 23673 39049 23707 39083
rect 24133 38981 24167 39015
rect 1959 38913 1993 38947
rect 3065 38913 3099 38947
rect 4077 38913 4111 38947
rect 4629 38913 4663 38947
rect 8367 38913 8401 38947
rect 11771 38913 11805 38947
rect 20637 38913 20671 38947
rect 20913 38913 20947 38947
rect 21649 38913 21683 38947
rect 22089 38913 22123 38947
rect 23581 38913 23615 38947
rect 23857 38913 23891 38947
rect 1685 38845 1719 38879
rect 3801 38845 3835 38879
rect 4353 38845 4387 38879
rect 4905 38845 4939 38879
rect 8125 38845 8159 38879
rect 11529 38845 11563 38879
rect 21833 38845 21867 38879
rect 2697 38709 2731 38743
rect 9137 38709 9171 38743
rect 12541 38709 12575 38743
rect 21465 38709 21499 38743
rect 23213 38709 23247 38743
rect 24409 38709 24443 38743
rect 13277 38505 13311 38539
rect 19901 38505 19935 38539
rect 22477 38505 22511 38539
rect 23673 38505 23707 38539
rect 6009 38437 6043 38471
rect 12081 38437 12115 38471
rect 23029 38437 23063 38471
rect 6402 38369 6436 38403
rect 12357 38369 12391 38403
rect 3801 38301 3835 38335
rect 4059 38271 4093 38305
rect 5365 38301 5399 38335
rect 5549 38301 5583 38335
rect 6285 38301 6319 38335
rect 6561 38301 6595 38335
rect 9137 38301 9171 38335
rect 9395 38271 9429 38305
rect 11437 38301 11471 38335
rect 11621 38301 11655 38335
rect 12474 38301 12508 38335
rect 12633 38301 12667 38335
rect 20085 38301 20119 38335
rect 22109 38301 22143 38335
rect 22661 38301 22695 38335
rect 22753 38301 22787 38335
rect 22937 38301 22971 38335
rect 23213 38301 23247 38335
rect 23489 38301 23523 38335
rect 23857 38301 23891 38335
rect 23949 38301 23983 38335
rect 1409 38233 1443 38267
rect 2237 38233 2271 38267
rect 2421 38233 2455 38267
rect 3157 38233 3191 38267
rect 4813 38165 4847 38199
rect 7205 38165 7239 38199
rect 10149 38165 10183 38199
rect 22201 38165 22235 38199
rect 22937 38165 22971 38199
rect 23305 38165 23339 38199
rect 24133 38165 24167 38199
rect 7389 37961 7423 37995
rect 13093 37961 13127 37995
rect 23857 37961 23891 37995
rect 3525 37893 3559 37927
rect 3893 37893 3927 37927
rect 4629 37893 4663 37927
rect 5825 37893 5859 37927
rect 8953 37893 8987 37927
rect 9229 37893 9263 37927
rect 9321 37893 9355 37927
rect 10057 37893 10091 37927
rect 23765 37893 23799 37927
rect 1409 37825 1443 37859
rect 2203 37825 2237 37859
rect 3801 37825 3835 37859
rect 4261 37825 4295 37859
rect 4997 37825 5031 37859
rect 5549 37825 5583 37859
rect 6651 37825 6685 37859
rect 9689 37825 9723 37859
rect 12355 37825 12389 37859
rect 21649 37825 21683 37859
rect 22107 37825 22141 37859
rect 23397 37825 23431 37859
rect 24041 37825 24075 37859
rect 24225 37825 24259 37859
rect 1685 37757 1719 37791
rect 1961 37757 1995 37791
rect 5273 37757 5307 37791
rect 6377 37757 6411 37791
rect 12081 37757 12115 37791
rect 21833 37757 21867 37791
rect 23213 37757 23247 37791
rect 2973 37689 3007 37723
rect 4813 37689 4847 37723
rect 21465 37689 21499 37723
rect 22845 37689 22879 37723
rect 23673 37689 23707 37723
rect 10241 37621 10275 37655
rect 24409 37621 24443 37655
rect 3433 37417 3467 37451
rect 22569 37417 22603 37451
rect 22845 37417 22879 37451
rect 21925 37349 21959 37383
rect 8217 37281 8251 37315
rect 8401 37281 8435 37315
rect 10057 37281 10091 37315
rect 24133 37281 24167 37315
rect 2513 37213 2547 37247
rect 3801 37213 3835 37247
rect 4721 37213 4755 37247
rect 4995 37213 5029 37247
rect 6561 37213 6595 37247
rect 6819 37183 6853 37217
rect 7941 37213 7975 37247
rect 8033 37213 8067 37247
rect 8309 37213 8343 37247
rect 8493 37213 8527 37247
rect 10331 37213 10365 37247
rect 20729 37213 20763 37247
rect 21833 37213 21867 37247
rect 22109 37213 22143 37247
rect 22753 37213 22787 37247
rect 23029 37213 23063 37247
rect 23305 37213 23339 37247
rect 23581 37213 23615 37247
rect 1409 37145 1443 37179
rect 2237 37145 2271 37179
rect 2789 37145 2823 37179
rect 3157 37145 3191 37179
rect 4077 37145 4111 37179
rect 23857 37145 23891 37179
rect 5733 37077 5767 37111
rect 7573 37077 7607 37111
rect 8217 37077 8251 37111
rect 11069 37077 11103 37111
rect 20545 37077 20579 37111
rect 21649 37077 21683 37111
rect 23121 37077 23155 37111
rect 23397 37077 23431 37111
rect 5917 36873 5951 36907
rect 7205 36873 7239 36907
rect 20361 36873 20395 36907
rect 20913 36873 20947 36907
rect 23949 36873 23983 36907
rect 1593 36805 1627 36839
rect 3433 36805 3467 36839
rect 3801 36805 3835 36839
rect 4537 36805 4571 36839
rect 23673 36805 23707 36839
rect 2143 36737 2177 36771
rect 3709 36737 3743 36771
rect 4169 36737 4203 36771
rect 5163 36737 5197 36771
rect 6929 36737 6963 36771
rect 7021 36737 7055 36771
rect 7389 36737 7423 36771
rect 7755 36737 7789 36771
rect 11771 36737 11805 36771
rect 17785 36737 17819 36771
rect 19165 36737 19199 36771
rect 19809 36737 19843 36771
rect 20269 36737 20303 36771
rect 20545 36737 20579 36771
rect 20821 36737 20855 36771
rect 21097 36737 21131 36771
rect 23029 36737 23063 36771
rect 23305 36737 23339 36771
rect 24133 36737 24167 36771
rect 24225 36737 24259 36771
rect 1869 36669 1903 36703
rect 4905 36669 4939 36703
rect 7481 36669 7515 36703
rect 11529 36669 11563 36703
rect 2881 36601 2915 36635
rect 18981 36601 19015 36635
rect 20085 36601 20119 36635
rect 20637 36601 20671 36635
rect 23121 36601 23155 36635
rect 1685 36533 1719 36567
rect 4721 36533 4755 36567
rect 8493 36533 8527 36567
rect 12541 36533 12575 36567
rect 17601 36533 17635 36567
rect 19625 36533 19659 36567
rect 22845 36533 22879 36567
rect 24409 36533 24443 36567
rect 7021 36329 7055 36363
rect 22385 36329 22419 36363
rect 23397 36329 23431 36363
rect 5733 36261 5767 36295
rect 10977 36261 11011 36295
rect 18521 36261 18555 36295
rect 21005 36261 21039 36295
rect 4721 36193 4755 36227
rect 6929 36193 6963 36227
rect 11253 36193 11287 36227
rect 1501 36125 1535 36159
rect 1775 36125 1809 36159
rect 2881 36125 2915 36159
rect 3801 36125 3835 36159
rect 5089 36125 5123 36159
rect 5273 36125 5307 36159
rect 6009 36125 6043 36159
rect 6126 36125 6160 36159
rect 6285 36125 6319 36159
rect 7205 36125 7239 36159
rect 8953 36125 8987 36159
rect 9227 36125 9261 36159
rect 10333 36125 10367 36159
rect 10517 36125 10551 36159
rect 11370 36125 11404 36159
rect 11539 36125 11573 36159
rect 17141 36125 17175 36159
rect 18797 36125 18831 36159
rect 21189 36125 21223 36159
rect 21833 36125 21867 36159
rect 22569 36125 22603 36159
rect 23581 36125 23615 36159
rect 23857 36125 23891 36159
rect 3157 36057 3191 36091
rect 4077 36057 4111 36091
rect 4445 36057 4479 36091
rect 12173 36057 12207 36091
rect 17386 36057 17420 36091
rect 24225 36057 24259 36091
rect 2513 35989 2547 36023
rect 9965 35989 9999 36023
rect 18613 35989 18647 36023
rect 21649 35989 21683 36023
rect 3341 35785 3375 35819
rect 6193 35785 6227 35819
rect 8217 35785 8251 35819
rect 14197 35785 14231 35819
rect 21097 35785 21131 35819
rect 21833 35785 21867 35819
rect 23121 35785 23155 35819
rect 23489 35785 23523 35819
rect 8585 35717 8619 35751
rect 9321 35717 9355 35751
rect 11713 35717 11747 35751
rect 11989 35717 12023 35751
rect 12081 35717 12115 35751
rect 12817 35717 12851 35751
rect 1501 35649 1535 35683
rect 2697 35649 2731 35683
rect 3433 35649 3467 35683
rect 8493 35649 8527 35683
rect 8953 35649 8987 35683
rect 9947 35679 9981 35713
rect 12449 35649 12483 35683
rect 13459 35649 13493 35683
rect 17843 35649 17877 35683
rect 18981 35649 19015 35683
rect 19349 35649 19383 35683
rect 19533 35649 19567 35683
rect 21281 35649 21315 35683
rect 22017 35649 22051 35683
rect 22569 35649 22603 35683
rect 22845 35649 22879 35683
rect 23305 35649 23339 35683
rect 23673 35649 23707 35683
rect 23949 35649 23983 35683
rect 24133 35649 24167 35683
rect 1685 35581 1719 35615
rect 2421 35581 2455 35615
rect 2559 35581 2593 35615
rect 3617 35581 3651 35615
rect 4353 35581 4387 35615
rect 4537 35581 4571 35615
rect 5273 35581 5307 35615
rect 5411 35581 5445 35615
rect 5549 35581 5583 35615
rect 9689 35581 9723 35615
rect 13185 35581 13219 35615
rect 17601 35581 17635 35615
rect 19257 35581 19291 35615
rect 19441 35581 19475 35615
rect 2145 35513 2179 35547
rect 4997 35513 5031 35547
rect 13001 35513 13035 35547
rect 18613 35513 18647 35547
rect 22661 35513 22695 35547
rect 9505 35445 9539 35479
rect 10701 35445 10735 35479
rect 19073 35445 19107 35479
rect 19165 35445 19199 35479
rect 22385 35445 22419 35479
rect 23765 35445 23799 35479
rect 24409 35445 24443 35479
rect 5273 35241 5307 35275
rect 6469 35241 6503 35275
rect 11713 35241 11747 35275
rect 12817 35241 12851 35275
rect 18245 35241 18279 35275
rect 23213 35241 23247 35275
rect 3341 35173 3375 35207
rect 16681 35173 16715 35207
rect 20821 35173 20855 35207
rect 1685 35105 1719 35139
rect 5457 35105 5491 35139
rect 10057 35105 10091 35139
rect 10517 35105 10551 35139
rect 10931 35105 10965 35139
rect 15669 35105 15703 35139
rect 1409 35037 1443 35071
rect 2329 35037 2363 35071
rect 2603 35037 2637 35071
rect 4261 35037 4295 35071
rect 5731 35037 5765 35071
rect 9873 35037 9907 35071
rect 10793 35037 10827 35071
rect 11069 35037 11103 35071
rect 11805 35037 11839 35071
rect 12079 35037 12113 35071
rect 14105 35037 14139 35071
rect 14379 35037 14413 35071
rect 15927 35007 15961 35041
rect 18153 35037 18187 35071
rect 19717 35037 19751 35071
rect 20085 35037 20119 35071
rect 21005 35037 21039 35071
rect 23397 35037 23431 35071
rect 23673 35037 23707 35071
rect 23949 35037 23983 35071
rect 4353 34969 4387 35003
rect 4721 34969 4755 35003
rect 3985 34901 4019 34935
rect 5089 34901 5123 34935
rect 15117 34901 15151 34935
rect 19533 34901 19567 34935
rect 19901 34901 19935 34935
rect 23489 34901 23523 34935
rect 24133 34901 24167 34935
rect 2421 34697 2455 34731
rect 4537 34697 4571 34731
rect 9045 34697 9079 34731
rect 15209 34697 15243 34731
rect 16957 34697 16991 34731
rect 18797 34697 18831 34731
rect 21465 34697 21499 34731
rect 23673 34697 23707 34731
rect 3065 34629 3099 34663
rect 19340 34629 19374 34663
rect 24133 34629 24167 34663
rect 1683 34561 1717 34595
rect 2789 34561 2823 34595
rect 3525 34561 3559 34595
rect 3799 34561 3833 34595
rect 4905 34561 4939 34595
rect 6619 34561 6653 34595
rect 8769 34561 8803 34595
rect 9321 34561 9355 34595
rect 9505 34561 9539 34595
rect 9597 34561 9631 34595
rect 10057 34561 10091 34595
rect 10299 34561 10333 34595
rect 14471 34571 14505 34605
rect 16682 34583 16716 34617
rect 17049 34561 17083 34595
rect 17325 34561 17359 34595
rect 17509 34561 17543 34595
rect 18981 34561 19015 34595
rect 20545 34561 20579 34595
rect 21005 34561 21039 34595
rect 21649 34561 21683 34595
rect 22091 34591 22125 34625
rect 23397 34561 23431 34595
rect 23857 34561 23891 34595
rect 1409 34493 1443 34527
rect 5089 34493 5123 34527
rect 6377 34493 6411 34527
rect 9045 34493 9079 34527
rect 14197 34493 14231 34527
rect 16957 34493 16991 34527
rect 17417 34493 17451 34527
rect 19073 34493 19107 34527
rect 20637 34493 20671 34527
rect 21833 34493 21867 34527
rect 24409 34493 24443 34527
rect 8861 34425 8895 34459
rect 9689 34425 9723 34459
rect 16773 34425 16807 34459
rect 17141 34425 17175 34459
rect 23213 34425 23247 34459
rect 7389 34357 7423 34391
rect 9413 34357 9447 34391
rect 11069 34357 11103 34391
rect 20453 34357 20487 34391
rect 20821 34357 20855 34391
rect 22845 34357 22879 34391
rect 9965 34153 9999 34187
rect 17325 34153 17359 34187
rect 21097 34153 21131 34187
rect 22385 34153 22419 34187
rect 7481 34085 7515 34119
rect 13553 34085 13587 34119
rect 17693 34085 17727 34119
rect 20637 34085 20671 34119
rect 23121 34085 23155 34119
rect 3065 34017 3099 34051
rect 6837 34017 6871 34051
rect 7021 34017 7055 34051
rect 7757 34017 7791 34051
rect 8953 34017 8987 34051
rect 12541 34017 12575 34051
rect 15945 34017 15979 34051
rect 21281 34017 21315 34051
rect 21465 34017 21499 34051
rect 1409 33949 1443 33983
rect 1683 33949 1717 33983
rect 2789 33949 2823 33983
rect 3801 33949 3835 33983
rect 4537 33949 4571 33983
rect 4779 33949 4813 33983
rect 7895 33949 7929 33983
rect 8033 33949 8067 33983
rect 9195 33949 9229 33983
rect 12815 33949 12849 33983
rect 14105 33949 14139 33983
rect 14363 33949 14397 33983
rect 16219 33949 16253 33983
rect 17509 33949 17543 33983
rect 17877 33949 17911 33983
rect 18153 33949 18187 33983
rect 19625 33949 19659 33983
rect 19899 33949 19933 33983
rect 21005 33949 21039 33983
rect 21373 33949 21407 33983
rect 21557 33949 21591 33983
rect 22569 33949 22603 33983
rect 22845 33949 22879 33983
rect 23305 33949 23339 33983
rect 23581 33949 23615 33983
rect 23857 33949 23891 33983
rect 23949 33949 23983 33983
rect 4077 33881 4111 33915
rect 2421 33813 2455 33847
rect 5549 33813 5583 33847
rect 8677 33813 8711 33847
rect 15117 33813 15151 33847
rect 16957 33813 16991 33847
rect 18245 33813 18279 33847
rect 21281 33813 21315 33847
rect 22661 33813 22695 33847
rect 23397 33813 23431 33847
rect 23673 33813 23707 33847
rect 24133 33813 24167 33847
rect 8861 33609 8895 33643
rect 9137 33609 9171 33643
rect 16957 33609 16991 33643
rect 18613 33609 18647 33643
rect 23213 33609 23247 33643
rect 3065 33541 3099 33575
rect 3341 33541 3375 33575
rect 4169 33541 4203 33575
rect 18981 33541 19015 33575
rect 24133 33541 24167 33575
rect 1759 33473 1793 33507
rect 3433 33473 3467 33507
rect 3801 33473 3835 33507
rect 4905 33473 4939 33507
rect 5163 33503 5197 33537
rect 8125 33473 8159 33507
rect 9045 33473 9079 33507
rect 9321 33473 9355 33507
rect 9763 33473 9797 33507
rect 11989 33473 12023 33507
rect 12725 33473 12759 33507
rect 15209 33473 15243 33507
rect 15467 33473 15501 33507
rect 17141 33473 17175 33507
rect 17233 33473 17267 33507
rect 17489 33473 17523 33507
rect 18705 33473 18739 33507
rect 18797 33473 18831 33507
rect 19073 33473 19107 33507
rect 19257 33473 19291 33507
rect 19533 33473 19567 33507
rect 21649 33473 21683 33507
rect 22089 33473 22123 33507
rect 23305 33473 23339 33507
rect 23673 33473 23707 33507
rect 23857 33473 23891 33507
rect 1501 33405 1535 33439
rect 6929 33405 6963 33439
rect 7113 33405 7147 33439
rect 7849 33405 7883 33439
rect 7966 33405 8000 33439
rect 8769 33405 8803 33439
rect 9505 33405 9539 33439
rect 11805 33405 11839 33439
rect 12842 33405 12876 33439
rect 13001 33405 13035 33439
rect 18981 33405 19015 33439
rect 21833 33405 21867 33439
rect 23581 33405 23615 33439
rect 23765 33405 23799 33439
rect 2513 33337 2547 33371
rect 4353 33337 4387 33371
rect 7573 33337 7607 33371
rect 12449 33337 12483 33371
rect 19165 33337 19199 33371
rect 19349 33337 19383 33371
rect 5917 33269 5951 33303
rect 10517 33269 10551 33303
rect 13645 33269 13679 33303
rect 16221 33269 16255 33303
rect 21465 33269 21499 33303
rect 23397 33269 23431 33303
rect 23489 33269 23523 33303
rect 24409 33269 24443 33303
rect 3341 33065 3375 33099
rect 8217 33065 8251 33099
rect 11805 33065 11839 33099
rect 12909 33065 12943 33099
rect 15945 33065 15979 33099
rect 18613 33065 18647 33099
rect 22293 33065 22327 33099
rect 14749 32997 14783 33031
rect 21925 32997 21959 33031
rect 23673 32997 23707 33031
rect 2329 32929 2363 32963
rect 7205 32929 7239 32963
rect 10149 32929 10183 32963
rect 10609 32929 10643 32963
rect 10885 32929 10919 32963
rect 11023 32929 11057 32963
rect 11897 32929 11931 32963
rect 17601 32929 17635 32963
rect 1409 32861 1443 32895
rect 2603 32861 2637 32895
rect 5273 32861 5307 32895
rect 5365 32861 5399 32895
rect 5733 32861 5767 32895
rect 7479 32861 7513 32895
rect 9965 32861 9999 32895
rect 11161 32861 11195 32895
rect 12171 32861 12205 32895
rect 14105 32861 14139 32895
rect 14289 32861 14323 32895
rect 15025 32861 15059 32895
rect 15142 32861 15176 32895
rect 15301 32861 15335 32895
rect 17843 32861 17877 32895
rect 22109 32861 22143 32895
rect 22201 32861 22235 32895
rect 23029 32861 23063 32895
rect 23581 32861 23615 32895
rect 23857 32861 23891 32895
rect 23949 32861 23983 32895
rect 1685 32793 1719 32827
rect 3801 32793 3835 32827
rect 4537 32793 4571 32827
rect 4997 32725 5031 32759
rect 6101 32725 6135 32759
rect 6285 32725 6319 32759
rect 22845 32725 22879 32759
rect 23397 32725 23431 32759
rect 24133 32725 24167 32759
rect 11069 32521 11103 32555
rect 15209 32521 15243 32555
rect 15393 32521 15427 32555
rect 22661 32521 22695 32555
rect 23673 32521 23707 32555
rect 3249 32453 3283 32487
rect 14105 32453 14139 32487
rect 14381 32453 14415 32487
rect 14473 32453 14507 32487
rect 2329 32385 2363 32419
rect 2446 32385 2480 32419
rect 2603 32385 2637 32419
rect 3341 32385 3375 32419
rect 3893 32385 3927 32419
rect 4629 32385 4663 32419
rect 8033 32385 8067 32419
rect 8307 32385 8341 32419
rect 10057 32385 10091 32419
rect 10331 32385 10365 32419
rect 14841 32385 14875 32419
rect 19165 32385 19199 32419
rect 19432 32385 19466 32419
rect 22017 32385 22051 32419
rect 22569 32385 22603 32419
rect 22845 32385 22879 32419
rect 23305 32385 23339 32419
rect 23581 32385 23615 32419
rect 23857 32385 23891 32419
rect 24133 32385 24167 32419
rect 24225 32385 24259 32419
rect 1409 32317 1443 32351
rect 1593 32317 1627 32351
rect 2053 32317 2087 32351
rect 3617 32317 3651 32351
rect 4077 32317 4111 32351
rect 21833 32249 21867 32283
rect 23397 32249 23431 32283
rect 9045 32181 9079 32215
rect 20545 32181 20579 32215
rect 22385 32181 22419 32215
rect 23121 32181 23155 32215
rect 23949 32181 23983 32215
rect 24409 32181 24443 32215
rect 2421 31977 2455 32011
rect 4721 31977 4755 32011
rect 15117 31977 15151 32011
rect 21649 31977 21683 32011
rect 23489 31977 23523 32011
rect 6837 31909 6871 31943
rect 16221 31909 16255 31943
rect 19533 31909 19567 31943
rect 20637 31909 20671 31943
rect 20913 31909 20947 31943
rect 21189 31909 21223 31943
rect 3065 31841 3099 31875
rect 3985 31841 4019 31875
rect 5825 31841 5859 31875
rect 11069 31841 11103 31875
rect 14105 31841 14139 31875
rect 16614 31841 16648 31875
rect 16773 31841 16807 31875
rect 17417 31841 17451 31875
rect 1409 31773 1443 31807
rect 1667 31743 1701 31777
rect 2789 31773 2823 31807
rect 3801 31773 3835 31807
rect 4905 31773 4939 31807
rect 6083 31743 6117 31777
rect 11343 31773 11377 31807
rect 13093 31773 13127 31807
rect 13185 31773 13219 31807
rect 14379 31773 14413 31807
rect 15577 31773 15611 31807
rect 15761 31773 15795 31807
rect 16497 31773 16531 31807
rect 19717 31773 19751 31807
rect 20085 31773 20119 31807
rect 20177 31773 20211 31807
rect 20821 31773 20855 31807
rect 21097 31773 21131 31807
rect 21373 31773 21407 31807
rect 21833 31773 21867 31807
rect 23213 31773 23247 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24225 31773 24259 31807
rect 12081 31637 12115 31671
rect 3893 31433 3927 31467
rect 7665 31433 7699 31467
rect 8677 31433 8711 31467
rect 4169 31365 4203 31399
rect 4445 31365 4479 31399
rect 4537 31365 4571 31399
rect 5273 31365 5307 31399
rect 6561 31365 6595 31399
rect 7297 31365 7331 31399
rect 8953 31365 8987 31399
rect 11621 31365 11655 31399
rect 12265 31365 12299 31399
rect 1683 31307 1717 31341
rect 3709 31297 3743 31331
rect 4905 31297 4939 31331
rect 6837 31297 6871 31331
rect 6929 31297 6963 31331
rect 9045 31297 9079 31331
rect 9413 31297 9447 31331
rect 9795 31297 9829 31331
rect 12541 31297 12575 31331
rect 12815 31297 12849 31331
rect 13921 31297 13955 31331
rect 14105 31297 14139 31331
rect 15391 31297 15425 31331
rect 16923 31297 16957 31331
rect 18245 31297 18279 31331
rect 18521 31297 18555 31331
rect 19775 31297 19809 31331
rect 21097 31297 21131 31331
rect 21465 31297 21499 31331
rect 22477 31297 22511 31331
rect 23121 31297 23155 31331
rect 23765 31297 23799 31331
rect 24133 31297 24167 31331
rect 24225 31297 24259 31331
rect 1409 31229 1443 31263
rect 2789 31229 2823 31263
rect 3065 31229 3099 31263
rect 15117 31229 15151 31263
rect 16681 31229 16715 31263
rect 19533 31229 19567 31263
rect 20913 31229 20947 31263
rect 12449 31161 12483 31195
rect 13553 31161 13587 31195
rect 18061 31161 18095 31195
rect 20545 31161 20579 31195
rect 21097 31161 21131 31195
rect 22293 31161 22327 31195
rect 22937 31161 22971 31195
rect 23581 31161 23615 31195
rect 2421 31093 2455 31127
rect 5457 31093 5491 31127
rect 7849 31093 7883 31127
rect 9965 31093 9999 31127
rect 11713 31093 11747 31127
rect 14013 31093 14047 31127
rect 16129 31093 16163 31127
rect 17693 31093 17727 31127
rect 18613 31093 18647 31127
rect 23949 31093 23983 31127
rect 24409 31093 24443 31127
rect 3341 30889 3375 30923
rect 5273 30889 5307 30923
rect 7389 30889 7423 30923
rect 9965 30889 9999 30923
rect 12541 30889 12575 30923
rect 12817 30889 12851 30923
rect 17601 30889 17635 30923
rect 19349 30889 19383 30923
rect 20729 30889 20763 30923
rect 23121 30889 23155 30923
rect 16405 30821 16439 30855
rect 19073 30821 19107 30855
rect 19901 30821 19935 30855
rect 22845 30821 22879 30855
rect 23489 30821 23523 30855
rect 2329 30753 2363 30787
rect 4261 30753 4295 30787
rect 6377 30753 6411 30787
rect 8953 30753 8987 30787
rect 11161 30753 11195 30787
rect 11437 30753 11471 30787
rect 11554 30753 11588 30787
rect 11713 30753 11747 30787
rect 16798 30753 16832 30787
rect 16957 30753 16991 30787
rect 17693 30753 17727 30787
rect 19533 30753 19567 30787
rect 19717 30753 19751 30787
rect 2603 30685 2637 30719
rect 3801 30685 3835 30719
rect 4535 30685 4569 30719
rect 6651 30685 6685 30719
rect 9227 30685 9261 30719
rect 10517 30685 10551 30719
rect 10701 30685 10735 30719
rect 12357 30685 12391 30719
rect 12725 30685 12759 30719
rect 13001 30685 13035 30719
rect 14105 30685 14139 30719
rect 14473 30685 14507 30719
rect 14933 30685 14967 30719
rect 15761 30685 15795 30719
rect 15945 30685 15979 30719
rect 16681 30685 16715 30719
rect 17949 30685 17983 30719
rect 19257 30685 19291 30719
rect 19625 30685 19659 30719
rect 19809 30685 19843 30719
rect 20085 30685 20119 30719
rect 20637 30685 20671 30719
rect 20821 30685 20855 30719
rect 22293 30685 22327 30719
rect 23029 30685 23063 30719
rect 23305 30685 23339 30719
rect 23673 30685 23707 30719
rect 1501 30617 1535 30651
rect 1685 30617 1719 30651
rect 15209 30617 15243 30651
rect 19533 30617 19567 30651
rect 23857 30617 23891 30651
rect 24225 30617 24259 30651
rect 3985 30549 4019 30583
rect 22109 30549 22143 30583
rect 10977 30345 11011 30379
rect 18981 30345 19015 30379
rect 23765 30345 23799 30379
rect 3341 30277 3375 30311
rect 24133 30277 24167 30311
rect 2697 30209 2731 30243
rect 3433 30209 3467 30243
rect 4427 30239 4461 30273
rect 7111 30209 7145 30243
rect 10239 30209 10273 30243
rect 14195 30209 14229 30243
rect 18243 30209 18277 30243
rect 20525 30209 20559 30243
rect 22107 30209 22141 30243
rect 23397 30209 23431 30243
rect 23673 30209 23707 30243
rect 23949 30209 23983 30243
rect 1501 30141 1535 30175
rect 1685 30141 1719 30175
rect 2145 30141 2179 30175
rect 2421 30141 2455 30175
rect 2559 30141 2593 30175
rect 4169 30141 4203 30175
rect 6837 30141 6871 30175
rect 9965 30141 9999 30175
rect 13921 30141 13955 30175
rect 17969 30141 18003 30175
rect 20269 30141 20303 30175
rect 21833 30141 21867 30175
rect 23489 30073 23523 30107
rect 3617 30005 3651 30039
rect 5181 30005 5215 30039
rect 7849 30005 7883 30039
rect 14933 30005 14967 30039
rect 21649 30005 21683 30039
rect 22845 30005 22879 30039
rect 23213 30005 23247 30039
rect 24409 30005 24443 30039
rect 2697 29801 2731 29835
rect 3249 29801 3283 29835
rect 3617 29801 3651 29835
rect 6285 29801 6319 29835
rect 8769 29801 8803 29835
rect 17417 29801 17451 29835
rect 1593 29733 1627 29767
rect 7573 29733 7607 29767
rect 11161 29733 11195 29767
rect 16221 29733 16255 29767
rect 23305 29733 23339 29767
rect 23581 29733 23615 29767
rect 3801 29665 3835 29699
rect 11437 29665 11471 29699
rect 11575 29665 11609 29699
rect 11713 29665 11747 29699
rect 12357 29665 12391 29699
rect 14197 29665 14231 29699
rect 15761 29665 15795 29699
rect 16497 29665 16531 29699
rect 16773 29665 16807 29699
rect 21741 29665 21775 29699
rect 22109 29665 22143 29699
rect 22293 29665 22327 29699
rect 22477 29665 22511 29699
rect 1409 29597 1443 29631
rect 1685 29597 1719 29631
rect 1959 29597 1993 29631
rect 3065 29597 3099 29631
rect 3433 29597 3467 29631
rect 4077 29597 4111 29631
rect 6929 29597 6963 29631
rect 7113 29597 7147 29631
rect 7849 29597 7883 29631
rect 7966 29597 8000 29631
rect 8125 29597 8159 29631
rect 10517 29597 10551 29631
rect 10701 29597 10735 29631
rect 12449 29597 12483 29631
rect 12691 29587 12725 29621
rect 14471 29597 14505 29631
rect 15577 29597 15611 29631
rect 16614 29597 16648 29631
rect 21189 29597 21223 29631
rect 21649 29597 21683 29631
rect 22017 29597 22051 29631
rect 22385 29597 22419 29631
rect 22569 29597 22603 29631
rect 23497 29597 23531 29631
rect 23765 29597 23799 29631
rect 23949 29597 23983 29631
rect 5273 29529 5307 29563
rect 5365 29529 5399 29563
rect 5733 29529 5767 29563
rect 22293 29529 22327 29563
rect 4997 29461 5031 29495
rect 6101 29461 6135 29495
rect 13461 29461 13495 29495
rect 15209 29461 15243 29495
rect 21005 29461 21039 29495
rect 24133 29461 24167 29495
rect 1593 29257 1627 29291
rect 3801 29257 3835 29291
rect 5917 29257 5951 29291
rect 8401 29257 8435 29291
rect 10885 29257 10919 29291
rect 14289 29257 14323 29291
rect 23121 29257 23155 29291
rect 1869 29189 1903 29223
rect 11621 29189 11655 29223
rect 14565 29189 14599 29223
rect 14657 29189 14691 29223
rect 15025 29189 15059 29223
rect 15393 29189 15427 29223
rect 1501 29121 1535 29155
rect 2511 29121 2545 29155
rect 3617 29121 3651 29155
rect 4905 29121 4939 29155
rect 5179 29121 5213 29155
rect 7663 29121 7697 29155
rect 9229 29121 9263 29155
rect 9503 29121 9537 29155
rect 10609 29121 10643 29155
rect 12541 29121 12575 29155
rect 12815 29121 12849 29155
rect 16955 29121 16989 29155
rect 19163 29121 19197 29155
rect 20269 29121 20303 29155
rect 20453 29121 20487 29155
rect 23305 29121 23339 29155
rect 23581 29121 23615 29155
rect 23857 29121 23891 29155
rect 24133 29121 24167 29155
rect 2237 29053 2271 29087
rect 7389 29053 7423 29087
rect 10885 29053 10919 29087
rect 16681 29053 16715 29087
rect 18889 29053 18923 29087
rect 2053 28985 2087 29019
rect 10241 28985 10275 29019
rect 10701 28985 10735 29019
rect 11805 28985 11839 29019
rect 15577 28985 15611 29019
rect 23397 28985 23431 29019
rect 23673 28985 23707 29019
rect 24409 28985 24443 29019
rect 3249 28917 3283 28951
rect 13553 28917 13587 28951
rect 17693 28917 17727 28951
rect 19901 28917 19935 28951
rect 20361 28917 20395 28951
rect 11161 28713 11195 28747
rect 11437 28713 11471 28747
rect 18889 28713 18923 28747
rect 22661 28713 22695 28747
rect 10793 28645 10827 28679
rect 18429 28645 18463 28679
rect 23213 28645 23247 28679
rect 1685 28577 1719 28611
rect 2329 28577 2363 28611
rect 8953 28577 8987 28611
rect 16681 28577 16715 28611
rect 17233 28577 17267 28611
rect 19349 28577 19383 28611
rect 19717 28577 19751 28611
rect 19901 28577 19935 28611
rect 19993 28577 20027 28611
rect 1409 28509 1443 28543
rect 2587 28479 2621 28513
rect 3893 28509 3927 28543
rect 4167 28509 4201 28543
rect 9211 28479 9245 28513
rect 10701 28509 10735 28543
rect 10977 28509 11011 28543
rect 11069 28509 11103 28543
rect 11345 28509 11379 28543
rect 11529 28509 11563 28543
rect 11713 28509 11747 28543
rect 11987 28509 12021 28543
rect 14105 28509 14139 28543
rect 14379 28509 14413 28543
rect 16037 28509 16071 28543
rect 16221 28509 16255 28543
rect 16957 28509 16991 28543
rect 17095 28509 17129 28543
rect 17877 28509 17911 28543
rect 18613 28509 18647 28543
rect 19073 28509 19107 28543
rect 19257 28509 19291 28543
rect 19625 28509 19659 28543
rect 20267 28509 20301 28543
rect 22845 28509 22879 28543
rect 23397 28509 23431 28543
rect 23673 28509 23707 28543
rect 23949 28509 23983 28543
rect 19901 28441 19935 28475
rect 3341 28373 3375 28407
rect 4905 28373 4939 28407
rect 9965 28373 9999 28407
rect 10517 28373 10551 28407
rect 12725 28373 12759 28407
rect 15117 28373 15151 28407
rect 21005 28373 21039 28407
rect 23489 28373 23523 28407
rect 24133 28373 24167 28407
rect 2513 28169 2547 28203
rect 3893 28169 3927 28203
rect 4077 28169 4111 28203
rect 5825 28169 5859 28203
rect 16221 28169 16255 28203
rect 19257 28169 19291 28203
rect 22109 28169 22143 28203
rect 23489 28169 23523 28203
rect 2789 28101 2823 28135
rect 3157 28101 3191 28135
rect 4537 28101 4571 28135
rect 4813 28101 4847 28135
rect 4905 28101 4939 28135
rect 5641 28101 5675 28135
rect 1501 28033 1535 28067
rect 1777 28033 1811 28067
rect 2329 28033 2363 28067
rect 3065 28033 3099 28067
rect 3525 28033 3559 28067
rect 5273 28033 5307 28067
rect 6651 28033 6685 28067
rect 10331 28033 10365 28067
rect 14013 28033 14047 28067
rect 15451 28033 15485 28067
rect 18133 28033 18167 28067
rect 19441 28033 19475 28067
rect 19697 28033 19731 28067
rect 20913 28033 20947 28067
rect 21281 28033 21315 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22293 28033 22327 28067
rect 22845 28033 22879 28067
rect 23121 28033 23155 28067
rect 23397 28033 23431 28067
rect 23673 28033 23707 28067
rect 23949 28033 23983 28067
rect 24133 28033 24167 28067
rect 6377 27965 6411 27999
rect 10057 27965 10091 27999
rect 12817 27965 12851 27999
rect 13001 27965 13035 27999
rect 13737 27965 13771 27999
rect 13854 27965 13888 27999
rect 15209 27965 15243 27999
rect 17877 27965 17911 27999
rect 21189 27965 21223 27999
rect 21925 27965 21959 27999
rect 1685 27897 1719 27931
rect 13461 27897 13495 27931
rect 21005 27897 21039 27931
rect 21373 27897 21407 27931
rect 22937 27897 22971 27931
rect 23213 27897 23247 27931
rect 1961 27829 1995 27863
rect 7389 27829 7423 27863
rect 11069 27829 11103 27863
rect 14657 27829 14691 27863
rect 20821 27829 20855 27863
rect 21097 27829 21131 27863
rect 22661 27829 22695 27863
rect 23765 27829 23799 27863
rect 24409 27829 24443 27863
rect 20913 27625 20947 27659
rect 22569 27625 22603 27659
rect 23581 27625 23615 27659
rect 5825 27557 5859 27591
rect 19993 27557 20027 27591
rect 22753 27557 22787 27591
rect 23121 27557 23155 27591
rect 1409 27489 1443 27523
rect 8953 27489 8987 27523
rect 9137 27489 9171 27523
rect 9597 27489 9631 27523
rect 10011 27489 10045 27523
rect 10149 27489 10183 27523
rect 16221 27489 16255 27523
rect 17601 27489 17635 27523
rect 22937 27489 22971 27523
rect 23397 27489 23431 27523
rect 1651 27421 1685 27455
rect 2789 27421 2823 27455
rect 3065 27421 3099 27455
rect 4813 27421 4847 27455
rect 5087 27421 5121 27455
rect 6745 27421 6779 27455
rect 9873 27421 9907 27455
rect 11529 27421 11563 27455
rect 11787 27421 11821 27455
rect 15209 27421 15243 27455
rect 16495 27411 16529 27445
rect 17843 27421 17877 27455
rect 20177 27421 20211 27455
rect 21097 27421 21131 27455
rect 21189 27421 21223 27455
rect 22661 27421 22695 27455
rect 23029 27421 23063 27455
rect 23305 27421 23339 27455
rect 23489 27421 23523 27455
rect 23765 27421 23799 27455
rect 23949 27421 23983 27455
rect 6653 27353 6687 27387
rect 7113 27353 7147 27387
rect 7481 27353 7515 27387
rect 10793 27353 10827 27387
rect 21434 27353 21468 27387
rect 2421 27285 2455 27319
rect 2973 27285 3007 27319
rect 3249 27285 3283 27319
rect 6377 27285 6411 27319
rect 7665 27285 7699 27319
rect 12541 27285 12575 27319
rect 15025 27285 15059 27319
rect 17233 27285 17267 27319
rect 18613 27285 18647 27319
rect 22937 27285 22971 27319
rect 24133 27285 24167 27319
rect 8769 27081 8803 27115
rect 22845 27081 22879 27115
rect 23305 27081 23339 27115
rect 23949 27081 23983 27115
rect 2053 27013 2087 27047
rect 3157 27013 3191 27047
rect 14657 27013 14691 27047
rect 2329 26945 2363 26979
rect 2421 26945 2455 26979
rect 2789 26945 2823 26979
rect 3525 26945 3559 26979
rect 4537 26945 4571 26979
rect 4811 26955 4845 26989
rect 7757 26945 7791 26979
rect 8031 26945 8065 26979
rect 13001 26945 13035 26979
rect 13854 26945 13888 26979
rect 15023 26945 15057 26979
rect 16681 26945 16715 26979
rect 17877 26945 17911 26979
rect 22107 26945 22141 26979
rect 23489 26945 23523 26979
rect 23765 26945 23799 26979
rect 24133 26945 24167 26979
rect 24225 26945 24259 26979
rect 12817 26877 12851 26911
rect 13461 26877 13495 26911
rect 13737 26877 13771 26911
rect 14013 26877 14047 26911
rect 14749 26877 14783 26911
rect 16865 26877 16899 26911
rect 17325 26877 17359 26911
rect 17601 26877 17635 26911
rect 17739 26877 17773 26911
rect 21833 26877 21867 26911
rect 3341 26809 3375 26843
rect 3709 26809 3743 26843
rect 23581 26809 23615 26843
rect 5549 26741 5583 26775
rect 15761 26741 15795 26775
rect 18521 26741 18555 26775
rect 24409 26741 24443 26775
rect 2605 26537 2639 26571
rect 3249 26537 3283 26571
rect 3341 26537 3375 26571
rect 4261 26537 4295 26571
rect 11069 26537 11103 26571
rect 15945 26537 15979 26571
rect 22753 26537 22787 26571
rect 9873 26469 9907 26503
rect 12817 26469 12851 26503
rect 19073 26469 19107 26503
rect 6561 26401 6595 26435
rect 9229 26401 9263 26435
rect 10287 26401 10321 26435
rect 16313 26401 16347 26435
rect 1593 26333 1627 26367
rect 1867 26333 1901 26367
rect 3525 26333 3559 26367
rect 3801 26333 3835 26367
rect 4077 26333 4111 26367
rect 6835 26333 6869 26367
rect 9413 26333 9447 26367
rect 10149 26333 10183 26367
rect 10425 26333 10459 26367
rect 11805 26333 11839 26367
rect 14933 26333 14967 26367
rect 15191 26303 15225 26337
rect 16497 26333 16531 26367
rect 16865 26333 16899 26367
rect 17693 26333 17727 26367
rect 17960 26333 17994 26367
rect 19441 26333 19475 26367
rect 22937 26333 22971 26367
rect 23489 26333 23523 26367
rect 23673 26333 23707 26367
rect 23857 26333 23891 26367
rect 11529 26265 11563 26299
rect 11897 26265 11931 26299
rect 12265 26265 12299 26299
rect 16773 26265 16807 26299
rect 24225 26265 24259 26299
rect 3985 26197 4019 26231
rect 7573 26197 7607 26231
rect 12633 26197 12667 26231
rect 19257 26197 19291 26231
rect 23673 26197 23707 26231
rect 3065 25993 3099 26027
rect 3341 25993 3375 26027
rect 8217 25993 8251 26027
rect 10885 25993 10919 26027
rect 15669 25993 15703 26027
rect 16037 25993 16071 26027
rect 22385 25993 22419 26027
rect 23489 25993 23523 26027
rect 23949 25993 23983 26027
rect 7113 25925 7147 25959
rect 24133 25925 24167 25959
rect 1501 25857 1535 25891
rect 1775 25857 1809 25891
rect 2881 25857 2915 25891
rect 3157 25857 3191 25891
rect 3433 25857 3467 25891
rect 3707 25857 3741 25891
rect 4813 25857 4847 25891
rect 5087 25857 5121 25891
rect 6837 25857 6871 25891
rect 7389 25857 7423 25891
rect 7481 25857 7515 25891
rect 7849 25857 7883 25891
rect 10082 25857 10116 25891
rect 11529 25857 11563 25891
rect 11787 25887 11821 25921
rect 13277 25857 13311 25891
rect 14289 25857 14323 25891
rect 14933 25857 14967 25891
rect 15485 25857 15519 25891
rect 15577 25857 15611 25891
rect 15853 25857 15887 25891
rect 16037 25857 16071 25891
rect 18613 25857 18647 25891
rect 18871 25887 18905 25921
rect 19993 25857 20027 25891
rect 20361 25857 20395 25891
rect 20545 25857 20579 25891
rect 21373 25857 21407 25891
rect 21557 25857 21591 25891
rect 22569 25857 22603 25891
rect 23029 25857 23063 25891
rect 23673 25857 23707 25891
rect 23765 25857 23799 25891
rect 9045 25789 9079 25823
rect 9229 25789 9263 25823
rect 9965 25789 9999 25823
rect 10241 25789 10275 25823
rect 13093 25789 13127 25823
rect 13737 25789 13771 25823
rect 14013 25789 14047 25823
rect 14130 25789 14164 25823
rect 20269 25789 20303 25823
rect 20453 25789 20487 25823
rect 9689 25721 9723 25755
rect 15301 25721 15335 25755
rect 19625 25721 19659 25755
rect 20177 25721 20211 25755
rect 2513 25653 2547 25687
rect 4445 25653 4479 25687
rect 5825 25653 5859 25687
rect 8401 25653 8435 25687
rect 12541 25653 12575 25687
rect 20085 25653 20119 25687
rect 21465 25653 21499 25687
rect 23121 25653 23155 25687
rect 24409 25653 24443 25687
rect 8309 25449 8343 25483
rect 10517 25449 10551 25483
rect 19349 25449 19383 25483
rect 21373 25449 21407 25483
rect 23489 25449 23523 25483
rect 1593 25381 1627 25415
rect 3341 25381 3375 25415
rect 12725 25381 12759 25415
rect 19625 25381 19659 25415
rect 23213 25381 23247 25415
rect 2329 25313 2363 25347
rect 7297 25313 7331 25347
rect 9505 25313 9539 25347
rect 16681 25313 16715 25347
rect 17325 25313 17359 25347
rect 17718 25313 17752 25347
rect 17877 25313 17911 25347
rect 20361 25313 20395 25347
rect 21833 25313 21867 25347
rect 23673 25313 23707 25347
rect 1409 25245 1443 25279
rect 1685 25245 1719 25279
rect 2145 25245 2179 25279
rect 2603 25245 2637 25279
rect 4353 25245 4387 25279
rect 5457 25245 5491 25279
rect 5715 25215 5749 25249
rect 7571 25245 7605 25279
rect 9779 25245 9813 25279
rect 16865 25245 16899 25279
rect 17601 25245 17635 25279
rect 19257 25245 19291 25279
rect 19809 25245 19843 25279
rect 20635 25245 20669 25279
rect 23397 25245 23431 25279
rect 4261 25177 4295 25211
rect 4721 25177 4755 25211
rect 5089 25177 5123 25211
rect 11437 25177 11471 25211
rect 11713 25177 11747 25211
rect 11805 25177 11839 25211
rect 12173 25177 12207 25211
rect 12541 25177 12575 25211
rect 22100 25177 22134 25211
rect 23857 25177 23891 25211
rect 24225 25177 24259 25211
rect 1869 25109 1903 25143
rect 1961 25109 1995 25143
rect 3985 25109 4019 25143
rect 5273 25109 5307 25143
rect 6469 25109 6503 25143
rect 18521 25109 18555 25143
rect 23673 25109 23707 25143
rect 1869 24905 1903 24939
rect 2145 24905 2179 24939
rect 2881 24905 2915 24939
rect 3999 24905 4033 24939
rect 17693 24905 17727 24939
rect 21833 24905 21867 24939
rect 23489 24905 23523 24939
rect 3617 24837 3651 24871
rect 1409 24769 1443 24803
rect 1685 24769 1719 24803
rect 1961 24769 1995 24803
rect 2237 24769 2271 24803
rect 3157 24769 3191 24803
rect 3249 24769 3283 24803
rect 4353 24769 4387 24803
rect 4537 24769 4571 24803
rect 5273 24769 5307 24803
rect 8493 24769 8527 24803
rect 8767 24769 8801 24803
rect 12431 24799 12465 24833
rect 16923 24769 16957 24803
rect 18335 24769 18369 24803
rect 19901 24769 19935 24803
rect 20157 24769 20191 24803
rect 21373 24769 21407 24803
rect 22017 24769 22051 24803
rect 22719 24769 22753 24803
rect 24133 24769 24167 24803
rect 5390 24701 5424 24735
rect 5549 24701 5583 24735
rect 12173 24701 12207 24735
rect 16681 24701 16715 24735
rect 18061 24701 18095 24735
rect 21649 24701 21683 24735
rect 22477 24701 22511 24735
rect 1593 24633 1627 24667
rect 4169 24633 4203 24667
rect 4997 24633 5031 24667
rect 9505 24633 9539 24667
rect 21281 24633 21315 24667
rect 2421 24565 2455 24599
rect 6193 24565 6227 24599
rect 13185 24565 13219 24599
rect 19073 24565 19107 24599
rect 21465 24565 21499 24599
rect 21557 24565 21591 24599
rect 24409 24565 24443 24599
rect 17969 24361 18003 24395
rect 21005 24361 21039 24395
rect 23397 24361 23431 24395
rect 23857 24361 23891 24395
rect 5825 24293 5859 24327
rect 9965 24293 9999 24327
rect 5181 24225 5215 24259
rect 6101 24225 6135 24259
rect 6377 24225 6411 24259
rect 7021 24225 7055 24259
rect 10609 24225 10643 24259
rect 12633 24225 12667 24259
rect 15025 24225 15059 24259
rect 15669 24225 15703 24259
rect 16062 24225 16096 24259
rect 16221 24225 16255 24259
rect 1869 24157 1903 24191
rect 5365 24157 5399 24191
rect 6218 24157 6252 24191
rect 7297 24157 7331 24191
rect 7481 24157 7515 24191
rect 7941 24157 7975 24191
rect 8953 24157 8987 24191
rect 9227 24157 9261 24191
rect 10883 24157 10917 24191
rect 12891 24127 12925 24161
rect 15209 24157 15243 24191
rect 15945 24157 15979 24191
rect 16957 24157 16991 24191
rect 17231 24157 17265 24191
rect 19717 24157 19751 24191
rect 19809 24157 19843 24191
rect 19993 24157 20027 24191
rect 20545 24157 20579 24191
rect 20913 24157 20947 24191
rect 23581 24157 23615 24191
rect 23673 24157 23707 24191
rect 23949 24157 23983 24191
rect 1593 24089 1627 24123
rect 1961 24089 1995 24123
rect 2329 24089 2363 24123
rect 2697 24021 2731 24055
rect 2881 24021 2915 24055
rect 7113 24021 7147 24055
rect 7573 24021 7607 24055
rect 7757 24021 7791 24055
rect 11621 24021 11655 24055
rect 13645 24021 13679 24055
rect 16865 24021 16899 24055
rect 19533 24021 19567 24055
rect 19901 24021 19935 24055
rect 20361 24021 20395 24055
rect 24133 24021 24167 24055
rect 3525 23817 3559 23851
rect 4077 23817 4111 23851
rect 10149 23817 10183 23851
rect 15669 23817 15703 23851
rect 19257 23817 19291 23851
rect 22845 23817 22879 23851
rect 8861 23749 8895 23783
rect 9137 23749 9171 23783
rect 9597 23749 9631 23783
rect 9965 23749 9999 23783
rect 24133 23749 24167 23783
rect 2513 23681 2547 23715
rect 2787 23681 2821 23715
rect 3893 23681 3927 23715
rect 7203 23681 7237 23715
rect 8309 23681 8343 23715
rect 8493 23681 8527 23715
rect 9229 23681 9263 23715
rect 11897 23681 11931 23715
rect 12633 23681 12667 23715
rect 13670 23681 13704 23715
rect 13829 23681 13863 23715
rect 14931 23681 14965 23715
rect 16221 23681 16255 23715
rect 17877 23681 17911 23715
rect 18133 23681 18167 23715
rect 19349 23681 19383 23715
rect 19623 23681 19657 23715
rect 23029 23681 23063 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 23489 23681 23523 23715
rect 23949 23681 23983 23715
rect 1409 23613 1443 23647
rect 1685 23613 1719 23647
rect 6929 23613 6963 23647
rect 12817 23613 12851 23647
rect 13277 23613 13311 23647
rect 13553 23613 13587 23647
rect 14657 23613 14691 23647
rect 23765 23545 23799 23579
rect 7941 23477 7975 23511
rect 8401 23477 8435 23511
rect 12081 23477 12115 23511
rect 14473 23477 14507 23511
rect 20361 23477 20395 23511
rect 23305 23477 23339 23511
rect 23581 23477 23615 23511
rect 24409 23477 24443 23511
rect 2237 23273 2271 23307
rect 3341 23273 3375 23307
rect 4813 23273 4847 23307
rect 9965 23273 9999 23307
rect 23765 23273 23799 23307
rect 18429 23205 18463 23239
rect 2329 23137 2363 23171
rect 3801 23137 3835 23171
rect 7849 23137 7883 23171
rect 14105 23137 14139 23171
rect 19349 23137 19383 23171
rect 19717 23137 19751 23171
rect 19901 23137 19935 23171
rect 2053 23069 2087 23103
rect 2603 23069 2637 23103
rect 4059 23039 4093 23073
rect 8033 23069 8067 23103
rect 8493 23069 8527 23103
rect 8953 23069 8987 23103
rect 9227 23069 9261 23103
rect 10885 23069 10919 23103
rect 10977 23069 11011 23103
rect 14379 23069 14413 23103
rect 18613 23069 18647 23103
rect 19257 23069 19291 23103
rect 19625 23069 19659 23103
rect 20637 23069 20671 23103
rect 22109 23069 22143 23103
rect 22385 23069 22419 23103
rect 23949 23069 23983 23103
rect 8769 23001 8803 23035
rect 10609 23001 10643 23035
rect 11345 23001 11379 23035
rect 20882 23001 20916 23035
rect 22641 23001 22675 23035
rect 11713 22933 11747 22967
rect 11897 22933 11931 22967
rect 15117 22933 15151 22967
rect 19901 22933 19935 22967
rect 22017 22933 22051 22967
rect 22201 22933 22235 22967
rect 24133 22933 24167 22967
rect 3341 22729 3375 22763
rect 11069 22729 11103 22763
rect 21097 22729 21131 22763
rect 24225 22729 24259 22763
rect 1409 22593 1443 22627
rect 1683 22593 1717 22627
rect 2973 22593 3007 22627
rect 3157 22593 3191 22627
rect 4443 22593 4477 22627
rect 6651 22593 6685 22627
rect 10057 22593 10091 22627
rect 10315 22623 10349 22657
rect 16865 22593 16899 22627
rect 17739 22593 17773 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 21649 22593 21683 22627
rect 21833 22593 21867 22627
rect 22107 22603 22141 22637
rect 23213 22593 23247 22627
rect 23487 22593 23521 22627
rect 4169 22525 4203 22559
rect 6377 22525 6411 22559
rect 16681 22525 16715 22559
rect 17601 22525 17635 22559
rect 17877 22525 17911 22559
rect 17325 22457 17359 22491
rect 2421 22389 2455 22423
rect 5181 22389 5215 22423
rect 7389 22389 7423 22423
rect 14841 22389 14875 22423
rect 18521 22389 18555 22423
rect 21557 22389 21591 22423
rect 22845 22389 22879 22423
rect 3065 22185 3099 22219
rect 3985 22185 4019 22219
rect 11069 22185 11103 22219
rect 12909 22185 12943 22219
rect 17325 22185 17359 22219
rect 22109 22185 22143 22219
rect 23213 22185 23247 22219
rect 6009 22117 6043 22151
rect 6561 22117 6595 22151
rect 22385 22117 22419 22151
rect 6653 22049 6687 22083
rect 10057 22049 10091 22083
rect 14749 22049 14783 22083
rect 15025 22049 15059 22083
rect 15301 22049 15335 22083
rect 19257 22049 19291 22083
rect 22293 22049 22327 22083
rect 23397 22049 23431 22083
rect 2145 21981 2179 22015
rect 2513 21981 2547 22015
rect 3249 21981 3283 22015
rect 3801 21981 3835 22015
rect 5457 21981 5491 22015
rect 5839 21981 5873 22015
rect 6927 21981 6961 22015
rect 10299 21981 10333 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 15142 21981 15176 22015
rect 16313 21981 16347 22015
rect 16587 21981 16621 22015
rect 18429 21981 18463 22015
rect 19524 21981 19558 22015
rect 20821 21981 20855 22015
rect 21005 21981 21039 22015
rect 22017 21981 22051 22015
rect 22569 21981 22603 22015
rect 23121 21981 23155 22015
rect 23581 21981 23615 22015
rect 24225 21981 24259 22015
rect 1777 21913 1811 21947
rect 2053 21913 2087 21947
rect 4721 21913 4755 21947
rect 4997 21913 5031 21947
rect 5089 21913 5123 21947
rect 11897 21913 11931 21947
rect 11989 21913 12023 21947
rect 12357 21913 12391 21947
rect 23949 21913 23983 21947
rect 2881 21845 2915 21879
rect 3433 21845 3467 21879
rect 7665 21845 7699 21879
rect 11621 21845 11655 21879
rect 12725 21845 12759 21879
rect 15945 21845 15979 21879
rect 18245 21845 18279 21879
rect 20637 21845 20671 21879
rect 21005 21845 21039 21879
rect 22293 21845 22327 21879
rect 23397 21845 23431 21879
rect 24041 21845 24075 21879
rect 2421 21641 2455 21675
rect 2973 21641 3007 21675
rect 3249 21641 3283 21675
rect 5733 21641 5767 21675
rect 8493 21641 8527 21675
rect 9597 21641 9631 21675
rect 9781 21641 9815 21675
rect 12817 21641 12851 21675
rect 14289 21641 14323 21675
rect 20913 21641 20947 21675
rect 22017 21641 22051 21675
rect 24409 21641 24443 21675
rect 6561 21573 6595 21607
rect 6837 21573 6871 21607
rect 6929 21573 6963 21607
rect 7665 21573 7699 21607
rect 24133 21573 24167 21607
rect 1409 21505 1443 21539
rect 1683 21505 1717 21539
rect 2789 21505 2823 21539
rect 3065 21505 3099 21539
rect 4721 21505 4755 21539
rect 4995 21505 5029 21539
rect 7297 21505 7331 21539
rect 8769 21505 8803 21539
rect 8861 21505 8895 21539
rect 9229 21505 9263 21539
rect 12047 21505 12081 21539
rect 13277 21505 13311 21539
rect 13551 21505 13585 21539
rect 15117 21505 15151 21539
rect 15391 21505 15425 21539
rect 17739 21505 17773 21539
rect 18521 21505 18555 21539
rect 18797 21505 18831 21539
rect 18889 21505 18923 21539
rect 19809 21505 19843 21539
rect 19901 21505 19935 21539
rect 20143 21505 20177 21539
rect 21281 21505 21315 21539
rect 21833 21505 21867 21539
rect 23397 21505 23431 21539
rect 23581 21505 23615 21539
rect 23673 21505 23707 21539
rect 11805 21437 11839 21471
rect 16727 21437 16761 21471
rect 16865 21437 16899 21471
rect 17325 21437 17359 21471
rect 17601 21437 17635 21471
rect 17877 21437 17911 21471
rect 21557 21437 21591 21471
rect 18613 21369 18647 21403
rect 21465 21369 21499 21403
rect 7849 21301 7883 21335
rect 15025 21301 15059 21335
rect 16129 21301 16163 21335
rect 18981 21301 19015 21335
rect 19625 21301 19659 21335
rect 21373 21301 21407 21335
rect 23489 21301 23523 21335
rect 23857 21301 23891 21335
rect 2513 21097 2547 21131
rect 8493 21097 8527 21131
rect 9965 21097 9999 21131
rect 17969 21097 18003 21131
rect 20453 21097 20487 21131
rect 2789 21029 2823 21063
rect 18981 21029 19015 21063
rect 20729 21029 20763 21063
rect 7481 20961 7515 20995
rect 8953 20961 8987 20995
rect 10333 20961 10367 20995
rect 11989 20961 12023 20995
rect 14749 20961 14783 20995
rect 15393 20961 15427 20995
rect 15669 20961 15703 20995
rect 15786 20961 15820 20995
rect 15945 20961 15979 20995
rect 16957 20961 16991 20995
rect 18889 20961 18923 20995
rect 22569 20961 22603 20995
rect 1409 20893 1443 20927
rect 1685 20893 1719 20927
rect 2329 20893 2363 20927
rect 2605 20893 2639 20927
rect 3801 20893 3835 20927
rect 4075 20893 4109 20927
rect 7739 20883 7773 20917
rect 9195 20893 9229 20927
rect 10575 20893 10609 20927
rect 12231 20893 12265 20927
rect 14933 20893 14967 20927
rect 17199 20893 17233 20927
rect 18616 20893 18650 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 20361 20893 20395 20927
rect 20913 20893 20947 20927
rect 24041 20893 24075 20927
rect 19073 20825 19107 20859
rect 19349 20825 19383 20859
rect 22814 20825 22848 20859
rect 4813 20757 4847 20791
rect 11345 20757 11379 20791
rect 13001 20757 13035 20791
rect 16589 20757 16623 20791
rect 23949 20757 23983 20791
rect 24133 20757 24167 20791
rect 15393 20553 15427 20587
rect 18797 20553 18831 20587
rect 22477 20553 22511 20587
rect 23765 20553 23799 20587
rect 9965 20485 9999 20519
rect 10241 20485 10275 20519
rect 10701 20485 10735 20519
rect 11069 20485 11103 20519
rect 14197 20485 14231 20519
rect 1683 20417 1717 20451
rect 3065 20417 3099 20451
rect 3801 20417 3835 20451
rect 3918 20417 3952 20451
rect 4077 20417 4111 20451
rect 4813 20417 4847 20451
rect 5087 20417 5121 20451
rect 10333 20417 10367 20451
rect 12541 20417 12575 20451
rect 13394 20417 13428 20451
rect 13553 20417 13587 20451
rect 14381 20417 14415 20451
rect 14655 20417 14689 20451
rect 17785 20417 17819 20451
rect 18059 20417 18093 20451
rect 22385 20417 22419 20451
rect 22661 20417 22695 20451
rect 22753 20417 22787 20451
rect 22995 20417 23029 20451
rect 24133 20417 24167 20451
rect 24225 20417 24259 20451
rect 1409 20349 1443 20383
rect 2881 20349 2915 20383
rect 12357 20349 12391 20383
rect 13001 20349 13035 20383
rect 13277 20349 13311 20383
rect 24409 20349 24443 20383
rect 3525 20281 3559 20315
rect 11253 20281 11287 20315
rect 22201 20281 22235 20315
rect 2421 20213 2455 20247
rect 4721 20213 4755 20247
rect 5825 20213 5859 20247
rect 24317 20213 24351 20247
rect 1593 20009 1627 20043
rect 3341 20009 3375 20043
rect 11161 20009 11195 20043
rect 13553 20009 13587 20043
rect 22109 20009 22143 20043
rect 23949 20009 23983 20043
rect 2329 19873 2363 19907
rect 10149 19873 10183 19907
rect 12541 19873 12575 19907
rect 16313 19873 16347 19907
rect 16589 19873 16623 19907
rect 16727 19873 16761 19907
rect 19257 19873 19291 19907
rect 22201 19873 22235 19907
rect 1501 19805 1535 19839
rect 2571 19805 2605 19839
rect 3801 19805 3835 19839
rect 4905 19805 4939 19839
rect 5457 19805 5491 19839
rect 5917 19805 5951 19839
rect 6653 19805 6687 19839
rect 6927 19805 6961 19839
rect 8217 19805 8251 19839
rect 10423 19805 10457 19839
rect 12783 19805 12817 19839
rect 15669 19805 15703 19839
rect 15853 19805 15887 19839
rect 16865 19805 16899 19839
rect 19073 19805 19107 19839
rect 20729 19805 20763 19839
rect 20985 19805 21019 19839
rect 22443 19805 22477 19839
rect 23673 19805 23707 19839
rect 5181 19737 5215 19771
rect 5549 19737 5583 19771
rect 19502 19737 19536 19771
rect 3985 19669 4019 19703
rect 6285 19669 6319 19703
rect 6469 19669 6503 19703
rect 7665 19669 7699 19703
rect 17509 19669 17543 19703
rect 18889 19669 18923 19703
rect 20637 19669 20671 19703
rect 23213 19669 23247 19703
rect 1593 19465 1627 19499
rect 3065 19465 3099 19499
rect 3525 19465 3559 19499
rect 5917 19465 5951 19499
rect 7113 19465 7147 19499
rect 8217 19465 8251 19499
rect 17693 19465 17727 19499
rect 20177 19465 20211 19499
rect 20821 19465 20855 19499
rect 21189 19465 21223 19499
rect 22385 19465 22419 19499
rect 7849 19397 7883 19431
rect 24133 19397 24167 19431
rect 1409 19329 1443 19363
rect 1685 19329 1719 19363
rect 1959 19329 1993 19363
rect 3249 19329 3283 19363
rect 3341 19329 3375 19363
rect 4905 19329 4939 19363
rect 5179 19329 5213 19363
rect 7389 19329 7423 19363
rect 7481 19329 7515 19363
rect 8861 19329 8895 19363
rect 9135 19329 9169 19363
rect 11803 19329 11837 19363
rect 13449 19329 13483 19363
rect 13703 19329 13737 19363
rect 16681 19329 16715 19363
rect 16923 19329 16957 19363
rect 19165 19329 19199 19363
rect 19439 19329 19473 19363
rect 20545 19329 20579 19363
rect 20913 19329 20947 19363
rect 21097 19329 21131 19363
rect 21373 19329 21407 19363
rect 21833 19329 21867 19363
rect 22109 19329 22143 19363
rect 22477 19329 22511 19363
rect 22661 19329 22695 19363
rect 23397 19329 23431 19363
rect 23581 19329 23615 19363
rect 11529 19261 11563 19295
rect 16497 19261 16531 19295
rect 20821 19261 20855 19295
rect 21005 19261 21039 19295
rect 22385 19261 22419 19295
rect 22569 19261 22603 19295
rect 24409 19261 24443 19295
rect 23213 19193 23247 19227
rect 2697 19125 2731 19159
rect 8401 19125 8435 19159
rect 9873 19125 9907 19159
rect 12541 19125 12575 19159
rect 14473 19125 14507 19159
rect 20637 19125 20671 19159
rect 21925 19125 21959 19159
rect 22201 19125 22235 19159
rect 23857 19125 23891 19159
rect 8125 18921 8159 18955
rect 17049 18921 17083 18955
rect 19717 18921 19751 18955
rect 3249 18853 3283 18887
rect 19993 18853 20027 18887
rect 22845 18853 22879 18887
rect 23581 18853 23615 18887
rect 1593 18785 1627 18819
rect 7113 18785 7147 18819
rect 16037 18785 16071 18819
rect 1867 18717 1901 18751
rect 3801 18717 3835 18751
rect 4075 18717 4109 18751
rect 7355 18717 7389 18751
rect 9413 18717 9447 18751
rect 9505 18717 9539 18751
rect 9873 18717 9907 18751
rect 10255 18717 10289 18751
rect 11253 18717 11287 18751
rect 11527 18717 11561 18751
rect 14565 18717 14599 18751
rect 15025 18717 15059 18751
rect 16311 18717 16345 18751
rect 17601 18717 17635 18751
rect 17843 18717 17877 18751
rect 19625 18717 19659 18751
rect 20177 18717 20211 18751
rect 22753 18717 22787 18751
rect 22937 18717 22971 18751
rect 23213 18717 23247 18751
rect 23397 18717 23431 18751
rect 23857 18717 23891 18751
rect 3065 18649 3099 18683
rect 9137 18649 9171 18683
rect 14289 18649 14323 18683
rect 14657 18649 14691 18683
rect 2605 18581 2639 18615
rect 4813 18581 4847 18615
rect 10425 18581 10459 18615
rect 12265 18581 12299 18615
rect 15393 18581 15427 18615
rect 15577 18581 15611 18615
rect 18613 18581 18647 18615
rect 23029 18581 23063 18615
rect 24133 18581 24167 18615
rect 5549 18377 5583 18411
rect 9229 18377 9263 18411
rect 11713 18377 11747 18411
rect 15209 18377 15243 18411
rect 3525 18309 3559 18343
rect 12081 18309 12115 18343
rect 12817 18309 12851 18343
rect 22814 18309 22848 18343
rect 24133 18309 24167 18343
rect 1501 18241 1535 18275
rect 2053 18241 2087 18275
rect 2327 18241 2361 18275
rect 3985 18241 4019 18275
rect 4259 18241 4293 18275
rect 5457 18241 5491 18275
rect 8217 18241 8251 18275
rect 8491 18241 8525 18275
rect 9871 18241 9905 18275
rect 11345 18241 11379 18275
rect 11989 18241 12023 18275
rect 12449 18241 12483 18275
rect 14197 18241 14231 18275
rect 14471 18241 14505 18275
rect 17141 18241 17175 18275
rect 18337 18241 18371 18275
rect 22569 18241 22603 18275
rect 9597 18173 9631 18207
rect 17325 18173 17359 18207
rect 18061 18173 18095 18207
rect 18199 18173 18233 18207
rect 13001 18105 13035 18139
rect 17785 18105 17819 18139
rect 1593 18037 1627 18071
rect 3065 18037 3099 18071
rect 3617 18037 3651 18071
rect 4997 18037 5031 18071
rect 10609 18037 10643 18071
rect 18981 18037 19015 18071
rect 23949 18037 23983 18071
rect 24409 18037 24443 18071
rect 18153 17833 18187 17867
rect 23765 17833 23799 17867
rect 2421 17765 2455 17799
rect 4445 17765 4479 17799
rect 10425 17765 10459 17799
rect 18705 17765 18739 17799
rect 1961 17697 1995 17731
rect 3801 17697 3835 17731
rect 4721 17697 4755 17731
rect 4859 17697 4893 17731
rect 9781 17697 9815 17731
rect 10818 17697 10852 17731
rect 12081 17697 12115 17731
rect 12725 17697 12759 17731
rect 13001 17697 13035 17731
rect 14289 17697 14323 17731
rect 17141 17697 17175 17731
rect 20729 17697 20763 17731
rect 22753 17697 22787 17731
rect 1409 17629 1443 17663
rect 1777 17629 1811 17663
rect 2697 17629 2731 17663
rect 2814 17629 2848 17663
rect 2973 17629 3007 17663
rect 3985 17629 4019 17663
rect 4997 17629 5031 17663
rect 5733 17629 5767 17663
rect 5991 17599 6025 17633
rect 9965 17629 9999 17663
rect 10701 17629 10735 17663
rect 10977 17629 11011 17663
rect 11621 17629 11655 17663
rect 11713 17629 11747 17663
rect 12265 17629 12299 17663
rect 13118 17629 13152 17663
rect 13277 17629 13311 17663
rect 17383 17629 17417 17663
rect 19257 17629 19291 17663
rect 22201 17629 22235 17663
rect 22661 17629 22695 17663
rect 23011 17599 23045 17633
rect 19502 17561 19536 17595
rect 20974 17561 21008 17595
rect 1593 17493 1627 17527
rect 3617 17493 3651 17527
rect 5641 17493 5675 17527
rect 6745 17493 6779 17527
rect 11897 17493 11931 17527
rect 13921 17493 13955 17527
rect 20637 17493 20671 17527
rect 22109 17493 22143 17527
rect 22293 17493 22327 17527
rect 22477 17493 22511 17527
rect 7849 17289 7883 17323
rect 8309 17289 8343 17323
rect 11069 17289 11103 17323
rect 13645 17289 13679 17323
rect 19533 17289 19567 17323
rect 20545 17289 20579 17323
rect 21005 17289 21039 17323
rect 23581 17289 23615 17323
rect 3525 17221 3559 17255
rect 6561 17221 6595 17255
rect 7665 17221 7699 17255
rect 1593 17153 1627 17187
rect 2881 17153 2915 17187
rect 3801 17153 3835 17187
rect 4905 17153 4939 17187
rect 5163 17183 5197 17217
rect 6837 17153 6871 17187
rect 6929 17153 6963 17187
rect 7297 17153 7331 17187
rect 10045 17153 10079 17187
rect 10331 17153 10365 17187
rect 12265 17153 12299 17187
rect 12633 17153 12667 17187
rect 12907 17153 12941 17187
rect 15451 17153 15485 17187
rect 16955 17153 16989 17187
rect 19717 17153 19751 17187
rect 20085 17153 20119 17187
rect 20729 17153 20763 17187
rect 21189 17153 21223 17187
rect 21465 17153 21499 17187
rect 21649 17153 21683 17187
rect 22075 17153 22109 17187
rect 23397 17153 23431 17187
rect 23857 17153 23891 17187
rect 24317 17153 24351 17187
rect 1685 17085 1719 17119
rect 1869 17085 1903 17119
rect 2329 17085 2363 17119
rect 2605 17085 2639 17119
rect 2743 17085 2777 17119
rect 15209 17085 15243 17119
rect 16681 17085 16715 17119
rect 21833 17085 21867 17119
rect 3617 17017 3651 17051
rect 5917 17017 5951 17051
rect 1409 16949 1443 16983
rect 12449 16949 12483 16983
rect 14473 16949 14507 16983
rect 16221 16949 16255 16983
rect 17693 16949 17727 16983
rect 20177 16949 20211 16983
rect 21557 16949 21591 16983
rect 22845 16949 22879 16983
rect 24133 16949 24167 16983
rect 24409 16949 24443 16983
rect 8769 16745 8803 16779
rect 15577 16745 15611 16779
rect 21281 16745 21315 16779
rect 22017 16745 22051 16779
rect 7573 16677 7607 16711
rect 13645 16677 13679 16711
rect 16405 16677 16439 16711
rect 22109 16677 22143 16711
rect 1777 16609 1811 16643
rect 2053 16609 2087 16643
rect 6929 16609 6963 16643
rect 7113 16609 7147 16643
rect 8125 16609 8159 16643
rect 12633 16609 12667 16643
rect 16798 16609 16832 16643
rect 16957 16609 16991 16643
rect 19809 16609 19843 16643
rect 21465 16609 21499 16643
rect 22201 16609 22235 16643
rect 1409 16541 1443 16575
rect 3617 16541 3651 16575
rect 7849 16541 7883 16575
rect 7987 16541 8021 16575
rect 12907 16541 12941 16575
rect 14565 16541 14599 16575
rect 15761 16541 15795 16575
rect 15945 16541 15979 16575
rect 16681 16541 16715 16575
rect 17601 16541 17635 16575
rect 17693 16541 17727 16575
rect 20067 16511 20101 16545
rect 21189 16541 21223 16575
rect 21925 16541 21959 16575
rect 23489 16541 23523 16575
rect 23673 16541 23707 16575
rect 2973 16473 3007 16507
rect 3893 16473 3927 16507
rect 14289 16473 14323 16507
rect 14657 16473 14691 16507
rect 15025 16473 15059 16507
rect 21465 16473 21499 16507
rect 24041 16473 24075 16507
rect 1593 16405 1627 16439
rect 3065 16405 3099 16439
rect 3433 16405 3467 16439
rect 3985 16405 4019 16439
rect 15393 16405 15427 16439
rect 17877 16405 17911 16439
rect 20821 16405 20855 16439
rect 23305 16405 23339 16439
rect 8493 16201 8527 16235
rect 13093 16201 13127 16235
rect 15393 16201 15427 16235
rect 19257 16201 19291 16235
rect 20821 16201 20855 16235
rect 24317 16201 24351 16235
rect 1685 16133 1719 16167
rect 2053 16133 2087 16167
rect 5365 16133 5399 16167
rect 18144 16133 18178 16167
rect 2145 16065 2179 16099
rect 2403 16095 2437 16129
rect 3525 16065 3559 16099
rect 4445 16065 4479 16099
rect 7723 16065 7757 16099
rect 8861 16065 8895 16099
rect 9135 16065 9169 16099
rect 10609 16065 10643 16099
rect 12081 16065 12115 16099
rect 12355 16065 12389 16099
rect 14655 16065 14689 16099
rect 19349 16065 19383 16099
rect 19809 16065 19843 16099
rect 20637 16065 20671 16099
rect 20821 16065 20855 16099
rect 22903 16065 22937 16099
rect 24041 16065 24075 16099
rect 24133 16065 24167 16099
rect 3709 15997 3743 16031
rect 4583 15997 4617 16031
rect 4721 15997 4755 16031
rect 7481 15997 7515 16031
rect 14381 15997 14415 16031
rect 17877 15997 17911 16031
rect 22661 15997 22695 16031
rect 24317 15997 24351 16031
rect 3157 15929 3191 15963
rect 4169 15929 4203 15963
rect 9873 15861 9907 15895
rect 10425 15861 10459 15895
rect 19441 15861 19475 15895
rect 19625 15861 19659 15895
rect 23673 15861 23707 15895
rect 1777 15657 1811 15691
rect 2881 15657 2915 15691
rect 4813 15657 4847 15691
rect 7849 15657 7883 15691
rect 10793 15657 10827 15691
rect 18337 15657 18371 15691
rect 24133 15657 24167 15691
rect 9597 15589 9631 15623
rect 5457 15521 5491 15555
rect 6837 15521 6871 15555
rect 9990 15521 10024 15555
rect 19257 15521 19291 15555
rect 22385 15521 22419 15555
rect 1685 15453 1719 15487
rect 2237 15453 2271 15487
rect 2789 15453 2823 15487
rect 3433 15453 3467 15487
rect 3801 15453 3835 15487
rect 4075 15453 4109 15487
rect 5699 15453 5733 15487
rect 7079 15453 7113 15487
rect 8953 15453 8987 15487
rect 9137 15453 9171 15487
rect 9873 15453 9907 15487
rect 10149 15453 10183 15487
rect 10885 15453 10919 15487
rect 11159 15453 11193 15487
rect 18521 15453 18555 15487
rect 19515 15423 19549 15457
rect 22293 15453 22327 15487
rect 23949 15453 23983 15487
rect 22630 15385 22664 15419
rect 2329 15317 2363 15351
rect 3249 15317 3283 15351
rect 6469 15317 6503 15351
rect 11897 15317 11931 15351
rect 20269 15317 20303 15351
rect 22109 15317 22143 15351
rect 23765 15317 23799 15351
rect 1593 15113 1627 15147
rect 3433 15113 3467 15147
rect 3985 15113 4019 15147
rect 10241 15113 10275 15147
rect 11713 15113 11747 15147
rect 12817 15113 12851 15147
rect 19717 15113 19751 15147
rect 3341 15045 3375 15079
rect 20536 15045 20570 15079
rect 23765 15045 23799 15079
rect 1777 14977 1811 15011
rect 1869 14977 1903 15011
rect 2143 14987 2177 15021
rect 3893 14977 3927 15011
rect 4627 14977 4661 15011
rect 6561 14977 6595 15011
rect 7435 14977 7469 15011
rect 9229 14977 9263 15011
rect 9487 14977 9521 15011
rect 11989 14977 12023 15011
rect 12081 14977 12115 15011
rect 12449 14977 12483 15011
rect 14163 14987 14197 15021
rect 17141 14977 17175 15011
rect 17408 14977 17442 15011
rect 19441 14977 19475 15011
rect 19533 14977 19567 15011
rect 19809 14977 19843 15011
rect 19993 14977 20027 15011
rect 20269 14977 20303 15011
rect 22075 14977 22109 15011
rect 23397 14977 23431 15011
rect 24225 14977 24259 15011
rect 4353 14909 4387 14943
rect 6377 14909 6411 14943
rect 7297 14909 7331 14943
rect 7573 14909 7607 14943
rect 13921 14909 13955 14943
rect 19717 14909 19751 14943
rect 19901 14909 19935 14943
rect 21833 14909 21867 14943
rect 24501 14909 24535 14943
rect 7021 14841 7055 14875
rect 22845 14841 22879 14875
rect 23489 14841 23523 14875
rect 24317 14841 24351 14875
rect 2881 14773 2915 14807
rect 5365 14773 5399 14807
rect 8217 14773 8251 14807
rect 13001 14773 13035 14807
rect 14933 14773 14967 14807
rect 18521 14773 18555 14807
rect 21649 14773 21683 14807
rect 24041 14773 24075 14807
rect 24409 14773 24443 14807
rect 4077 14569 4111 14603
rect 7849 14569 7883 14603
rect 12265 14569 12299 14603
rect 18061 14569 18095 14603
rect 2421 14501 2455 14535
rect 5549 14501 5583 14535
rect 21557 14501 21591 14535
rect 21925 14501 21959 14535
rect 23581 14501 23615 14535
rect 2835 14433 2869 14467
rect 4629 14433 4663 14467
rect 5963 14433 5997 14467
rect 6837 14433 6871 14467
rect 11253 14433 11287 14467
rect 14473 14433 14507 14467
rect 14933 14433 14967 14467
rect 15209 14433 15243 14467
rect 15347 14433 15381 14467
rect 16865 14433 16899 14467
rect 17141 14433 17175 14467
rect 17258 14433 17292 14467
rect 22109 14433 22143 14467
rect 22569 14433 22603 14467
rect 1777 14365 1811 14399
rect 1961 14365 1995 14399
rect 2697 14365 2731 14399
rect 2973 14365 3007 14399
rect 3985 14365 4019 14399
rect 4261 14365 4295 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 5825 14365 5859 14399
rect 6101 14365 6135 14399
rect 7095 14335 7129 14369
rect 11495 14365 11529 14399
rect 12633 14365 12667 14399
rect 12907 14365 12941 14399
rect 14289 14365 14323 14399
rect 15485 14365 15519 14399
rect 16221 14365 16255 14399
rect 16405 14365 16439 14399
rect 17417 14365 17451 14399
rect 18337 14365 18371 14399
rect 18429 14365 18463 14399
rect 18889 14365 18923 14399
rect 21097 14365 21131 14399
rect 21465 14365 21499 14399
rect 21833 14365 21867 14399
rect 22377 14365 22411 14399
rect 22477 14365 22511 14399
rect 22661 14365 22695 14399
rect 23305 14365 23339 14399
rect 23397 14365 23431 14399
rect 23857 14365 23891 14399
rect 16129 14297 16163 14331
rect 3617 14229 3651 14263
rect 3801 14229 3835 14263
rect 6745 14229 6779 14263
rect 13645 14229 13679 14263
rect 18153 14229 18187 14263
rect 18521 14229 18555 14263
rect 18705 14229 18739 14263
rect 20913 14229 20947 14263
rect 22109 14229 22143 14263
rect 22201 14229 22235 14263
rect 23121 14229 23155 14263
rect 24133 14229 24167 14263
rect 3249 14025 3283 14059
rect 3801 14025 3835 14059
rect 5917 14025 5951 14059
rect 10609 14025 10643 14059
rect 14289 14025 14323 14059
rect 15669 14025 15703 14059
rect 17693 14025 17727 14059
rect 23213 14025 23247 14059
rect 1501 13957 1535 13991
rect 23857 13957 23891 13991
rect 24133 13957 24167 13991
rect 2145 13889 2179 13923
rect 2511 13889 2545 13923
rect 3709 13889 3743 13923
rect 4353 13889 4387 13923
rect 4629 13889 4663 13923
rect 4905 13889 4939 13923
rect 5179 13889 5213 13923
rect 7111 13889 7145 13923
rect 8217 13889 8251 13923
rect 8491 13889 8525 13923
rect 9597 13889 9631 13923
rect 9855 13919 9889 13953
rect 12449 13889 12483 13923
rect 13645 13889 13679 13923
rect 14899 13889 14933 13923
rect 16955 13889 16989 13923
rect 18303 13889 18337 13923
rect 19441 13889 19475 13923
rect 19625 13889 19659 13923
rect 22753 13889 22787 13923
rect 22928 13895 22962 13929
rect 23029 13889 23063 13923
rect 23213 13889 23247 13923
rect 23489 13889 23523 13923
rect 1777 13821 1811 13855
rect 2237 13821 2271 13855
rect 6837 13821 6871 13855
rect 12633 13821 12667 13855
rect 13093 13821 13127 13855
rect 13369 13821 13403 13855
rect 13507 13821 13541 13855
rect 14657 13821 14691 13855
rect 16681 13821 16715 13855
rect 18061 13821 18095 13855
rect 22845 13821 22879 13855
rect 23581 13821 23615 13855
rect 23489 13753 23523 13787
rect 1961 13685 1995 13719
rect 4169 13685 4203 13719
rect 4445 13685 4479 13719
rect 7849 13685 7883 13719
rect 9229 13685 9263 13719
rect 19073 13685 19107 13719
rect 19533 13685 19567 13719
rect 24409 13685 24443 13719
rect 2697 13481 2731 13515
rect 3249 13481 3283 13515
rect 11621 13481 11655 13515
rect 13645 13481 13679 13515
rect 16497 13481 16531 13515
rect 18613 13481 18647 13515
rect 22293 13481 22327 13515
rect 22661 13481 22695 13515
rect 9321 13413 9355 13447
rect 10425 13413 10459 13447
rect 18705 13413 18739 13447
rect 1777 13345 1811 13379
rect 9965 13345 9999 13379
rect 10839 13345 10873 13379
rect 15485 13345 15519 13379
rect 18797 13345 18831 13379
rect 20453 13345 20487 13379
rect 22845 13345 22879 13379
rect 1501 13277 1535 13311
rect 2053 13277 2087 13311
rect 3801 13277 3835 13311
rect 4075 13277 4109 13311
rect 9505 13277 9539 13311
rect 9781 13277 9815 13311
rect 10701 13277 10735 13311
rect 10977 13277 11011 13311
rect 12633 13277 12667 13311
rect 12907 13277 12941 13311
rect 15727 13277 15761 13311
rect 18521 13277 18555 13311
rect 19717 13277 19751 13311
rect 19901 13277 19935 13311
rect 20361 13277 20395 13311
rect 20637 13277 20671 13311
rect 20821 13277 20855 13311
rect 22477 13277 22511 13311
rect 22569 13277 22603 13311
rect 2421 13209 2455 13243
rect 2605 13209 2639 13243
rect 3157 13209 3191 13243
rect 20177 13209 20211 13243
rect 20269 13209 20303 13243
rect 20729 13209 20763 13243
rect 23112 13209 23146 13243
rect 4813 13141 4847 13175
rect 24225 13141 24259 13175
rect 1777 12937 1811 12971
rect 9873 12937 9907 12971
rect 11069 12937 11103 12971
rect 21005 12937 21039 12971
rect 22201 12937 22235 12971
rect 23397 12937 23431 12971
rect 23949 12869 23983 12903
rect 1685 12801 1719 12835
rect 2603 12811 2637 12845
rect 3709 12801 3743 12835
rect 4905 12801 4939 12835
rect 6377 12801 6411 12835
rect 6619 12801 6653 12835
rect 8217 12801 8251 12835
rect 8953 12801 8987 12835
rect 9229 12801 9263 12835
rect 10057 12801 10091 12835
rect 10331 12801 10365 12835
rect 11987 12801 12021 12835
rect 13921 12801 13955 12835
rect 14195 12801 14229 12835
rect 17015 12801 17049 12835
rect 18487 12801 18521 12835
rect 19625 12801 19659 12835
rect 19892 12801 19926 12835
rect 21281 12801 21315 12835
rect 21557 12801 21591 12835
rect 22109 12801 22143 12835
rect 22385 12801 22419 12835
rect 22643 12831 22677 12865
rect 2329 12733 2363 12767
rect 3893 12733 3927 12767
rect 4353 12733 4387 12767
rect 4647 12733 4681 12767
rect 4746 12733 4780 12767
rect 8033 12733 8067 12767
rect 9070 12733 9104 12767
rect 11713 12733 11747 12767
rect 16773 12733 16807 12767
rect 18245 12733 18279 12767
rect 8677 12665 8711 12699
rect 19257 12665 19291 12699
rect 21373 12665 21407 12699
rect 3341 12597 3375 12631
rect 5549 12597 5583 12631
rect 7389 12597 7423 12631
rect 12725 12597 12759 12631
rect 14933 12597 14967 12631
rect 17785 12597 17819 12631
rect 21097 12597 21131 12631
rect 24225 12597 24259 12631
rect 4169 12393 4203 12427
rect 8677 12393 8711 12427
rect 15577 12393 15611 12427
rect 22661 12393 22695 12427
rect 24133 12393 24167 12427
rect 23305 12325 23339 12359
rect 23765 12325 23799 12359
rect 1777 12257 1811 12291
rect 1961 12257 1995 12291
rect 2421 12257 2455 12291
rect 2973 12257 3007 12291
rect 3617 12257 3651 12291
rect 4905 12257 4939 12291
rect 5549 12257 5583 12291
rect 5825 12257 5859 12291
rect 5963 12257 5997 12291
rect 6837 12257 6871 12291
rect 7481 12257 7515 12291
rect 7757 12257 7791 12291
rect 7895 12257 7929 12291
rect 17049 12257 17083 12291
rect 17442 12257 17476 12291
rect 17601 12257 17635 12291
rect 19901 12257 19935 12291
rect 21281 12257 21315 12291
rect 2697 12189 2731 12223
rect 2835 12189 2869 12223
rect 3893 12189 3927 12223
rect 5089 12189 5123 12223
rect 6101 12189 6135 12223
rect 7021 12189 7055 12223
rect 8033 12189 8067 12223
rect 11897 12189 11931 12223
rect 14657 12189 14691 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 17325 12189 17359 12223
rect 20143 12189 20177 12223
rect 22753 12189 22787 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 23489 12189 23523 12223
rect 23581 12189 23615 12223
rect 23949 12189 23983 12223
rect 4445 12121 4479 12155
rect 11805 12121 11839 12155
rect 12265 12121 12299 12155
rect 14565 12121 14599 12155
rect 15025 12121 15059 12155
rect 21548 12121 21582 12155
rect 4537 12053 4571 12087
rect 6745 12053 6779 12087
rect 11529 12053 11563 12087
rect 12633 12053 12667 12087
rect 12817 12053 12851 12087
rect 14289 12053 14323 12087
rect 15393 12053 15427 12087
rect 18245 12053 18279 12087
rect 20913 12053 20947 12087
rect 22845 12053 22879 12087
rect 23121 12053 23155 12087
rect 2881 11849 2915 11883
rect 4537 11849 4571 11883
rect 5917 11849 5951 11883
rect 7941 11849 7975 11883
rect 12541 11849 12575 11883
rect 13921 11849 13955 11883
rect 15945 11849 15979 11883
rect 17693 11849 17727 11883
rect 21465 11849 21499 11883
rect 2143 11713 2177 11747
rect 3433 11713 3467 11747
rect 3525 11713 3559 11747
rect 3799 11723 3833 11757
rect 5163 11743 5197 11777
rect 7203 11713 7237 11747
rect 8583 11713 8617 11747
rect 11529 11713 11563 11747
rect 11803 11713 11837 11747
rect 13183 11713 13217 11747
rect 14933 11713 14967 11747
rect 15207 11713 15241 11747
rect 16923 11713 16957 11747
rect 18061 11713 18095 11747
rect 18319 11743 18353 11777
rect 21649 11713 21683 11747
rect 21925 11713 21959 11747
rect 22385 11713 22419 11747
rect 22753 11713 22787 11747
rect 23305 11713 23339 11747
rect 23581 11713 23615 11747
rect 23673 11713 23707 11747
rect 24133 11713 24167 11747
rect 1869 11645 1903 11679
rect 4905 11645 4939 11679
rect 6929 11645 6963 11679
rect 8309 11645 8343 11679
rect 12909 11645 12943 11679
rect 16681 11645 16715 11679
rect 22661 11577 22695 11611
rect 23121 11577 23155 11611
rect 3249 11509 3283 11543
rect 9321 11509 9355 11543
rect 19073 11509 19107 11543
rect 23397 11509 23431 11543
rect 23857 11509 23891 11543
rect 24409 11509 24443 11543
rect 2145 11305 2179 11339
rect 3433 11305 3467 11339
rect 4537 11305 4571 11339
rect 5089 11305 5123 11339
rect 7665 11305 7699 11339
rect 11069 11305 11103 11339
rect 11529 11305 11563 11339
rect 18153 11305 18187 11339
rect 23765 11305 23799 11339
rect 1685 11237 1719 11271
rect 2605 11237 2639 11271
rect 5457 11237 5491 11271
rect 9597 11237 9631 11271
rect 15853 11237 15887 11271
rect 17049 11237 17083 11271
rect 18705 11237 18739 11271
rect 20729 11237 20763 11271
rect 8953 11169 8987 11203
rect 15393 11169 15427 11203
rect 16246 11169 16280 11203
rect 16405 11169 16439 11203
rect 18889 11169 18923 11203
rect 22753 11169 22787 11203
rect 1501 11101 1535 11135
rect 2789 11101 2823 11135
rect 3617 11101 3651 11135
rect 3893 11101 3927 11135
rect 4997 11101 5031 11135
rect 5641 11101 5675 11135
rect 6653 11101 6687 11135
rect 6927 11101 6961 11135
rect 8493 11101 8527 11135
rect 9137 11101 9171 11135
rect 9873 11101 9907 11135
rect 9990 11101 10024 11135
rect 10149 11101 10183 11135
rect 15209 11101 15243 11135
rect 16129 11101 16163 11135
rect 17141 11101 17175 11135
rect 17415 11101 17449 11135
rect 18705 11101 18739 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 20085 11101 20119 11135
rect 20269 11101 20303 11135
rect 20729 11101 20763 11135
rect 22995 11101 23029 11135
rect 2053 11033 2087 11067
rect 2973 11033 3007 11067
rect 4445 11033 4479 11067
rect 10793 11033 10827 11067
rect 19073 11033 19107 11067
rect 19349 11033 19383 11067
rect 3065 10965 3099 10999
rect 3985 10965 4019 10999
rect 1593 10761 1627 10795
rect 3801 10761 3835 10795
rect 10241 10761 10275 10795
rect 10977 10761 11011 10795
rect 14933 10761 14967 10795
rect 20269 10761 20303 10795
rect 20729 10761 20763 10795
rect 1501 10693 1535 10727
rect 13645 10693 13679 10727
rect 13921 10693 13955 10727
rect 14381 10693 14415 10727
rect 14749 10693 14783 10727
rect 2145 10625 2179 10659
rect 2495 10655 2529 10689
rect 3985 10625 4019 10659
rect 4351 10625 4385 10659
rect 6619 10625 6653 10659
rect 9471 10625 9505 10659
rect 10793 10625 10827 10659
rect 12355 10625 12389 10659
rect 14013 10625 14047 10659
rect 17693 10625 17727 10659
rect 17785 10625 17819 10659
rect 18041 10625 18075 10659
rect 19531 10625 19565 10659
rect 20637 10625 20671 10659
rect 20821 10625 20855 10659
rect 21097 10625 21131 10659
rect 22661 10625 22695 10659
rect 22753 10625 22787 10659
rect 22995 10625 23029 10659
rect 2237 10557 2271 10591
rect 4077 10557 4111 10591
rect 6377 10557 6411 10591
rect 9229 10557 9263 10591
rect 12081 10557 12115 10591
rect 19257 10557 19291 10591
rect 13093 10489 13127 10523
rect 20913 10489 20947 10523
rect 1961 10421 1995 10455
rect 3249 10421 3283 10455
rect 5089 10421 5123 10455
rect 7389 10421 7423 10455
rect 17509 10421 17543 10455
rect 19165 10421 19199 10455
rect 22477 10421 22511 10455
rect 23765 10421 23799 10455
rect 3617 10217 3651 10251
rect 7573 10217 7607 10251
rect 15117 10217 15151 10251
rect 18429 10217 18463 10251
rect 20177 10217 20211 10251
rect 10977 10149 11011 10183
rect 20361 10149 20395 10183
rect 1961 10081 1995 10115
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 3985 10081 4019 10115
rect 4445 10081 4479 10115
rect 4721 10081 4755 10115
rect 4838 10081 4872 10115
rect 4997 10081 5031 10115
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 6770 10081 6804 10115
rect 6929 10081 6963 10115
rect 20821 10081 20855 10115
rect 1777 10013 1811 10047
rect 2835 10013 2869 10047
rect 2973 10013 3007 10047
rect 3801 10013 3835 10047
rect 5733 10013 5767 10047
rect 5917 10013 5951 10047
rect 9965 10013 9999 10047
rect 10239 10013 10273 10047
rect 11897 10013 11931 10047
rect 14105 10013 14139 10047
rect 14363 9983 14397 10017
rect 18337 10013 18371 10047
rect 19073 10013 19107 10047
rect 20085 10013 20119 10047
rect 20545 10013 20579 10047
rect 21063 10013 21097 10047
rect 22477 10013 22511 10047
rect 22753 10013 22787 10047
rect 22995 10013 23029 10047
rect 11805 9945 11839 9979
rect 12265 9945 12299 9979
rect 5641 9877 5675 9911
rect 11529 9877 11563 9911
rect 12633 9877 12667 9911
rect 12817 9877 12851 9911
rect 18889 9877 18923 9911
rect 21833 9877 21867 9911
rect 22293 9877 22327 9911
rect 23765 9877 23799 9911
rect 2697 9673 2731 9707
rect 4537 9673 4571 9707
rect 5917 9673 5951 9707
rect 11253 9673 11287 9707
rect 12817 9673 12851 9707
rect 21097 9673 21131 9707
rect 1593 9537 1627 9571
rect 1927 9537 1961 9571
rect 3249 9537 3283 9571
rect 3767 9537 3801 9571
rect 5147 9537 5181 9571
rect 7665 9537 7699 9571
rect 8401 9537 8435 9571
rect 8663 9537 8697 9571
rect 9321 9537 9355 9571
rect 9413 9537 9447 9571
rect 10333 9537 10367 9571
rect 10471 9537 10505 9571
rect 10609 9537 10643 9571
rect 11805 9537 11839 9571
rect 12079 9537 12113 9571
rect 18337 9537 18371 9571
rect 18595 9567 18629 9601
rect 19984 9537 20018 9571
rect 21833 9537 21867 9571
rect 22109 9537 22143 9571
rect 22293 9537 22327 9571
rect 22569 9537 22603 9571
rect 22995 9537 23029 9571
rect 24317 9537 24351 9571
rect 1685 9469 1719 9503
rect 3513 9469 3547 9503
rect 4905 9469 4939 9503
rect 7481 9469 7515 9503
rect 8539 9469 8573 9503
rect 9597 9469 9631 9503
rect 19717 9469 19751 9503
rect 22753 9469 22787 9503
rect 8125 9401 8159 9435
rect 10057 9401 10091 9435
rect 22385 9401 22419 9435
rect 23765 9401 23799 9435
rect 1409 9333 1443 9367
rect 3065 9333 3099 9367
rect 19349 9333 19383 9367
rect 21925 9333 21959 9367
rect 22201 9333 22235 9367
rect 24133 9333 24167 9367
rect 2697 9129 2731 9163
rect 4077 9129 4111 9163
rect 8493 9129 8527 9163
rect 10793 9129 10827 9163
rect 22661 9129 22695 9163
rect 23397 9129 23431 9163
rect 23949 9129 23983 9163
rect 1685 9061 1719 9095
rect 2237 9061 2271 9095
rect 9781 8993 9815 9027
rect 14105 8993 14139 9027
rect 21281 8993 21315 9027
rect 2053 8925 2087 8959
rect 3157 8925 3191 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 7481 8925 7515 8959
rect 7755 8925 7789 8959
rect 10055 8925 10089 8959
rect 14347 8925 14381 8959
rect 15485 8925 15519 8959
rect 15759 8925 15793 8959
rect 16865 8925 16899 8959
rect 17107 8925 17141 8959
rect 22937 8925 22971 8959
rect 23673 8925 23707 8959
rect 1501 8857 1535 8891
rect 2605 8857 2639 8891
rect 21548 8857 21582 8891
rect 23121 8857 23155 8891
rect 3249 8789 3283 8823
rect 3801 8789 3835 8823
rect 15117 8789 15151 8823
rect 16497 8789 16531 8823
rect 17877 8789 17911 8823
rect 22753 8789 22787 8823
rect 2697 8585 2731 8619
rect 7113 8585 7147 8619
rect 8401 8585 8435 8619
rect 10149 8585 10183 8619
rect 13001 8585 13035 8619
rect 17141 8585 17175 8619
rect 19625 8585 19659 8619
rect 1501 8517 1535 8551
rect 2421 8517 2455 8551
rect 2605 8517 2639 8551
rect 11713 8517 11747 8551
rect 12817 8517 12851 8551
rect 13829 8517 13863 8551
rect 14197 8517 14231 8551
rect 14933 8517 14967 8551
rect 17417 8517 17451 8551
rect 17509 8517 17543 8551
rect 18245 8517 18279 8551
rect 1869 8449 1903 8483
rect 2053 8449 2087 8483
rect 3157 8449 3191 8483
rect 3709 8449 3743 8483
rect 7297 8449 7331 8483
rect 7663 8449 7697 8483
rect 9379 8449 9413 8483
rect 11989 8449 12023 8483
rect 12081 8449 12115 8483
rect 12449 8449 12483 8483
rect 14105 8449 14139 8483
rect 14565 8449 14599 8483
rect 17877 8449 17911 8483
rect 18855 8449 18889 8483
rect 19993 8449 20027 8483
rect 20177 8449 20211 8483
rect 22201 8449 22235 8483
rect 22661 8449 22695 8483
rect 23489 8449 23523 8483
rect 24041 8449 24075 8483
rect 24501 8449 24535 8483
rect 7389 8381 7423 8415
rect 9137 8381 9171 8415
rect 18613 8381 18647 8415
rect 22017 8381 22051 8415
rect 23305 8381 23339 8415
rect 23949 8381 23983 8415
rect 3341 8313 3375 8347
rect 3893 8313 3927 8347
rect 15117 8313 15151 8347
rect 22661 8313 22695 8347
rect 18429 8245 18463 8279
rect 20085 8245 20119 8279
rect 24317 8245 24351 8279
rect 1593 8041 1627 8075
rect 3341 8041 3375 8075
rect 8125 8041 8159 8075
rect 10885 8041 10919 8075
rect 12265 8041 12299 8075
rect 13645 8041 13679 8075
rect 18245 8041 18279 8075
rect 19901 8041 19935 8075
rect 22661 8041 22695 8075
rect 3801 7973 3835 8007
rect 5917 7973 5951 8007
rect 6929 7973 6963 8007
rect 15945 7973 15979 8007
rect 19441 7973 19475 8007
rect 21097 7973 21131 8007
rect 6285 7905 6319 7939
rect 7205 7905 7239 7939
rect 12633 7905 12667 7939
rect 16338 7905 16372 7939
rect 16497 7905 16531 7939
rect 18889 7905 18923 7939
rect 1961 7837 1995 7871
rect 2235 7837 2269 7871
rect 3525 7837 3559 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4905 7837 4939 7871
rect 5179 7837 5213 7871
rect 6469 7837 6503 7871
rect 7343 7837 7377 7871
rect 7481 7837 7515 7871
rect 9873 7837 9907 7871
rect 10147 7837 10181 7871
rect 11253 7837 11287 7871
rect 11527 7837 11561 7871
rect 12875 7837 12909 7871
rect 15301 7837 15335 7871
rect 15485 7837 15519 7871
rect 16221 7837 16255 7871
rect 17233 7837 17267 7871
rect 17491 7807 17525 7841
rect 18797 7837 18831 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 20085 7837 20119 7871
rect 20361 7837 20395 7871
rect 20637 7837 20671 7871
rect 21097 7837 21131 7871
rect 22477 7837 22511 7871
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 1501 7769 1535 7803
rect 19809 7769 19843 7803
rect 23112 7769 23146 7803
rect 2973 7701 3007 7735
rect 4077 7701 4111 7735
rect 17141 7701 17175 7735
rect 22293 7701 22327 7735
rect 24225 7701 24259 7735
rect 1777 7497 1811 7531
rect 2145 7497 2179 7531
rect 4261 7497 4295 7531
rect 7481 7497 7515 7531
rect 19533 7497 19567 7531
rect 19993 7497 20027 7531
rect 21557 7497 21591 7531
rect 23305 7497 23339 7531
rect 24133 7497 24167 7531
rect 1685 7429 1719 7463
rect 13277 7429 13311 7463
rect 13553 7429 13587 7463
rect 14381 7429 14415 7463
rect 23857 7429 23891 7463
rect 2329 7361 2363 7395
rect 2605 7361 2639 7395
rect 3341 7361 3375 7395
rect 3617 7361 3651 7395
rect 5411 7361 5445 7395
rect 5549 7361 5583 7395
rect 6743 7361 6777 7395
rect 8291 7391 8325 7425
rect 9413 7361 9447 7395
rect 9687 7361 9721 7395
rect 13645 7361 13679 7395
rect 14013 7361 14047 7395
rect 18153 7361 18187 7395
rect 18420 7361 18454 7395
rect 19901 7361 19935 7395
rect 20444 7361 20478 7395
rect 22017 7361 22051 7395
rect 22567 7361 22601 7395
rect 24501 7361 24535 7395
rect 2421 7293 2455 7327
rect 3065 7293 3099 7327
rect 3479 7293 3513 7327
rect 4353 7293 4387 7327
rect 4537 7293 4571 7327
rect 5273 7293 5307 7327
rect 6469 7293 6503 7327
rect 8033 7293 8067 7327
rect 20177 7293 20211 7327
rect 22293 7293 22327 7327
rect 4997 7225 5031 7259
rect 14565 7225 14599 7259
rect 24317 7225 24351 7259
rect 6193 7157 6227 7191
rect 9045 7157 9079 7191
rect 10425 7157 10459 7191
rect 21833 7157 21867 7191
rect 1593 6953 1627 6987
rect 3341 6953 3375 6987
rect 5549 6953 5583 6987
rect 13553 6953 13587 6987
rect 18613 6953 18647 6987
rect 20729 6953 20763 6987
rect 21097 6953 21131 6987
rect 9597 6885 9631 6919
rect 20361 6885 20395 6919
rect 21741 6885 21775 6919
rect 22661 6885 22695 6919
rect 2329 6817 2363 6851
rect 4537 6817 4571 6851
rect 8953 6817 8987 6851
rect 10149 6817 10183 6851
rect 21373 6817 21407 6851
rect 24041 6817 24075 6851
rect 2237 6749 2271 6783
rect 2603 6749 2637 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 4811 6749 4845 6783
rect 9137 6749 9171 6783
rect 9873 6749 9907 6783
rect 9990 6749 10024 6783
rect 12541 6749 12575 6783
rect 12799 6719 12833 6753
rect 18797 6749 18831 6783
rect 19349 6749 19383 6783
rect 19623 6749 19657 6783
rect 20913 6749 20947 6783
rect 21005 6749 21039 6783
rect 21189 6749 21223 6783
rect 21281 6749 21315 6783
rect 21557 6749 21591 6783
rect 22017 6749 22051 6783
rect 22385 6749 22419 6783
rect 22753 6749 22787 6783
rect 23397 6749 23431 6783
rect 23489 6749 23523 6783
rect 23949 6749 23983 6783
rect 24133 6749 24167 6783
rect 1501 6681 1535 6715
rect 2053 6613 2087 6647
rect 3801 6613 3835 6647
rect 4077 6613 4111 6647
rect 10793 6613 10827 6647
rect 23213 6613 23247 6647
rect 23581 6613 23615 6647
rect 3433 6409 3467 6443
rect 4997 6409 5031 6443
rect 8309 6409 8343 6443
rect 10701 6409 10735 6443
rect 14473 6409 14507 6443
rect 17969 6409 18003 6443
rect 19809 6409 19843 6443
rect 23305 6409 23339 6443
rect 23949 6409 23983 6443
rect 24317 6409 24351 6443
rect 2237 6341 2271 6375
rect 3341 6341 3375 6375
rect 1685 6273 1719 6307
rect 2605 6273 2639 6307
rect 2789 6273 2823 6307
rect 4259 6273 4293 6307
rect 5549 6273 5583 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7414 6273 7448 6307
rect 7573 6273 7607 6307
rect 8217 6273 8251 6307
rect 8493 6273 8527 6307
rect 8861 6273 8895 6307
rect 9919 6273 9953 6307
rect 11529 6273 11563 6307
rect 12725 6273 12759 6307
rect 13719 6303 13753 6337
rect 14933 6273 14967 6307
rect 15207 6273 15241 6307
rect 17693 6273 17727 6307
rect 19993 6273 20027 6307
rect 20269 6273 20303 6307
rect 20361 6273 20395 6307
rect 20821 6273 20855 6307
rect 20913 6273 20947 6307
rect 21189 6273 21223 6307
rect 21649 6273 21683 6307
rect 21833 6273 21867 6307
rect 22075 6273 22109 6307
rect 23213 6273 23247 6307
rect 23397 6273 23431 6307
rect 23673 6273 23707 6307
rect 23765 6273 23799 6307
rect 24041 6273 24075 6307
rect 24501 6273 24535 6307
rect 3985 6205 4019 6239
rect 7297 6205 7331 6239
rect 9045 6205 9079 6239
rect 9781 6205 9815 6239
rect 10057 6205 10091 6239
rect 11713 6205 11747 6239
rect 12449 6205 12483 6239
rect 12587 6205 12621 6239
rect 13461 6205 13495 6239
rect 17969 6205 18003 6239
rect 7021 6137 7055 6171
rect 9505 6137 9539 6171
rect 12173 6137 12207 6171
rect 13369 6137 13403 6171
rect 17785 6137 17819 6171
rect 20545 6137 20579 6171
rect 20637 6137 20671 6171
rect 21465 6137 21499 6171
rect 22845 6137 22879 6171
rect 1777 6069 1811 6103
rect 2881 6069 2915 6103
rect 5365 6069 5399 6103
rect 15945 6069 15979 6103
rect 20085 6069 20119 6103
rect 21097 6069 21131 6103
rect 21281 6069 21315 6103
rect 23489 6069 23523 6103
rect 24133 6069 24167 6103
rect 1593 5865 1627 5899
rect 2145 5865 2179 5899
rect 3249 5865 3283 5899
rect 5641 5865 5675 5899
rect 7113 5865 7147 5899
rect 8493 5865 8527 5899
rect 10885 5865 10919 5899
rect 18245 5865 18279 5899
rect 22937 5865 22971 5899
rect 12265 5797 12299 5831
rect 15945 5797 15979 5831
rect 20913 5797 20947 5831
rect 21465 5797 21499 5831
rect 23949 5797 23983 5831
rect 3985 5729 4019 5763
rect 6101 5729 6135 5763
rect 7481 5729 7515 5763
rect 15301 5729 15335 5763
rect 16221 5729 16255 5763
rect 16338 5729 16372 5763
rect 16497 5729 16531 5763
rect 19257 5729 19291 5763
rect 2605 5661 2639 5695
rect 3157 5661 3191 5695
rect 4259 5661 4293 5695
rect 5549 5661 5583 5695
rect 5825 5661 5859 5695
rect 6359 5631 6393 5665
rect 7755 5661 7789 5695
rect 9873 5661 9907 5695
rect 10147 5661 10181 5695
rect 11253 5661 11287 5695
rect 11527 5661 11561 5695
rect 15485 5661 15519 5695
rect 17233 5661 17267 5695
rect 17507 5661 17541 5695
rect 19499 5661 19533 5695
rect 20729 5661 20763 5695
rect 21005 5661 21039 5695
rect 21281 5637 21315 5671
rect 21557 5661 21591 5695
rect 23305 5661 23339 5695
rect 23673 5661 23707 5695
rect 23949 5661 23983 5695
rect 1501 5593 1535 5627
rect 2053 5593 2087 5627
rect 21802 5593 21836 5627
rect 2881 5525 2915 5559
rect 4997 5525 5031 5559
rect 5365 5525 5399 5559
rect 17141 5525 17175 5559
rect 20269 5525 20303 5559
rect 21189 5525 21223 5559
rect 6193 5321 6227 5355
rect 10241 5321 10275 5355
rect 17693 5321 17727 5355
rect 18153 5321 18187 5355
rect 18429 5321 18463 5355
rect 18613 5321 18647 5355
rect 24501 5321 24535 5355
rect 19533 5253 19567 5287
rect 1409 5185 1443 5219
rect 1667 5215 1701 5249
rect 3063 5185 3097 5219
rect 4353 5185 4387 5219
rect 5390 5185 5424 5219
rect 6377 5185 6411 5219
rect 6651 5185 6685 5219
rect 9503 5195 9537 5229
rect 12725 5185 12759 5219
rect 13645 5185 13679 5219
rect 13921 5185 13955 5219
rect 14657 5185 14691 5219
rect 15715 5185 15749 5219
rect 16955 5185 16989 5219
rect 18061 5185 18095 5219
rect 18337 5185 18371 5219
rect 18521 5185 18555 5219
rect 18797 5185 18831 5219
rect 19165 5185 19199 5219
rect 19349 5185 19383 5219
rect 19867 5185 19901 5219
rect 21189 5185 21223 5219
rect 21465 5185 21499 5219
rect 21557 5185 21591 5219
rect 22201 5185 22235 5219
rect 23388 5185 23422 5219
rect 2789 5117 2823 5151
rect 4537 5117 4571 5151
rect 4997 5117 5031 5151
rect 5273 5117 5307 5151
rect 5549 5117 5583 5151
rect 9229 5117 9263 5151
rect 12909 5117 12943 5151
rect 13783 5117 13817 5151
rect 14841 5117 14875 5151
rect 15577 5117 15611 5151
rect 15853 5117 15887 5151
rect 16681 5117 16715 5151
rect 19625 5117 19659 5151
rect 21005 5117 21039 5151
rect 22385 5117 22419 5151
rect 23121 5117 23155 5151
rect 13369 5049 13403 5083
rect 15301 5049 15335 5083
rect 19165 5049 19199 5083
rect 20637 5049 20671 5083
rect 2421 4981 2455 5015
rect 3801 4981 3835 5015
rect 7389 4981 7423 5015
rect 14565 4981 14599 5015
rect 16497 4981 16531 5015
rect 1501 4777 1535 4811
rect 3801 4777 3835 4811
rect 5549 4777 5583 4811
rect 13645 4777 13679 4811
rect 16405 4777 16439 4811
rect 19625 4777 19659 4811
rect 21281 4777 21315 4811
rect 24041 4777 24075 4811
rect 18797 4709 18831 4743
rect 18889 4709 18923 4743
rect 19349 4709 19383 4743
rect 19809 4709 19843 4743
rect 21005 4709 21039 4743
rect 22017 4709 22051 4743
rect 1961 4641 1995 4675
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 2835 4641 2869 4675
rect 12633 4641 12667 4675
rect 15393 4641 15427 4675
rect 17417 4641 17451 4675
rect 1685 4573 1719 4607
rect 1777 4573 1811 4607
rect 2973 4573 3007 4607
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 4537 4573 4571 4607
rect 4811 4573 4845 4607
rect 12907 4573 12941 4607
rect 15651 4543 15685 4577
rect 19073 4573 19107 4607
rect 19257 4573 19291 4607
rect 19533 4573 19567 4607
rect 19717 4573 19751 4607
rect 19993 4573 20027 4607
rect 20085 4573 20119 4607
rect 20269 4573 20303 4607
rect 20545 4573 20579 4607
rect 20821 4573 20855 4607
rect 20913 4573 20947 4607
rect 21189 4573 21223 4607
rect 21373 4573 21407 4607
rect 21649 4573 21683 4607
rect 21833 4573 21867 4607
rect 22293 4573 22327 4607
rect 22477 4573 22511 4607
rect 22751 4573 22785 4607
rect 17684 4505 17718 4539
rect 23949 4505 23983 4539
rect 3617 4437 3651 4471
rect 4077 4437 4111 4471
rect 20269 4437 20303 4471
rect 20361 4437 20395 4471
rect 20637 4437 20671 4471
rect 21465 4437 21499 4471
rect 22109 4437 22143 4471
rect 23489 4437 23523 4471
rect 15577 4233 15611 4267
rect 21465 4233 21499 4267
rect 1685 4165 1719 4199
rect 19257 4165 19291 4199
rect 24317 4165 24351 4199
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 3341 4097 3375 4131
rect 3479 4097 3513 4131
rect 3617 4097 3651 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 6745 4097 6779 4131
rect 7019 4097 7053 4131
rect 9321 4097 9355 4131
rect 10331 4097 10365 4131
rect 11529 4097 11563 4131
rect 11803 4097 11837 4131
rect 14565 4097 14599 4131
rect 14839 4097 14873 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 18797 4097 18831 4131
rect 19073 4097 19107 4131
rect 19901 4097 19935 4131
rect 20352 4097 20386 4131
rect 22385 4097 22419 4131
rect 22661 4097 22695 4131
rect 23029 4097 23063 4131
rect 24501 4097 24535 4131
rect 1961 4029 1995 4063
rect 2421 4029 2455 4063
rect 8125 4029 8159 4063
rect 8309 4029 8343 4063
rect 9045 4029 9079 4063
rect 9183 4029 9217 4063
rect 10057 4029 10091 4063
rect 20085 4029 20119 4063
rect 22017 4029 22051 4063
rect 23857 4029 23891 4063
rect 3065 3961 3099 3995
rect 8769 3961 8803 3995
rect 17693 3961 17727 3995
rect 18613 3961 18647 3995
rect 19717 3961 19751 3995
rect 22661 3961 22695 3995
rect 2145 3893 2179 3927
rect 4353 3893 4387 3927
rect 7757 3893 7791 3927
rect 9965 3893 9999 3927
rect 11069 3893 11103 3927
rect 12541 3893 12575 3927
rect 18337 3893 18371 3927
rect 18889 3893 18923 3927
rect 19349 3893 19383 3927
rect 1593 3689 1627 3723
rect 2145 3689 2179 3723
rect 2697 3689 2731 3723
rect 4905 3689 4939 3723
rect 15117 3689 15151 3723
rect 18245 3689 18279 3723
rect 20637 3689 20671 3723
rect 7205 3621 7239 3655
rect 8493 3621 8527 3655
rect 9597 3621 9631 3655
rect 13553 3621 13587 3655
rect 18521 3621 18555 3655
rect 23673 3621 23707 3655
rect 6929 3553 6963 3587
rect 7481 3553 7515 3587
rect 8953 3553 8987 3587
rect 9873 3553 9907 3587
rect 10011 3553 10045 3587
rect 21281 3553 21315 3587
rect 22661 3553 22695 3587
rect 1501 3485 1535 3519
rect 2513 3485 2547 3519
rect 5089 3485 5123 3519
rect 5363 3485 5397 3519
rect 7389 3485 7423 3519
rect 7755 3485 7789 3519
rect 9137 3485 9171 3519
rect 10149 3485 10183 3519
rect 11529 3485 11563 3519
rect 11805 3485 11839 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 14379 3485 14413 3519
rect 17233 3485 17267 3519
rect 17969 3485 18003 3519
rect 18061 3485 18095 3519
rect 18337 3485 18371 3519
rect 19257 3485 19291 3519
rect 19524 3485 19558 3519
rect 20821 3485 20855 3519
rect 21555 3485 21589 3519
rect 22935 3485 22969 3519
rect 24225 3485 24259 3519
rect 2053 3417 2087 3451
rect 4813 3417 4847 3451
rect 12081 3417 12115 3451
rect 12357 3417 12391 3451
rect 12449 3417 12483 3451
rect 12817 3417 12851 3451
rect 18705 3417 18739 3451
rect 19073 3417 19107 3451
rect 6101 3349 6135 3383
rect 10793 3349 10827 3383
rect 11345 3349 11379 3383
rect 11621 3349 11655 3383
rect 13185 3349 13219 3383
rect 13369 3349 13403 3383
rect 17049 3349 17083 3383
rect 17785 3349 17819 3383
rect 20913 3349 20947 3383
rect 22293 3349 22327 3383
rect 24041 3349 24075 3383
rect 1777 3145 1811 3179
rect 3341 3145 3375 3179
rect 3709 3145 3743 3179
rect 4537 3145 4571 3179
rect 6561 3145 6595 3179
rect 8033 3145 8067 3179
rect 11253 3145 11287 3179
rect 13185 3145 13219 3179
rect 18521 3145 18555 3179
rect 19165 3145 19199 3179
rect 24317 3145 24351 3179
rect 7665 3077 7699 3111
rect 9413 3077 9447 3111
rect 9965 3077 9999 3111
rect 10220 3077 10254 3111
rect 10333 3077 10367 3111
rect 11069 3077 11103 3111
rect 18705 3077 18739 3111
rect 21925 3077 21959 3111
rect 23090 3077 23124 3111
rect 1501 3009 1535 3043
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 3249 3009 3283 3043
rect 3525 3009 3559 3043
rect 4445 3009 4479 3043
rect 6837 3009 6871 3043
rect 6929 3009 6963 3043
rect 7297 3009 7331 3043
rect 8217 3009 8251 3043
rect 8493 3009 8527 3043
rect 9137 3009 9171 3043
rect 10701 3009 10735 3043
rect 11713 3009 11747 3043
rect 12081 3009 12115 3043
rect 12431 3039 12465 3073
rect 15669 3009 15703 3043
rect 16957 3009 16991 3043
rect 17417 3009 17451 3043
rect 17693 3009 17727 3043
rect 17969 3009 18003 3043
rect 18061 3009 18095 3043
rect 18337 3009 18371 3043
rect 19349 3009 19383 3043
rect 20821 3009 20855 3043
rect 22477 3009 22511 3043
rect 22845 3009 22879 3043
rect 24501 3009 24535 3043
rect 12173 2941 12207 2975
rect 19533 2941 19567 2975
rect 19809 2941 19843 2975
rect 21005 2941 21039 2975
rect 1685 2873 1719 2907
rect 7849 2873 7883 2907
rect 24225 2873 24259 2907
rect 2053 2805 2087 2839
rect 8309 2805 8343 2839
rect 8953 2805 8987 2839
rect 11529 2805 11563 2839
rect 11897 2805 11931 2839
rect 15485 2805 15519 2839
rect 17233 2805 17267 2839
rect 17509 2805 17543 2839
rect 17785 2805 17819 2839
rect 18245 2805 18279 2839
rect 18797 2805 18831 2839
rect 22017 2805 22051 2839
rect 22569 2805 22603 2839
rect 1961 2601 1995 2635
rect 3249 2601 3283 2635
rect 3985 2601 4019 2635
rect 4721 2601 4755 2635
rect 6837 2601 6871 2635
rect 10885 2601 10919 2635
rect 13277 2601 13311 2635
rect 14933 2601 14967 2635
rect 16681 2601 16715 2635
rect 16773 2601 16807 2635
rect 23213 2601 23247 2635
rect 1685 2533 1719 2567
rect 5549 2533 5583 2567
rect 11621 2533 11655 2567
rect 13369 2533 13403 2567
rect 23857 2533 23891 2567
rect 5825 2465 5859 2499
rect 9873 2465 9907 2499
rect 16405 2465 16439 2499
rect 21097 2465 21131 2499
rect 21833 2465 21867 2499
rect 23489 2465 23523 2499
rect 24041 2465 24075 2499
rect 1777 2397 1811 2431
rect 2237 2397 2271 2431
rect 2511 2397 2545 2431
rect 3801 2397 3835 2431
rect 4537 2397 4571 2431
rect 4997 2397 5031 2431
rect 5457 2397 5491 2431
rect 5733 2397 5767 2431
rect 6099 2397 6133 2431
rect 7573 2397 7607 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 8309 2397 8343 2431
rect 8769 2397 8803 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 10147 2397 10181 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 12081 2397 12115 2431
rect 12449 2397 12483 2431
rect 12909 2397 12943 2431
rect 13553 2397 13587 2431
rect 13829 2397 13863 2431
rect 15393 2397 15427 2431
rect 15669 2397 15703 2431
rect 15945 2397 15979 2431
rect 16497 2397 16531 2431
rect 16957 2397 16991 2431
rect 17233 2397 17267 2431
rect 18705 2397 18739 2431
rect 19441 2397 19475 2431
rect 20637 2397 20671 2431
rect 21741 2397 21775 2431
rect 23397 2397 23431 2431
rect 23581 2397 23615 2431
rect 23857 2397 23891 2431
rect 1501 2329 1535 2363
rect 17601 2329 17635 2363
rect 18153 2329 18187 2363
rect 20177 2329 20211 2363
rect 22078 2329 22112 2363
rect 24225 2329 24259 2363
rect 4813 2261 4847 2295
rect 5273 2261 5307 2295
rect 7389 2261 7423 2295
rect 7665 2261 7699 2295
rect 7941 2261 7975 2295
rect 8401 2261 8435 2295
rect 8585 2261 8619 2295
rect 8953 2261 8987 2295
rect 9505 2261 9539 2295
rect 11345 2261 11379 2295
rect 11897 2261 11931 2295
rect 12725 2261 12759 2295
rect 13645 2261 13679 2295
rect 15209 2261 15243 2295
rect 15485 2261 15519 2295
rect 15761 2261 15795 2295
rect 17049 2261 17083 2295
rect 17693 2261 17727 2295
rect 18245 2261 18279 2295
rect 18797 2261 18831 2295
rect 21557 2261 21591 2295
rect 1593 2057 1627 2091
rect 2697 2057 2731 2091
rect 4261 2057 4295 2091
rect 4997 2057 5031 2091
rect 5365 2057 5399 2091
rect 6837 2057 6871 2091
rect 7573 2057 7607 2091
rect 9137 2057 9171 2091
rect 10517 2057 10551 2091
rect 15209 2057 15243 2091
rect 18337 2057 18371 2091
rect 22385 2057 22419 2091
rect 5641 1989 5675 2023
rect 5825 1989 5859 2023
rect 6009 1989 6043 2023
rect 11805 1989 11839 2023
rect 12357 1989 12391 2023
rect 17325 1989 17359 2023
rect 17877 1989 17911 2023
rect 21465 1989 21499 2023
rect 22753 1989 22787 2023
rect 24317 1989 24351 2023
rect 1409 1921 1443 1955
rect 1685 1921 1719 1955
rect 1943 1951 1977 1985
rect 3433 1921 3467 1955
rect 3709 1921 3743 1955
rect 3801 1921 3835 1955
rect 4169 1921 4203 1955
rect 4445 1921 4479 1955
rect 4813 1921 4847 1955
rect 5273 1921 5307 1955
rect 6193 1921 6227 1955
rect 6561 1921 6595 1955
rect 6653 1921 6687 1955
rect 7113 1921 7147 1955
rect 7481 1921 7515 1955
rect 7849 1921 7883 1955
rect 8033 1921 8067 1955
rect 8125 1921 8159 1955
rect 8399 1921 8433 1955
rect 9779 1921 9813 1955
rect 10977 1921 11011 1955
rect 13093 1921 13127 1955
rect 13553 1921 13587 1955
rect 13829 1921 13863 1955
rect 14289 1921 14323 1955
rect 14473 1921 14507 1955
rect 14841 1921 14875 1955
rect 15393 1921 15427 1955
rect 15669 1921 15703 1955
rect 16129 1921 16163 1955
rect 16773 1921 16807 1955
rect 18521 1921 18555 1955
rect 19717 1921 19751 1955
rect 20821 1921 20855 1955
rect 21925 1921 21959 1955
rect 22201 1921 22235 1955
rect 9505 1853 9539 1887
rect 18613 1853 18647 1887
rect 18889 1853 18923 1887
rect 19901 1853 19935 1887
rect 3985 1785 4019 1819
rect 6377 1785 6411 1819
rect 7297 1785 7331 1819
rect 13369 1785 13403 1819
rect 14105 1785 14139 1819
rect 3249 1717 3283 1751
rect 3525 1717 3559 1751
rect 4629 1717 4663 1751
rect 11069 1717 11103 1751
rect 11897 1717 11931 1751
rect 12633 1717 12667 1751
rect 13645 1717 13679 1751
rect 14657 1717 14691 1751
rect 15025 1717 15059 1751
rect 15761 1717 15795 1751
rect 16313 1717 16347 1751
rect 16865 1717 16899 1751
rect 17417 1717 17451 1751
rect 17969 1717 18003 1751
rect 22017 1717 22051 1751
rect 2789 1513 2823 1547
rect 4169 1513 4203 1547
rect 14289 1513 14323 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 16865 1513 16899 1547
rect 17417 1513 17451 1547
rect 18521 1513 18555 1547
rect 23121 1513 23155 1547
rect 23857 1513 23891 1547
rect 8953 1445 8987 1479
rect 13645 1445 13679 1479
rect 18061 1445 18095 1479
rect 18889 1445 18923 1479
rect 20545 1445 20579 1479
rect 9965 1377 9999 1411
rect 11253 1377 11287 1411
rect 12541 1377 12575 1411
rect 1409 1309 1443 1343
rect 1685 1309 1719 1343
rect 4905 1309 4939 1343
rect 5273 1309 5307 1343
rect 5549 1309 5583 1343
rect 6561 1309 6595 1343
rect 7389 1309 7423 1343
rect 7757 1309 7791 1343
rect 8125 1309 8159 1343
rect 8493 1309 8527 1343
rect 9137 1309 9171 1343
rect 9413 1309 9447 1343
rect 9689 1309 9723 1343
rect 10425 1309 10459 1343
rect 10977 1309 11011 1343
rect 11713 1309 11747 1343
rect 11805 1309 11839 1343
rect 12909 1309 12943 1343
rect 13277 1309 13311 1343
rect 13829 1309 13863 1343
rect 14657 1309 14691 1343
rect 15301 1309 15335 1343
rect 15853 1309 15887 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 17325 1309 17359 1343
rect 17877 1309 17911 1343
rect 18429 1309 18463 1343
rect 19073 1309 19107 1343
rect 21649 1309 21683 1343
rect 23673 1309 23707 1343
rect 23949 1309 23983 1343
rect 24133 1309 24167 1343
rect 2329 1241 2363 1275
rect 2513 1241 2547 1275
rect 2697 1241 2731 1275
rect 3065 1241 3099 1275
rect 3433 1241 3467 1275
rect 3617 1241 3651 1275
rect 3893 1241 3927 1275
rect 4629 1241 4663 1275
rect 6745 1241 6779 1275
rect 6929 1241 6963 1275
rect 7113 1241 7147 1275
rect 12265 1241 12299 1275
rect 14197 1241 14231 1275
rect 19257 1241 19291 1275
rect 21189 1241 21223 1275
rect 21373 1241 21407 1275
rect 21833 1241 21867 1275
rect 1593 1173 1627 1207
rect 1869 1173 1903 1207
rect 3157 1173 3191 1207
rect 4721 1173 4755 1207
rect 5089 1173 5123 1207
rect 6377 1173 6411 1207
rect 7205 1173 7239 1207
rect 7573 1173 7607 1207
rect 7941 1173 7975 1207
rect 8309 1173 8343 1207
rect 8677 1173 8711 1207
rect 10517 1173 10551 1207
rect 11529 1173 11563 1207
rect 11989 1173 12023 1207
rect 13093 1173 13127 1207
rect 13461 1173 13495 1207
rect 14841 1173 14875 1207
rect 21465 1173 21499 1207
rect 24133 1173 24167 1207
<< metal1 >>
rect 18138 43800 18144 43852
rect 18196 43840 18202 43852
rect 21266 43840 21272 43852
rect 18196 43812 21272 43840
rect 18196 43800 18202 43812
rect 21266 43800 21272 43812
rect 21324 43800 21330 43852
rect 21726 43800 21732 43852
rect 21784 43840 21790 43852
rect 22922 43840 22928 43852
rect 21784 43812 22928 43840
rect 21784 43800 21790 43812
rect 22922 43800 22928 43812
rect 22980 43800 22986 43852
rect 20714 43732 20720 43784
rect 20772 43772 20778 43784
rect 22554 43772 22560 43784
rect 20772 43744 22560 43772
rect 20772 43732 20778 43744
rect 22554 43732 22560 43744
rect 22612 43732 22618 43784
rect 5258 43664 5264 43716
rect 5316 43704 5322 43716
rect 16022 43704 16028 43716
rect 5316 43676 16028 43704
rect 5316 43664 5322 43676
rect 16022 43664 16028 43676
rect 16080 43664 16086 43716
rect 18506 43664 18512 43716
rect 18564 43704 18570 43716
rect 20990 43704 20996 43716
rect 18564 43676 20996 43704
rect 18564 43664 18570 43676
rect 20990 43664 20996 43676
rect 21048 43664 21054 43716
rect 3602 43596 3608 43648
rect 3660 43636 3666 43648
rect 10502 43636 10508 43648
rect 3660 43608 10508 43636
rect 3660 43596 3666 43608
rect 10502 43596 10508 43608
rect 10560 43596 10566 43648
rect 17494 43596 17500 43648
rect 17552 43636 17558 43648
rect 22370 43636 22376 43648
rect 17552 43608 22376 43636
rect 17552 43596 17558 43608
rect 22370 43596 22376 43608
rect 22428 43596 22434 43648
rect 1104 43546 25000 43568
rect 1104 43494 6884 43546
rect 6936 43494 6948 43546
rect 7000 43494 7012 43546
rect 7064 43494 7076 43546
rect 7128 43494 7140 43546
rect 7192 43494 12818 43546
rect 12870 43494 12882 43546
rect 12934 43494 12946 43546
rect 12998 43494 13010 43546
rect 13062 43494 13074 43546
rect 13126 43494 18752 43546
rect 18804 43494 18816 43546
rect 18868 43494 18880 43546
rect 18932 43494 18944 43546
rect 18996 43494 19008 43546
rect 19060 43494 24686 43546
rect 24738 43494 24750 43546
rect 24802 43494 24814 43546
rect 24866 43494 24878 43546
rect 24930 43494 24942 43546
rect 24994 43494 25000 43546
rect 1104 43472 25000 43494
rect 1854 43392 1860 43444
rect 1912 43392 1918 43444
rect 2777 43435 2835 43441
rect 2777 43401 2789 43435
rect 2823 43432 2835 43435
rect 2958 43432 2964 43444
rect 2823 43404 2964 43432
rect 2823 43401 2835 43404
rect 2777 43395 2835 43401
rect 2958 43392 2964 43404
rect 3016 43392 3022 43444
rect 3145 43435 3203 43441
rect 3145 43401 3157 43435
rect 3191 43401 3203 43435
rect 3145 43395 3203 43401
rect 382 43324 388 43376
rect 440 43364 446 43376
rect 3160 43364 3188 43395
rect 4338 43392 4344 43444
rect 4396 43432 4402 43444
rect 4617 43435 4675 43441
rect 4617 43432 4629 43435
rect 4396 43404 4629 43432
rect 4396 43392 4402 43404
rect 4617 43401 4629 43404
rect 4663 43401 4675 43435
rect 4617 43395 4675 43401
rect 5534 43392 5540 43444
rect 5592 43392 5598 43444
rect 6089 43435 6147 43441
rect 6089 43401 6101 43435
rect 6135 43432 6147 43435
rect 6270 43432 6276 43444
rect 6135 43404 6276 43432
rect 6135 43401 6147 43404
rect 6089 43395 6147 43401
rect 6270 43392 6276 43404
rect 6328 43392 6334 43444
rect 6365 43435 6423 43441
rect 6365 43401 6377 43435
rect 6411 43401 6423 43435
rect 6365 43395 6423 43401
rect 6380 43364 6408 43395
rect 6638 43392 6644 43444
rect 6696 43432 6702 43444
rect 7009 43435 7067 43441
rect 7009 43432 7021 43435
rect 6696 43404 7021 43432
rect 6696 43392 6702 43404
rect 7009 43401 7021 43404
rect 7055 43401 7067 43435
rect 7009 43395 7067 43401
rect 7377 43435 7435 43441
rect 7377 43401 7389 43435
rect 7423 43432 7435 43435
rect 7650 43432 7656 43444
rect 7423 43404 7656 43432
rect 7423 43401 7435 43404
rect 7377 43395 7435 43401
rect 7650 43392 7656 43404
rect 7708 43392 7714 43444
rect 7745 43435 7803 43441
rect 7745 43401 7757 43435
rect 7791 43432 7803 43435
rect 7926 43432 7932 43444
rect 7791 43404 7932 43432
rect 7791 43401 7803 43404
rect 7745 43395 7803 43401
rect 7926 43392 7932 43404
rect 7984 43392 7990 43444
rect 8297 43435 8355 43441
rect 8297 43401 8309 43435
rect 8343 43432 8355 43435
rect 8478 43432 8484 43444
rect 8343 43404 8484 43432
rect 8343 43401 8355 43404
rect 8297 43395 8355 43401
rect 8478 43392 8484 43404
rect 8536 43392 8542 43444
rect 8665 43435 8723 43441
rect 8665 43401 8677 43435
rect 8711 43432 8723 43435
rect 9030 43432 9036 43444
rect 8711 43404 9036 43432
rect 8711 43401 8723 43404
rect 8665 43395 8723 43401
rect 9030 43392 9036 43404
rect 9088 43392 9094 43444
rect 9217 43435 9275 43441
rect 9217 43401 9229 43435
rect 9263 43432 9275 43435
rect 9582 43432 9588 43444
rect 9263 43404 9588 43432
rect 9263 43401 9275 43404
rect 9217 43395 9275 43401
rect 9582 43392 9588 43404
rect 9640 43392 9646 43444
rect 9769 43435 9827 43441
rect 9769 43401 9781 43435
rect 9815 43432 9827 43435
rect 9858 43432 9864 43444
rect 9815 43404 9864 43432
rect 9815 43401 9827 43404
rect 9769 43395 9827 43401
rect 9858 43392 9864 43404
rect 9916 43392 9922 43444
rect 10502 43392 10508 43444
rect 10560 43392 10566 43444
rect 12253 43435 12311 43441
rect 12253 43401 12265 43435
rect 12299 43432 12311 43435
rect 13998 43432 14004 43444
rect 12299 43404 14004 43432
rect 12299 43401 12311 43404
rect 12253 43395 12311 43401
rect 13998 43392 14004 43404
rect 14056 43392 14062 43444
rect 17034 43392 17040 43444
rect 17092 43432 17098 43444
rect 17092 43404 18000 43432
rect 17092 43392 17098 43404
rect 6733 43367 6791 43373
rect 6733 43364 6745 43367
rect 440 43336 3188 43364
rect 3896 43336 6224 43364
rect 6380 43336 6745 43364
rect 440 43324 446 43336
rect 658 43256 664 43308
rect 716 43296 722 43308
rect 1581 43299 1639 43305
rect 1581 43296 1593 43299
rect 716 43268 1593 43296
rect 716 43256 722 43268
rect 1581 43265 1593 43268
rect 1627 43265 1639 43299
rect 1581 43259 1639 43265
rect 1765 43299 1823 43305
rect 1765 43265 1777 43299
rect 1811 43265 1823 43299
rect 1765 43259 1823 43265
rect 1780 43228 1808 43259
rect 2498 43256 2504 43308
rect 2556 43256 2562 43308
rect 3053 43299 3111 43305
rect 3053 43265 3065 43299
rect 3099 43296 3111 43299
rect 3896 43296 3924 43336
rect 3099 43268 3924 43296
rect 3973 43299 4031 43305
rect 3099 43265 3111 43268
rect 3053 43259 3111 43265
rect 3973 43265 3985 43299
rect 4019 43296 4031 43299
rect 4338 43296 4344 43308
rect 4019 43268 4344 43296
rect 4019 43265 4031 43268
rect 3973 43259 4031 43265
rect 4338 43256 4344 43268
rect 4396 43256 4402 43308
rect 4525 43299 4583 43305
rect 4525 43265 4537 43299
rect 4571 43265 4583 43299
rect 4525 43259 4583 43265
rect 5261 43299 5319 43305
rect 5261 43265 5273 43299
rect 5307 43296 5319 43299
rect 5442 43296 5448 43308
rect 5307 43268 5448 43296
rect 5307 43265 5319 43268
rect 5261 43259 5319 43265
rect 2958 43228 2964 43240
rect 1780 43200 2964 43228
rect 2958 43188 2964 43200
rect 3016 43188 3022 43240
rect 4246 43188 4252 43240
rect 4304 43228 4310 43240
rect 4540 43228 4568 43259
rect 5442 43256 5448 43268
rect 5500 43256 5506 43308
rect 5534 43256 5540 43308
rect 5592 43296 5598 43308
rect 5905 43299 5963 43305
rect 5905 43296 5917 43299
rect 5592 43268 5917 43296
rect 5592 43256 5598 43268
rect 5905 43265 5917 43268
rect 5951 43265 5963 43299
rect 5905 43259 5963 43265
rect 4304 43200 4568 43228
rect 4304 43188 4310 43200
rect 3789 43163 3847 43169
rect 3789 43129 3801 43163
rect 3835 43160 3847 43163
rect 4706 43160 4712 43172
rect 3835 43132 4712 43160
rect 3835 43129 3847 43132
rect 3789 43123 3847 43129
rect 4706 43120 4712 43132
rect 4764 43120 4770 43172
rect 1397 43095 1455 43101
rect 1397 43061 1409 43095
rect 1443 43092 1455 43095
rect 1762 43092 1768 43104
rect 1443 43064 1768 43092
rect 1443 43061 1455 43064
rect 1397 43055 1455 43061
rect 1762 43052 1768 43064
rect 1820 43052 1826 43104
rect 4341 43095 4399 43101
rect 4341 43061 4353 43095
rect 4387 43092 4399 43095
rect 4430 43092 4436 43104
rect 4387 43064 4436 43092
rect 4387 43061 4399 43064
rect 4341 43055 4399 43061
rect 4430 43052 4436 43064
rect 4488 43052 4494 43104
rect 6196 43092 6224 43336
rect 6733 43333 6745 43336
rect 6779 43333 6791 43367
rect 6733 43327 6791 43333
rect 8021 43367 8079 43373
rect 8021 43333 8033 43367
rect 8067 43364 8079 43367
rect 8938 43364 8944 43376
rect 8067 43336 8944 43364
rect 8067 43333 8079 43336
rect 8021 43327 8079 43333
rect 8938 43324 8944 43336
rect 8996 43324 9002 43376
rect 9398 43324 9404 43376
rect 9456 43364 9462 43376
rect 11146 43364 11152 43376
rect 9456 43336 11152 43364
rect 9456 43324 9462 43336
rect 11146 43324 11152 43336
rect 11204 43324 11210 43376
rect 12434 43324 12440 43376
rect 12492 43324 12498 43376
rect 12802 43324 12808 43376
rect 12860 43324 12866 43376
rect 13354 43324 13360 43376
rect 13412 43364 13418 43376
rect 14185 43367 14243 43373
rect 14185 43364 14197 43367
rect 13412 43336 14197 43364
rect 13412 43324 13418 43336
rect 14185 43333 14197 43336
rect 14231 43333 14243 43367
rect 14185 43327 14243 43333
rect 14734 43324 14740 43376
rect 14792 43324 14798 43376
rect 14826 43324 14832 43376
rect 14884 43364 14890 43376
rect 15105 43367 15163 43373
rect 15105 43364 15117 43367
rect 14884 43336 15117 43364
rect 14884 43324 14890 43336
rect 15105 43333 15117 43336
rect 15151 43333 15163 43367
rect 15105 43327 15163 43333
rect 15930 43324 15936 43376
rect 15988 43364 15994 43376
rect 16301 43367 16359 43373
rect 16301 43364 16313 43367
rect 15988 43336 16313 43364
rect 15988 43324 15994 43336
rect 16301 43333 16313 43336
rect 16347 43333 16359 43367
rect 16301 43327 16359 43333
rect 16390 43324 16396 43376
rect 16448 43364 16454 43376
rect 16761 43367 16819 43373
rect 16761 43364 16773 43367
rect 16448 43336 16773 43364
rect 16448 43324 16454 43336
rect 16761 43333 16773 43336
rect 16807 43333 16819 43367
rect 16761 43327 16819 43333
rect 16850 43324 16856 43376
rect 16908 43364 16914 43376
rect 16908 43336 17816 43364
rect 16908 43324 16914 43336
rect 6270 43256 6276 43308
rect 6328 43296 6334 43308
rect 6549 43299 6607 43305
rect 6549 43296 6561 43299
rect 6328 43268 6561 43296
rect 6328 43256 6334 43268
rect 6549 43265 6561 43268
rect 6595 43265 6607 43299
rect 6549 43259 6607 43265
rect 7193 43299 7251 43305
rect 7193 43265 7205 43299
rect 7239 43296 7251 43299
rect 7282 43296 7288 43308
rect 7239 43268 7288 43296
rect 7239 43265 7251 43268
rect 7193 43259 7251 43265
rect 7282 43256 7288 43268
rect 7340 43256 7346 43308
rect 7561 43299 7619 43305
rect 7561 43265 7573 43299
rect 7607 43265 7619 43299
rect 7561 43259 7619 43265
rect 8481 43299 8539 43305
rect 8481 43265 8493 43299
rect 8527 43265 8539 43299
rect 8481 43259 8539 43265
rect 9033 43299 9091 43305
rect 9033 43265 9045 43299
rect 9079 43265 9091 43299
rect 9033 43259 9091 43265
rect 7576 43228 7604 43259
rect 8110 43228 8116 43240
rect 7576 43200 8116 43228
rect 8110 43188 8116 43200
rect 8168 43188 8174 43240
rect 8496 43160 8524 43259
rect 9048 43228 9076 43259
rect 9490 43256 9496 43308
rect 9548 43256 9554 43308
rect 9950 43256 9956 43308
rect 10008 43256 10014 43308
rect 10318 43256 10324 43308
rect 10376 43256 10382 43308
rect 10686 43256 10692 43308
rect 10744 43256 10750 43308
rect 11054 43256 11060 43308
rect 11112 43256 11118 43308
rect 11238 43256 11244 43308
rect 11296 43296 11302 43308
rect 11517 43299 11575 43305
rect 11517 43296 11529 43299
rect 11296 43268 11529 43296
rect 11296 43256 11302 43268
rect 11517 43265 11529 43268
rect 11563 43265 11575 43299
rect 11517 43259 11575 43265
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 13630 43256 13636 43308
rect 13688 43256 13694 43308
rect 15470 43256 15476 43308
rect 15528 43256 15534 43308
rect 15838 43256 15844 43308
rect 15896 43256 15902 43308
rect 16022 43256 16028 43308
rect 16080 43296 16086 43308
rect 16485 43299 16543 43305
rect 16485 43296 16497 43299
rect 16080 43268 16497 43296
rect 16080 43256 16086 43268
rect 16485 43265 16497 43268
rect 16531 43265 16543 43299
rect 16485 43259 16543 43265
rect 17402 43256 17408 43308
rect 17460 43296 17466 43308
rect 17788 43305 17816 43336
rect 17497 43299 17555 43305
rect 17497 43296 17509 43299
rect 17460 43268 17509 43296
rect 17460 43256 17466 43268
rect 17497 43265 17509 43268
rect 17543 43265 17555 43299
rect 17497 43259 17555 43265
rect 17773 43299 17831 43305
rect 17773 43265 17785 43299
rect 17819 43265 17831 43299
rect 17972 43296 18000 43404
rect 18138 43392 18144 43444
rect 18196 43432 18202 43444
rect 20073 43435 20131 43441
rect 18196 43404 19472 43432
rect 18196 43392 18202 43404
rect 18230 43324 18236 43376
rect 18288 43364 18294 43376
rect 18288 43336 18644 43364
rect 18288 43324 18294 43336
rect 18616 43305 18644 43336
rect 18049 43299 18107 43305
rect 18049 43296 18061 43299
rect 17972 43268 18061 43296
rect 17773 43259 17831 43265
rect 18049 43265 18061 43268
rect 18095 43265 18107 43299
rect 18049 43259 18107 43265
rect 18325 43299 18383 43305
rect 18325 43265 18337 43299
rect 18371 43265 18383 43299
rect 18325 43259 18383 43265
rect 18601 43299 18659 43305
rect 18601 43265 18613 43299
rect 18647 43265 18659 43299
rect 18601 43259 18659 43265
rect 18877 43299 18935 43305
rect 18877 43265 18889 43299
rect 18923 43296 18935 43299
rect 19334 43296 19340 43308
rect 18923 43268 19340 43296
rect 18923 43265 18935 43268
rect 18877 43259 18935 43265
rect 9674 43228 9680 43240
rect 9048 43200 9680 43228
rect 9674 43188 9680 43200
rect 9732 43188 9738 43240
rect 17310 43188 17316 43240
rect 17368 43228 17374 43240
rect 18340 43228 18368 43259
rect 19334 43256 19340 43268
rect 19392 43256 19398 43308
rect 19444 43305 19472 43404
rect 20073 43401 20085 43435
rect 20119 43432 20131 43435
rect 20346 43432 20352 43444
rect 20119 43404 20352 43432
rect 20119 43401 20131 43404
rect 20073 43395 20131 43401
rect 20346 43392 20352 43404
rect 20404 43392 20410 43444
rect 20622 43392 20628 43444
rect 20680 43432 20686 43444
rect 20993 43435 21051 43441
rect 20993 43432 21005 43435
rect 20680 43404 21005 43432
rect 20680 43392 20686 43404
rect 20993 43401 21005 43404
rect 21039 43401 21051 43435
rect 20993 43395 21051 43401
rect 21174 43392 21180 43444
rect 21232 43432 21238 43444
rect 22005 43435 22063 43441
rect 22005 43432 22017 43435
rect 21232 43404 22017 43432
rect 21232 43392 21238 43404
rect 22005 43401 22017 43404
rect 22051 43401 22063 43435
rect 22373 43435 22431 43441
rect 22373 43432 22385 43435
rect 22005 43395 22063 43401
rect 22204 43404 22385 43432
rect 20530 43324 20536 43376
rect 20588 43364 20594 43376
rect 20588 43336 21404 43364
rect 20588 43324 20594 43336
rect 19429 43299 19487 43305
rect 19429 43265 19441 43299
rect 19475 43265 19487 43299
rect 19429 43259 19487 43265
rect 19705 43299 19763 43305
rect 19705 43265 19717 43299
rect 19751 43265 19763 43299
rect 19705 43259 19763 43265
rect 17368 43200 18368 43228
rect 19720 43228 19748 43259
rect 19886 43256 19892 43308
rect 19944 43256 19950 43308
rect 20349 43299 20407 43305
rect 20349 43265 20361 43299
rect 20395 43265 20407 43299
rect 20349 43259 20407 43265
rect 19978 43228 19984 43240
rect 19720 43200 19984 43228
rect 17368 43188 17374 43200
rect 19978 43188 19984 43200
rect 20036 43188 20042 43240
rect 20364 43228 20392 43259
rect 20622 43256 20628 43308
rect 20680 43296 20686 43308
rect 21376 43305 21404 43336
rect 21542 43324 21548 43376
rect 21600 43364 21606 43376
rect 22204 43364 22232 43404
rect 22373 43401 22385 43404
rect 22419 43401 22431 43435
rect 22373 43395 22431 43401
rect 22922 43392 22928 43444
rect 22980 43392 22986 43444
rect 23106 43392 23112 43444
rect 23164 43432 23170 43444
rect 23477 43435 23535 43441
rect 23477 43432 23489 43435
rect 23164 43404 23489 43432
rect 23164 43392 23170 43404
rect 23477 43401 23489 43404
rect 23523 43401 23535 43435
rect 23477 43395 23535 43401
rect 23014 43364 23020 43376
rect 21600 43336 22232 43364
rect 22388 43336 23020 43364
rect 21600 43324 21606 43336
rect 20901 43299 20959 43305
rect 20901 43296 20913 43299
rect 20680 43268 20913 43296
rect 20680 43256 20686 43268
rect 20901 43265 20913 43268
rect 20947 43265 20959 43299
rect 20901 43259 20959 43265
rect 21361 43299 21419 43305
rect 21361 43265 21373 43299
rect 21407 43265 21419 43299
rect 21361 43259 21419 43265
rect 21634 43256 21640 43308
rect 21692 43296 21698 43308
rect 21821 43299 21879 43305
rect 21821 43296 21833 43299
rect 21692 43268 21833 43296
rect 21692 43256 21698 43268
rect 21821 43265 21833 43268
rect 21867 43265 21879 43299
rect 21821 43259 21879 43265
rect 22281 43299 22339 43305
rect 22281 43265 22293 43299
rect 22327 43296 22339 43299
rect 22388 43296 22416 43336
rect 23014 43324 23020 43336
rect 23072 43324 23078 43376
rect 22327 43268 22416 43296
rect 22327 43265 22339 43268
rect 22281 43259 22339 43265
rect 22462 43256 22468 43308
rect 22520 43296 22526 43308
rect 22833 43299 22891 43305
rect 22833 43296 22845 43299
rect 22520 43268 22845 43296
rect 22520 43256 22526 43268
rect 22833 43265 22845 43268
rect 22879 43265 22891 43299
rect 22833 43259 22891 43265
rect 22922 43256 22928 43308
rect 22980 43296 22986 43308
rect 23385 43299 23443 43305
rect 23385 43296 23397 43299
rect 22980 43268 23397 43296
rect 22980 43256 22986 43268
rect 23385 43265 23397 43268
rect 23431 43265 23443 43299
rect 23385 43259 23443 43265
rect 23937 43299 23995 43305
rect 23937 43265 23949 43299
rect 23983 43265 23995 43299
rect 23937 43259 23995 43265
rect 22186 43228 22192 43240
rect 20364 43200 22192 43228
rect 22186 43188 22192 43200
rect 22244 43188 22250 43240
rect 22646 43188 22652 43240
rect 22704 43228 22710 43240
rect 23952 43228 23980 43259
rect 22704 43200 23980 43228
rect 22704 43188 22710 43200
rect 10594 43160 10600 43172
rect 8496 43132 10600 43160
rect 10594 43120 10600 43132
rect 10652 43120 10658 43172
rect 13630 43120 13636 43172
rect 13688 43160 13694 43172
rect 13688 43132 14412 43160
rect 13688 43120 13694 43132
rect 9766 43092 9772 43104
rect 6196 43064 9772 43092
rect 9766 43052 9772 43064
rect 9824 43052 9830 43104
rect 10134 43052 10140 43104
rect 10192 43052 10198 43104
rect 10873 43095 10931 43101
rect 10873 43061 10885 43095
rect 10919 43092 10931 43095
rect 10962 43092 10968 43104
rect 10919 43064 10968 43092
rect 10919 43061 10931 43064
rect 10873 43055 10931 43061
rect 10962 43052 10968 43064
rect 11020 43052 11026 43104
rect 11238 43052 11244 43104
rect 11296 43052 11302 43104
rect 11701 43095 11759 43101
rect 11701 43061 11713 43095
rect 11747 43092 11759 43095
rect 11974 43092 11980 43104
rect 11747 43064 11980 43092
rect 11747 43061 11759 43064
rect 11701 43055 11759 43061
rect 11974 43052 11980 43064
rect 12032 43052 12038 43104
rect 12526 43052 12532 43104
rect 12584 43052 12590 43104
rect 12894 43052 12900 43104
rect 12952 43052 12958 43104
rect 13817 43095 13875 43101
rect 13817 43061 13829 43095
rect 13863 43092 13875 43095
rect 14182 43092 14188 43104
rect 13863 43064 14188 43092
rect 13863 43061 13875 43064
rect 13817 43055 13875 43061
rect 14182 43052 14188 43064
rect 14240 43052 14246 43104
rect 14274 43052 14280 43104
rect 14332 43052 14338 43104
rect 14384 43092 14412 43132
rect 14918 43120 14924 43172
rect 14976 43120 14982 43172
rect 17865 43163 17923 43169
rect 17865 43160 17877 43163
rect 17696 43132 17877 43160
rect 17696 43104 17724 43132
rect 17865 43129 17877 43132
rect 17911 43129 17923 43163
rect 17865 43123 17923 43129
rect 18322 43120 18328 43172
rect 18380 43160 18386 43172
rect 19245 43163 19303 43169
rect 19245 43160 19257 43163
rect 18380 43132 19257 43160
rect 18380 43120 18386 43132
rect 19245 43129 19257 43132
rect 19291 43129 19303 43163
rect 19245 43123 19303 43129
rect 20625 43163 20683 43169
rect 20625 43129 20637 43163
rect 20671 43160 20683 43163
rect 20714 43160 20720 43172
rect 20671 43132 20720 43160
rect 20671 43129 20683 43132
rect 20625 43123 20683 43129
rect 20714 43120 20720 43132
rect 20772 43120 20778 43172
rect 20898 43120 20904 43172
rect 20956 43160 20962 43172
rect 21545 43163 21603 43169
rect 21545 43160 21557 43163
rect 20956 43132 21557 43160
rect 20956 43120 20962 43132
rect 21545 43129 21557 43132
rect 21591 43129 21603 43163
rect 21545 43123 21603 43129
rect 15197 43095 15255 43101
rect 15197 43092 15209 43095
rect 14384 43064 15209 43092
rect 15197 43061 15209 43064
rect 15243 43061 15255 43095
rect 15197 43055 15255 43061
rect 15286 43052 15292 43104
rect 15344 43092 15350 43104
rect 15657 43095 15715 43101
rect 15657 43092 15669 43095
rect 15344 43064 15669 43092
rect 15344 43052 15350 43064
rect 15657 43061 15669 43064
rect 15703 43061 15715 43095
rect 15657 43055 15715 43061
rect 15838 43052 15844 43104
rect 15896 43092 15902 43104
rect 16025 43095 16083 43101
rect 16025 43092 16037 43095
rect 15896 43064 16037 43092
rect 15896 43052 15902 43064
rect 16025 43061 16037 43064
rect 16071 43061 16083 43095
rect 16025 43055 16083 43061
rect 16850 43052 16856 43104
rect 16908 43052 16914 43104
rect 17313 43095 17371 43101
rect 17313 43061 17325 43095
rect 17359 43092 17371 43095
rect 17494 43092 17500 43104
rect 17359 43064 17500 43092
rect 17359 43061 17371 43064
rect 17313 43055 17371 43061
rect 17494 43052 17500 43064
rect 17552 43052 17558 43104
rect 17586 43052 17592 43104
rect 17644 43052 17650 43104
rect 17678 43052 17684 43104
rect 17736 43052 17742 43104
rect 18138 43052 18144 43104
rect 18196 43052 18202 43104
rect 18414 43052 18420 43104
rect 18472 43052 18478 43104
rect 18506 43052 18512 43104
rect 18564 43092 18570 43104
rect 18693 43095 18751 43101
rect 18693 43092 18705 43095
rect 18564 43064 18705 43092
rect 18564 43052 18570 43064
rect 18693 43061 18705 43064
rect 18739 43061 18751 43095
rect 18693 43055 18751 43061
rect 19518 43052 19524 43104
rect 19576 43052 19582 43104
rect 24118 43052 24124 43104
rect 24176 43052 24182 43104
rect 1104 43002 24840 43024
rect 1104 42950 3917 43002
rect 3969 42950 3981 43002
rect 4033 42950 4045 43002
rect 4097 42950 4109 43002
rect 4161 42950 4173 43002
rect 4225 42950 9851 43002
rect 9903 42950 9915 43002
rect 9967 42950 9979 43002
rect 10031 42950 10043 43002
rect 10095 42950 10107 43002
rect 10159 42950 15785 43002
rect 15837 42950 15849 43002
rect 15901 42950 15913 43002
rect 15965 42950 15977 43002
rect 16029 42950 16041 43002
rect 16093 42950 21719 43002
rect 21771 42950 21783 43002
rect 21835 42950 21847 43002
rect 21899 42950 21911 43002
rect 21963 42950 21975 43002
rect 22027 42950 24840 43002
rect 1104 42928 24840 42950
rect 2222 42848 2228 42900
rect 2280 42848 2286 42900
rect 3326 42848 3332 42900
rect 3384 42848 3390 42900
rect 3786 42848 3792 42900
rect 3844 42888 3850 42900
rect 4157 42891 4215 42897
rect 4157 42888 4169 42891
rect 3844 42860 4169 42888
rect 3844 42848 3850 42860
rect 4157 42857 4169 42860
rect 4203 42857 4215 42891
rect 4157 42851 4215 42857
rect 6086 42848 6092 42900
rect 6144 42848 6150 42900
rect 6822 42848 6828 42900
rect 6880 42848 6886 42900
rect 7374 42848 7380 42900
rect 7432 42848 7438 42900
rect 9490 42848 9496 42900
rect 9548 42848 9554 42900
rect 9674 42848 9680 42900
rect 9732 42888 9738 42900
rect 10321 42891 10379 42897
rect 10321 42888 10333 42891
rect 9732 42860 10333 42888
rect 9732 42848 9738 42860
rect 10321 42857 10333 42860
rect 10367 42857 10379 42891
rect 10321 42851 10379 42857
rect 10594 42848 10600 42900
rect 10652 42848 10658 42900
rect 16301 42891 16359 42897
rect 16301 42888 16313 42891
rect 10980 42860 16313 42888
rect 8386 42820 8392 42832
rect 2148 42792 8392 42820
rect 1394 42712 1400 42764
rect 1452 42752 1458 42764
rect 1765 42755 1823 42761
rect 1765 42752 1777 42755
rect 1452 42724 1777 42752
rect 1452 42712 1458 42724
rect 1765 42721 1777 42724
rect 1811 42721 1823 42755
rect 1765 42715 1823 42721
rect 2148 42693 2176 42792
rect 8386 42780 8392 42792
rect 8444 42780 8450 42832
rect 8941 42823 8999 42829
rect 8941 42789 8953 42823
rect 8987 42820 8999 42823
rect 9508 42820 9536 42848
rect 10980 42820 11008 42860
rect 16301 42857 16313 42860
rect 16347 42857 16359 42891
rect 16301 42851 16359 42857
rect 16850 42848 16856 42900
rect 16908 42848 16914 42900
rect 17678 42848 17684 42900
rect 17736 42848 17742 42900
rect 18138 42888 18144 42900
rect 17880 42860 18144 42888
rect 8987 42792 9260 42820
rect 9508 42792 11008 42820
rect 8987 42789 8999 42792
rect 8941 42783 8999 42789
rect 2774 42712 2780 42764
rect 2832 42752 2838 42764
rect 2961 42755 3019 42761
rect 2961 42752 2973 42755
rect 2832 42724 2973 42752
rect 2832 42712 2838 42724
rect 2961 42721 2973 42724
rect 3007 42721 3019 42755
rect 2961 42715 3019 42721
rect 4890 42712 4896 42764
rect 4948 42752 4954 42764
rect 5353 42755 5411 42761
rect 5353 42752 5365 42755
rect 4948 42724 5365 42752
rect 4948 42712 4954 42724
rect 5353 42721 5365 42724
rect 5399 42721 5411 42755
rect 5353 42715 5411 42721
rect 8665 42755 8723 42761
rect 8665 42721 8677 42755
rect 8711 42752 8723 42755
rect 8754 42752 8760 42764
rect 8711 42724 8760 42752
rect 8711 42721 8723 42724
rect 8665 42715 8723 42721
rect 8754 42712 8760 42724
rect 8812 42712 8818 42764
rect 2133 42687 2191 42693
rect 2133 42653 2145 42687
rect 2179 42653 2191 42687
rect 2133 42647 2191 42653
rect 4246 42644 4252 42696
rect 4304 42684 4310 42696
rect 4525 42687 4583 42693
rect 4525 42684 4537 42687
rect 4304 42656 4537 42684
rect 4304 42644 4310 42656
rect 4525 42653 4537 42656
rect 4571 42653 4583 42687
rect 4525 42647 4583 42653
rect 4706 42644 4712 42696
rect 4764 42684 4770 42696
rect 5077 42687 5135 42693
rect 5077 42684 5089 42687
rect 4764 42656 5089 42684
rect 4764 42644 4770 42656
rect 5077 42653 5089 42656
rect 5123 42653 5135 42687
rect 5077 42647 5135 42653
rect 5537 42687 5595 42693
rect 5537 42653 5549 42687
rect 5583 42653 5595 42687
rect 5537 42647 5595 42653
rect 1489 42619 1547 42625
rect 1489 42585 1501 42619
rect 1535 42616 1547 42619
rect 2590 42616 2596 42628
rect 1535 42588 2596 42616
rect 1535 42585 1547 42588
rect 1489 42579 1547 42585
rect 2590 42576 2596 42588
rect 2648 42576 2654 42628
rect 2685 42619 2743 42625
rect 2685 42585 2697 42619
rect 2731 42616 2743 42619
rect 2731 42588 3096 42616
rect 2731 42585 2743 42588
rect 2685 42579 2743 42585
rect 3068 42560 3096 42588
rect 3234 42576 3240 42628
rect 3292 42576 3298 42628
rect 3878 42576 3884 42628
rect 3936 42616 3942 42628
rect 4065 42619 4123 42625
rect 4065 42616 4077 42619
rect 3936 42588 4077 42616
rect 3936 42576 3942 42588
rect 4065 42585 4077 42588
rect 4111 42585 4123 42619
rect 4065 42579 4123 42585
rect 3050 42508 3056 42560
rect 3108 42508 3114 42560
rect 3142 42508 3148 42560
rect 3200 42548 3206 42560
rect 4154 42548 4160 42560
rect 3200 42520 4160 42548
rect 3200 42508 3206 42520
rect 4154 42508 4160 42520
rect 4212 42508 4218 42560
rect 4614 42508 4620 42560
rect 4672 42548 4678 42560
rect 4709 42551 4767 42557
rect 4709 42548 4721 42551
rect 4672 42520 4721 42548
rect 4672 42508 4678 42520
rect 4709 42517 4721 42520
rect 4755 42517 4767 42551
rect 4709 42511 4767 42517
rect 4798 42508 4804 42560
rect 4856 42548 4862 42560
rect 5552 42548 5580 42647
rect 7742 42644 7748 42696
rect 7800 42644 7806 42696
rect 9122 42644 9128 42696
rect 9180 42644 9186 42696
rect 9232 42684 9260 42792
rect 11146 42780 11152 42832
rect 11204 42820 11210 42832
rect 16868 42820 16896 42848
rect 11204 42792 16896 42820
rect 11204 42780 11210 42792
rect 9306 42712 9312 42764
rect 9364 42752 9370 42764
rect 9769 42755 9827 42761
rect 9769 42752 9781 42755
rect 9364 42724 9781 42752
rect 9364 42712 9370 42724
rect 9769 42721 9781 42724
rect 9815 42721 9827 42755
rect 9769 42715 9827 42721
rect 12250 42712 12256 42764
rect 12308 42752 12314 42764
rect 12308 42724 13216 42752
rect 12308 42712 12314 42724
rect 9493 42687 9551 42693
rect 9493 42684 9505 42687
rect 9232 42656 9505 42684
rect 9493 42653 9505 42656
rect 9539 42653 9551 42687
rect 9493 42647 9551 42653
rect 9582 42644 9588 42696
rect 9640 42684 9646 42696
rect 10045 42687 10103 42693
rect 10045 42684 10057 42687
rect 9640 42656 10057 42684
rect 9640 42644 9646 42656
rect 10045 42653 10057 42656
rect 10091 42653 10103 42687
rect 10045 42647 10103 42653
rect 10505 42687 10563 42693
rect 10505 42653 10517 42687
rect 10551 42653 10563 42687
rect 10505 42647 10563 42653
rect 5994 42576 6000 42628
rect 6052 42576 6058 42628
rect 6730 42576 6736 42628
rect 6788 42576 6794 42628
rect 7282 42576 7288 42628
rect 7340 42576 7346 42628
rect 8389 42619 8447 42625
rect 7392 42588 8294 42616
rect 4856 42520 5580 42548
rect 4856 42508 4862 42520
rect 5718 42508 5724 42560
rect 5776 42508 5782 42560
rect 5902 42508 5908 42560
rect 5960 42548 5966 42560
rect 7392 42548 7420 42588
rect 5960 42520 7420 42548
rect 5960 42508 5966 42520
rect 7466 42508 7472 42560
rect 7524 42548 7530 42560
rect 7929 42551 7987 42557
rect 7929 42548 7941 42551
rect 7524 42520 7941 42548
rect 7524 42508 7530 42520
rect 7929 42517 7941 42520
rect 7975 42517 7987 42551
rect 8266 42548 8294 42588
rect 8389 42585 8401 42619
rect 8435 42616 8447 42619
rect 8754 42616 8760 42628
rect 8435 42588 8760 42616
rect 8435 42585 8447 42588
rect 8389 42579 8447 42585
rect 8754 42576 8760 42588
rect 8812 42576 8818 42628
rect 10520 42616 10548 42647
rect 10778 42644 10784 42696
rect 10836 42644 10842 42696
rect 11606 42644 11612 42696
rect 11664 42644 11670 42696
rect 11882 42644 11888 42696
rect 11940 42644 11946 42696
rect 12713 42687 12771 42693
rect 12713 42653 12725 42687
rect 12759 42653 12771 42687
rect 12713 42647 12771 42653
rect 12728 42616 12756 42647
rect 12986 42644 12992 42696
rect 13044 42644 13050 42696
rect 13078 42616 13084 42628
rect 9600 42588 10548 42616
rect 10612 42588 12434 42616
rect 12728 42588 13084 42616
rect 8662 42548 8668 42560
rect 8266 42520 8668 42548
rect 7929 42511 7987 42517
rect 8662 42508 8668 42520
rect 8720 42508 8726 42560
rect 9306 42508 9312 42560
rect 9364 42548 9370 42560
rect 9600 42548 9628 42588
rect 9364 42520 9628 42548
rect 9364 42508 9370 42520
rect 9766 42508 9772 42560
rect 9824 42548 9830 42560
rect 10229 42551 10287 42557
rect 10229 42548 10241 42551
rect 9824 42520 10241 42548
rect 9824 42508 9830 42520
rect 10229 42517 10241 42520
rect 10275 42517 10287 42551
rect 10229 42511 10287 42517
rect 10318 42508 10324 42560
rect 10376 42548 10382 42560
rect 10612 42548 10640 42588
rect 10376 42520 10640 42548
rect 10376 42508 10382 42520
rect 11790 42508 11796 42560
rect 11848 42508 11854 42560
rect 12066 42508 12072 42560
rect 12124 42508 12130 42560
rect 12406 42548 12434 42588
rect 13078 42576 13084 42588
rect 13136 42576 13142 42628
rect 13188 42557 13216 42724
rect 13814 42712 13820 42764
rect 13872 42752 13878 42764
rect 13872 42724 14688 42752
rect 13872 42712 13878 42724
rect 14090 42644 14096 42696
rect 14148 42644 14154 42696
rect 14366 42644 14372 42696
rect 14424 42644 14430 42696
rect 14660 42693 14688 42724
rect 15194 42712 15200 42764
rect 15252 42752 15258 42764
rect 17696 42752 17724 42848
rect 15252 42724 15608 42752
rect 15252 42712 15258 42724
rect 15580 42693 15608 42724
rect 17420 42724 17724 42752
rect 14645 42687 14703 42693
rect 14645 42653 14657 42687
rect 14691 42653 14703 42687
rect 14645 42647 14703 42653
rect 15289 42687 15347 42693
rect 15289 42653 15301 42687
rect 15335 42653 15347 42687
rect 15289 42647 15347 42653
rect 15565 42687 15623 42693
rect 15565 42653 15577 42687
rect 15611 42653 15623 42687
rect 15565 42647 15623 42653
rect 14918 42616 14924 42628
rect 14292 42588 14924 42616
rect 14292 42557 14320 42588
rect 14918 42576 14924 42588
rect 14976 42576 14982 42628
rect 15304 42616 15332 42647
rect 16482 42644 16488 42696
rect 16540 42644 16546 42696
rect 16574 42644 16580 42696
rect 16632 42644 16638 42696
rect 17420 42693 17448 42724
rect 17129 42687 17187 42693
rect 17129 42653 17141 42687
rect 17175 42653 17187 42687
rect 17129 42647 17187 42653
rect 17405 42687 17463 42693
rect 17405 42653 17417 42687
rect 17451 42653 17463 42687
rect 17405 42647 17463 42653
rect 16114 42616 16120 42628
rect 15304 42588 16120 42616
rect 16114 42576 16120 42588
rect 16172 42576 16178 42628
rect 17144 42616 17172 42647
rect 17586 42644 17592 42696
rect 17644 42644 17650 42696
rect 17681 42687 17739 42693
rect 17681 42653 17693 42687
rect 17727 42684 17739 42687
rect 17880 42684 17908 42860
rect 18138 42848 18144 42860
rect 18196 42848 18202 42900
rect 18874 42848 18880 42900
rect 18932 42848 18938 42900
rect 18966 42848 18972 42900
rect 19024 42888 19030 42900
rect 20806 42888 20812 42900
rect 19024 42860 20812 42888
rect 19024 42848 19030 42860
rect 20806 42848 20812 42860
rect 20864 42848 20870 42900
rect 18046 42780 18052 42832
rect 18104 42780 18110 42832
rect 18414 42752 18420 42764
rect 17972 42724 18420 42752
rect 17972 42693 18000 42724
rect 18414 42712 18420 42724
rect 18472 42712 18478 42764
rect 18524 42724 19196 42752
rect 17727 42656 17908 42684
rect 17957 42687 18015 42693
rect 17727 42653 17739 42656
rect 17681 42647 17739 42653
rect 17957 42653 17969 42687
rect 18003 42653 18015 42687
rect 17957 42647 18015 42653
rect 18233 42687 18291 42693
rect 18233 42653 18245 42687
rect 18279 42684 18291 42687
rect 18322 42684 18328 42696
rect 18279 42656 18328 42684
rect 18279 42653 18291 42656
rect 18233 42647 18291 42653
rect 18322 42644 18328 42656
rect 18380 42644 18386 42696
rect 18524 42693 18552 42724
rect 18509 42687 18567 42693
rect 18509 42653 18521 42687
rect 18555 42653 18567 42687
rect 18509 42647 18567 42653
rect 18785 42687 18843 42693
rect 18785 42653 18797 42687
rect 18831 42684 18843 42687
rect 18966 42684 18972 42696
rect 18831 42656 18972 42684
rect 18831 42653 18843 42656
rect 18785 42647 18843 42653
rect 18966 42644 18972 42656
rect 19024 42644 19030 42696
rect 19061 42687 19119 42693
rect 19061 42653 19073 42687
rect 19107 42653 19119 42687
rect 19061 42647 19119 42653
rect 17604 42616 17632 42644
rect 17144 42588 17632 42616
rect 18248 42588 18736 42616
rect 18248 42560 18276 42588
rect 12897 42551 12955 42557
rect 12897 42548 12909 42551
rect 12406 42520 12909 42548
rect 12897 42517 12909 42520
rect 12943 42517 12955 42551
rect 12897 42511 12955 42517
rect 13173 42551 13231 42557
rect 13173 42517 13185 42551
rect 13219 42517 13231 42551
rect 13173 42511 13231 42517
rect 14277 42551 14335 42557
rect 14277 42517 14289 42551
rect 14323 42517 14335 42551
rect 14277 42511 14335 42517
rect 14550 42508 14556 42560
rect 14608 42508 14614 42560
rect 14826 42508 14832 42560
rect 14884 42508 14890 42560
rect 15470 42508 15476 42560
rect 15528 42508 15534 42560
rect 15562 42508 15568 42560
rect 15620 42548 15626 42560
rect 15749 42551 15807 42557
rect 15749 42548 15761 42551
rect 15620 42520 15761 42548
rect 15620 42508 15626 42520
rect 15749 42517 15761 42520
rect 15795 42517 15807 42551
rect 15749 42511 15807 42517
rect 16390 42508 16396 42560
rect 16448 42548 16454 42560
rect 16761 42551 16819 42557
rect 16761 42548 16773 42551
rect 16448 42520 16773 42548
rect 16448 42508 16454 42520
rect 16761 42517 16773 42520
rect 16807 42517 16819 42551
rect 16761 42511 16819 42517
rect 16942 42508 16948 42560
rect 17000 42508 17006 42560
rect 17218 42508 17224 42560
rect 17276 42508 17282 42560
rect 17310 42508 17316 42560
rect 17368 42548 17374 42560
rect 17497 42551 17555 42557
rect 17497 42548 17509 42551
rect 17368 42520 17509 42548
rect 17368 42508 17374 42520
rect 17497 42517 17509 42520
rect 17543 42517 17555 42551
rect 17497 42511 17555 42517
rect 17770 42508 17776 42560
rect 17828 42508 17834 42560
rect 18230 42508 18236 42560
rect 18288 42508 18294 42560
rect 18322 42508 18328 42560
rect 18380 42508 18386 42560
rect 18598 42508 18604 42560
rect 18656 42508 18662 42560
rect 18708 42548 18736 42588
rect 19076 42548 19104 42647
rect 19168 42616 19196 42724
rect 21358 42712 21364 42764
rect 21416 42752 21422 42764
rect 23477 42755 23535 42761
rect 21416 42724 23244 42752
rect 21416 42712 21422 42724
rect 19242 42644 19248 42696
rect 19300 42644 19306 42696
rect 21266 42644 21272 42696
rect 21324 42644 21330 42696
rect 21910 42644 21916 42696
rect 21968 42644 21974 42696
rect 22370 42644 22376 42696
rect 22428 42684 22434 42696
rect 23216 42693 23244 42724
rect 23477 42721 23489 42755
rect 23523 42752 23535 42755
rect 25130 42752 25136 42764
rect 23523 42724 25136 42752
rect 23523 42721 23535 42724
rect 23477 42715 23535 42721
rect 25130 42712 25136 42724
rect 25188 42712 25194 42764
rect 22649 42687 22707 42693
rect 22649 42684 22661 42687
rect 22428 42656 22661 42684
rect 22428 42644 22434 42656
rect 22649 42653 22661 42656
rect 22695 42653 22707 42687
rect 22649 42647 22707 42653
rect 23201 42687 23259 42693
rect 23201 42653 23213 42687
rect 23247 42653 23259 42687
rect 23201 42647 23259 42653
rect 24121 42687 24179 42693
rect 24121 42653 24133 42687
rect 24167 42684 24179 42687
rect 24210 42684 24216 42696
rect 24167 42656 24216 42684
rect 24167 42653 24179 42656
rect 24121 42647 24179 42653
rect 24210 42644 24216 42656
rect 24268 42644 24274 42696
rect 24578 42644 24584 42696
rect 24636 42644 24642 42696
rect 19168 42588 21128 42616
rect 18708 42520 19104 42548
rect 20530 42508 20536 42560
rect 20588 42508 20594 42560
rect 21100 42557 21128 42588
rect 21542 42576 21548 42628
rect 21600 42576 21606 42628
rect 22097 42619 22155 42625
rect 22097 42585 22109 42619
rect 22143 42585 22155 42619
rect 22097 42579 22155 42585
rect 22465 42619 22523 42625
rect 22465 42585 22477 42619
rect 22511 42616 22523 42619
rect 22511 42588 23520 42616
rect 22511 42585 22523 42588
rect 22465 42579 22523 42585
rect 21085 42551 21143 42557
rect 21085 42517 21097 42551
rect 21131 42517 21143 42551
rect 21085 42511 21143 42517
rect 21174 42508 21180 42560
rect 21232 42548 21238 42560
rect 22112 42548 22140 42579
rect 21232 42520 22140 42548
rect 21232 42508 21238 42520
rect 22278 42508 22284 42560
rect 22336 42548 22342 42560
rect 22741 42551 22799 42557
rect 22741 42548 22753 42551
rect 22336 42520 22753 42548
rect 22336 42508 22342 42520
rect 22741 42517 22753 42520
rect 22787 42517 22799 42551
rect 23492 42548 23520 42588
rect 23750 42576 23756 42628
rect 23808 42576 23814 42628
rect 24596 42548 24624 42644
rect 23492 42520 24624 42548
rect 22741 42511 22799 42517
rect 1104 42458 25000 42480
rect 1104 42406 6884 42458
rect 6936 42406 6948 42458
rect 7000 42406 7012 42458
rect 7064 42406 7076 42458
rect 7128 42406 7140 42458
rect 7192 42406 12818 42458
rect 12870 42406 12882 42458
rect 12934 42406 12946 42458
rect 12998 42406 13010 42458
rect 13062 42406 13074 42458
rect 13126 42406 18752 42458
rect 18804 42406 18816 42458
rect 18868 42406 18880 42458
rect 18932 42406 18944 42458
rect 18996 42406 19008 42458
rect 19060 42406 24686 42458
rect 24738 42406 24750 42458
rect 24802 42406 24814 42458
rect 24866 42406 24878 42458
rect 24930 42406 24942 42458
rect 24994 42406 25000 42458
rect 1104 42384 25000 42406
rect 474 42304 480 42356
rect 532 42344 538 42356
rect 1581 42347 1639 42353
rect 1581 42344 1593 42347
rect 532 42316 1593 42344
rect 532 42304 538 42316
rect 1581 42313 1593 42316
rect 1627 42313 1639 42347
rect 2314 42344 2320 42356
rect 1581 42307 1639 42313
rect 1964 42316 2320 42344
rect 1489 42279 1547 42285
rect 1489 42245 1501 42279
rect 1535 42276 1547 42279
rect 1964 42276 1992 42316
rect 2314 42304 2320 42316
rect 2372 42304 2378 42356
rect 2501 42347 2559 42353
rect 2501 42313 2513 42347
rect 2547 42344 2559 42347
rect 3142 42344 3148 42356
rect 2547 42316 3148 42344
rect 2547 42313 2559 42316
rect 2501 42307 2559 42313
rect 3142 42304 3148 42316
rect 3200 42304 3206 42356
rect 3234 42304 3240 42356
rect 3292 42344 3298 42356
rect 3421 42347 3479 42353
rect 3421 42344 3433 42347
rect 3292 42316 3433 42344
rect 3292 42304 3298 42316
rect 3421 42313 3433 42316
rect 3467 42313 3479 42347
rect 3421 42307 3479 42313
rect 3697 42347 3755 42353
rect 3697 42313 3709 42347
rect 3743 42344 3755 42347
rect 3743 42316 4200 42344
rect 3743 42313 3755 42316
rect 3697 42307 3755 42313
rect 1535 42248 1992 42276
rect 1535 42245 1547 42248
rect 1489 42239 1547 42245
rect 2038 42236 2044 42288
rect 2096 42236 2102 42288
rect 4172 42276 4200 42316
rect 4890 42304 4896 42356
rect 4948 42344 4954 42356
rect 4985 42347 5043 42353
rect 4985 42344 4997 42347
rect 4948 42316 4997 42344
rect 4948 42304 4954 42316
rect 4985 42313 4997 42316
rect 5031 42313 5043 42347
rect 4985 42307 5043 42313
rect 5169 42347 5227 42353
rect 5169 42313 5181 42347
rect 5215 42313 5227 42347
rect 5902 42344 5908 42356
rect 5169 42307 5227 42313
rect 5368 42316 5908 42344
rect 4172 42248 4844 42276
rect 3712 42220 3924 42232
rect 2130 42168 2136 42220
rect 2188 42208 2194 42220
rect 2685 42211 2743 42217
rect 2685 42208 2697 42211
rect 2188 42180 2697 42208
rect 2188 42168 2194 42180
rect 2685 42177 2697 42180
rect 2731 42177 2743 42211
rect 2685 42171 2743 42177
rect 2774 42168 2780 42220
rect 2832 42168 2838 42220
rect 3326 42168 3332 42220
rect 3384 42208 3390 42220
rect 3605 42211 3663 42217
rect 3605 42208 3617 42211
rect 3384 42180 3617 42208
rect 3384 42168 3390 42180
rect 3605 42177 3617 42180
rect 3651 42177 3663 42211
rect 3605 42171 3663 42177
rect 3694 42168 3700 42220
rect 3752 42217 3924 42220
rect 3752 42211 3939 42217
rect 3752 42204 3893 42211
rect 3752 42168 3758 42204
rect 3881 42177 3893 42204
rect 3927 42177 3939 42211
rect 3881 42171 3939 42177
rect 3970 42168 3976 42220
rect 4028 42168 4034 42220
rect 4062 42168 4068 42220
rect 4120 42208 4126 42220
rect 4120 42180 4200 42208
rect 4120 42168 4126 42180
rect 3510 42140 3516 42152
rect 2976 42112 3516 42140
rect 2976 42081 3004 42112
rect 3510 42100 3516 42112
rect 3568 42100 3574 42152
rect 4172 42081 4200 42180
rect 4706 42168 4712 42220
rect 4764 42168 4770 42220
rect 4816 42217 4844 42248
rect 5184 42220 5212 42307
rect 4801 42211 4859 42217
rect 4801 42177 4813 42211
rect 4847 42177 4859 42211
rect 4801 42171 4859 42177
rect 5166 42168 5172 42220
rect 5224 42168 5230 42220
rect 5368 42217 5396 42316
rect 5902 42304 5908 42316
rect 5960 42304 5966 42356
rect 5997 42347 6055 42353
rect 5997 42313 6009 42347
rect 6043 42344 6055 42347
rect 6270 42344 6276 42356
rect 6043 42316 6276 42344
rect 6043 42313 6055 42316
rect 5997 42307 6055 42313
rect 6270 42304 6276 42316
rect 6328 42304 6334 42356
rect 7190 42304 7196 42356
rect 7248 42344 7254 42356
rect 7374 42344 7380 42356
rect 7248 42316 7380 42344
rect 7248 42304 7254 42316
rect 7374 42304 7380 42316
rect 7432 42304 7438 42356
rect 8202 42304 8208 42356
rect 8260 42344 8266 42356
rect 8481 42347 8539 42353
rect 8481 42344 8493 42347
rect 8260 42316 8493 42344
rect 8260 42304 8266 42316
rect 8481 42313 8493 42316
rect 8527 42313 8539 42347
rect 9953 42347 10011 42353
rect 9953 42344 9965 42347
rect 8481 42307 8539 42313
rect 9692 42316 9965 42344
rect 5442 42236 5448 42288
rect 5500 42236 5506 42288
rect 5810 42236 5816 42288
rect 5868 42276 5874 42288
rect 5868 42248 8524 42276
rect 5868 42236 5874 42248
rect 5353 42211 5411 42217
rect 5353 42177 5365 42211
rect 5399 42177 5411 42211
rect 5353 42171 5411 42177
rect 4982 42100 4988 42152
rect 5040 42140 5046 42152
rect 5460 42140 5488 42236
rect 5721 42211 5779 42217
rect 5721 42177 5733 42211
rect 5767 42208 5779 42211
rect 6181 42211 6239 42217
rect 6181 42208 6193 42211
rect 5767 42180 6193 42208
rect 5767 42177 5779 42180
rect 5721 42171 5779 42177
rect 6181 42177 6193 42180
rect 6227 42208 6239 42211
rect 6549 42211 6607 42217
rect 6227 42180 6316 42208
rect 6227 42177 6239 42180
rect 6181 42171 6239 42177
rect 6288 42152 6316 42180
rect 6549 42177 6561 42211
rect 6595 42177 6607 42211
rect 6549 42171 6607 42177
rect 6825 42211 6883 42217
rect 6825 42177 6837 42211
rect 6871 42208 6883 42211
rect 6871 42180 7236 42208
rect 6871 42177 6883 42180
rect 6825 42171 6883 42177
rect 5040 42112 5488 42140
rect 5040 42100 5046 42112
rect 6270 42100 6276 42152
rect 6328 42100 6334 42152
rect 6564 42140 6592 42171
rect 6914 42140 6920 42152
rect 6564 42112 6920 42140
rect 6914 42100 6920 42112
rect 6972 42100 6978 42152
rect 7208 42149 7236 42180
rect 7466 42168 7472 42220
rect 7524 42168 7530 42220
rect 7650 42168 7656 42220
rect 7708 42208 7714 42220
rect 7929 42211 7987 42217
rect 7929 42208 7941 42211
rect 7708 42180 7941 42208
rect 7708 42168 7714 42180
rect 7929 42177 7941 42180
rect 7975 42177 7987 42211
rect 7929 42171 7987 42177
rect 8202 42168 8208 42220
rect 8260 42168 8266 42220
rect 8389 42211 8447 42217
rect 8389 42177 8401 42211
rect 8435 42177 8447 42211
rect 8496 42208 8524 42248
rect 8570 42236 8576 42288
rect 8628 42276 8634 42288
rect 9122 42276 9128 42288
rect 8628 42248 9128 42276
rect 8628 42236 8634 42248
rect 9122 42236 9128 42248
rect 9180 42236 9186 42288
rect 8846 42208 8852 42220
rect 8496 42180 8852 42208
rect 8389 42171 8447 42177
rect 7193 42143 7251 42149
rect 7193 42109 7205 42143
rect 7239 42140 7251 42143
rect 7239 42112 7788 42140
rect 7239 42109 7251 42112
rect 7193 42103 7251 42109
rect 2961 42075 3019 42081
rect 2961 42041 2973 42075
rect 3007 42041 3019 42075
rect 2961 42035 3019 42041
rect 4157 42075 4215 42081
rect 4157 42041 4169 42075
rect 4203 42041 4215 42075
rect 4157 42035 4215 42041
rect 5810 42032 5816 42084
rect 5868 42072 5874 42084
rect 6365 42075 6423 42081
rect 6365 42072 6377 42075
rect 5868 42044 6377 42072
rect 5868 42032 5874 42044
rect 6365 42041 6377 42044
rect 6411 42041 6423 42075
rect 6365 42035 6423 42041
rect 6641 42075 6699 42081
rect 6641 42041 6653 42075
rect 6687 42072 6699 42075
rect 7558 42072 7564 42084
rect 6687 42044 7564 42072
rect 6687 42041 6699 42044
rect 6641 42035 6699 42041
rect 7558 42032 7564 42044
rect 7616 42032 7622 42084
rect 7760 42072 7788 42112
rect 7834 42100 7840 42152
rect 7892 42140 7898 42152
rect 8404 42140 8432 42171
rect 8846 42168 8852 42180
rect 8904 42168 8910 42220
rect 9030 42168 9036 42220
rect 9088 42168 9094 42220
rect 9401 42211 9459 42217
rect 9401 42177 9413 42211
rect 9447 42208 9459 42211
rect 9490 42208 9496 42220
rect 9447 42180 9496 42208
rect 9447 42177 9459 42180
rect 9401 42171 9459 42177
rect 9490 42168 9496 42180
rect 9548 42168 9554 42220
rect 9692 42208 9720 42316
rect 9953 42313 9965 42316
rect 9999 42313 10011 42347
rect 17218 42344 17224 42356
rect 9953 42307 10011 42313
rect 16776 42316 17224 42344
rect 9766 42236 9772 42288
rect 9824 42276 9830 42288
rect 9824 42248 9904 42276
rect 9824 42236 9830 42248
rect 9876 42217 9904 42248
rect 14734 42236 14740 42288
rect 14792 42276 14798 42288
rect 16390 42276 16396 42288
rect 14792 42248 16396 42276
rect 14792 42236 14798 42248
rect 16390 42236 16396 42248
rect 16448 42236 16454 42288
rect 16776 42285 16804 42316
rect 17218 42304 17224 42316
rect 17276 42304 17282 42356
rect 17310 42304 17316 42356
rect 17368 42304 17374 42356
rect 17770 42304 17776 42356
rect 17828 42304 17834 42356
rect 18322 42304 18328 42356
rect 18380 42304 18386 42356
rect 19705 42347 19763 42353
rect 18432 42316 19012 42344
rect 16761 42279 16819 42285
rect 16761 42245 16773 42279
rect 16807 42245 16819 42279
rect 16761 42239 16819 42245
rect 16942 42236 16948 42288
rect 17000 42236 17006 42288
rect 17129 42279 17187 42285
rect 17129 42245 17141 42279
rect 17175 42276 17187 42279
rect 17328 42276 17356 42304
rect 17175 42248 17356 42276
rect 17497 42279 17555 42285
rect 17175 42245 17187 42248
rect 17129 42239 17187 42245
rect 17497 42245 17509 42279
rect 17543 42276 17555 42279
rect 17788 42276 17816 42304
rect 17543 42248 17816 42276
rect 17865 42279 17923 42285
rect 17543 42245 17555 42248
rect 17497 42239 17555 42245
rect 17865 42245 17877 42279
rect 17911 42276 17923 42279
rect 18046 42276 18052 42288
rect 17911 42248 18052 42276
rect 17911 42245 17923 42248
rect 17865 42239 17923 42245
rect 18046 42236 18052 42248
rect 18104 42236 18110 42288
rect 18233 42279 18291 42285
rect 18233 42245 18245 42279
rect 18279 42276 18291 42279
rect 18340 42276 18368 42304
rect 18432 42288 18460 42316
rect 18279 42248 18368 42276
rect 18279 42245 18291 42248
rect 18233 42239 18291 42245
rect 18414 42236 18420 42288
rect 18472 42236 18478 42288
rect 18598 42236 18604 42288
rect 18656 42236 18662 42288
rect 18984 42285 19012 42316
rect 19705 42313 19717 42347
rect 19751 42313 19763 42347
rect 19705 42307 19763 42313
rect 19981 42347 20039 42353
rect 19981 42313 19993 42347
rect 20027 42344 20039 42347
rect 20533 42347 20591 42353
rect 20027 42316 20484 42344
rect 20027 42313 20039 42316
rect 19981 42307 20039 42313
rect 18969 42279 19027 42285
rect 18969 42245 18981 42279
rect 19015 42245 19027 42279
rect 18969 42239 19027 42245
rect 19337 42279 19395 42285
rect 19337 42245 19349 42279
rect 19383 42276 19395 42279
rect 19518 42276 19524 42288
rect 19383 42248 19524 42276
rect 19383 42245 19395 42248
rect 19337 42239 19395 42245
rect 19518 42236 19524 42248
rect 19576 42236 19582 42288
rect 19720 42276 19748 42307
rect 19720 42248 20208 42276
rect 9600 42180 9720 42208
rect 9861 42211 9919 42217
rect 7892 42112 8432 42140
rect 7892 42100 7898 42112
rect 8754 42100 8760 42152
rect 8812 42140 8818 42152
rect 9600 42140 9628 42180
rect 9861 42177 9873 42211
rect 9907 42177 9919 42211
rect 9861 42171 9919 42177
rect 10137 42211 10195 42217
rect 10137 42177 10149 42211
rect 10183 42177 10195 42211
rect 10137 42171 10195 42177
rect 16117 42211 16175 42217
rect 16117 42177 16129 42211
rect 16163 42208 16175 42211
rect 16960 42208 16988 42236
rect 16163 42180 16988 42208
rect 16163 42177 16175 42180
rect 16117 42171 16175 42177
rect 10152 42140 10180 42171
rect 17034 42168 17040 42220
rect 17092 42208 17098 42220
rect 20180 42217 20208 42248
rect 20456 42217 20484 42316
rect 20533 42313 20545 42347
rect 20579 42344 20591 42347
rect 20622 42344 20628 42356
rect 20579 42316 20628 42344
rect 20579 42313 20591 42316
rect 20533 42307 20591 42313
rect 20622 42304 20628 42316
rect 20680 42304 20686 42356
rect 20806 42304 20812 42356
rect 20864 42304 20870 42356
rect 21634 42304 21640 42356
rect 21692 42344 21698 42356
rect 21821 42347 21879 42353
rect 21821 42344 21833 42347
rect 21692 42316 21833 42344
rect 21692 42304 21698 42316
rect 21821 42313 21833 42316
rect 21867 42313 21879 42347
rect 21821 42307 21879 42313
rect 22557 42347 22615 42353
rect 22557 42313 22569 42347
rect 22603 42344 22615 42347
rect 23109 42347 23167 42353
rect 22603 42316 23060 42344
rect 22603 42313 22615 42316
rect 22557 42307 22615 42313
rect 22738 42276 22744 42288
rect 21652 42248 22744 42276
rect 19889 42211 19947 42217
rect 19889 42208 19901 42211
rect 17092 42180 19901 42208
rect 17092 42168 17098 42180
rect 19889 42177 19901 42180
rect 19935 42177 19947 42211
rect 19889 42171 19947 42177
rect 20165 42211 20223 42217
rect 20165 42177 20177 42211
rect 20211 42177 20223 42211
rect 20165 42171 20223 42177
rect 20441 42211 20499 42217
rect 20441 42177 20453 42211
rect 20487 42177 20499 42211
rect 20441 42171 20499 42177
rect 20717 42211 20775 42217
rect 20717 42177 20729 42211
rect 20763 42177 20775 42211
rect 20717 42171 20775 42177
rect 8812 42112 9628 42140
rect 9884 42112 10180 42140
rect 8812 42100 8818 42112
rect 9677 42075 9735 42081
rect 7760 42044 8984 42072
rect 1302 41964 1308 42016
rect 1360 42004 1366 42016
rect 2133 42007 2191 42013
rect 2133 42004 2145 42007
rect 1360 41976 2145 42004
rect 1360 41964 1366 41976
rect 2133 41973 2145 41976
rect 2179 41973 2191 42007
rect 2133 41967 2191 41973
rect 3326 41964 3332 42016
rect 3384 42004 3390 42016
rect 4430 42004 4436 42016
rect 3384 41976 4436 42004
rect 3384 41964 3390 41976
rect 4430 41964 4436 41976
rect 4488 41964 4494 42016
rect 4522 41964 4528 42016
rect 4580 41964 4586 42016
rect 4890 41964 4896 42016
rect 4948 42004 4954 42016
rect 7098 42004 7104 42016
rect 4948 41976 7104 42004
rect 4948 41964 4954 41976
rect 7098 41964 7104 41976
rect 7156 41964 7162 42016
rect 7285 42007 7343 42013
rect 7285 41973 7297 42007
rect 7331 42004 7343 42007
rect 7374 42004 7380 42016
rect 7331 41976 7380 42004
rect 7331 41973 7343 41976
rect 7285 41967 7343 41973
rect 7374 41964 7380 41976
rect 7432 41964 7438 42016
rect 7745 42007 7803 42013
rect 7745 41973 7757 42007
rect 7791 42004 7803 42007
rect 7926 42004 7932 42016
rect 7791 41976 7932 42004
rect 7791 41973 7803 41976
rect 7745 41967 7803 41973
rect 7926 41964 7932 41976
rect 7984 41964 7990 42016
rect 8018 41964 8024 42016
rect 8076 41964 8082 42016
rect 8846 41964 8852 42016
rect 8904 41964 8910 42016
rect 8956 42004 8984 42044
rect 9677 42041 9689 42075
rect 9723 42072 9735 42075
rect 9884 42072 9912 42112
rect 11698 42100 11704 42152
rect 11756 42140 11762 42152
rect 11756 42112 18644 42140
rect 11756 42100 11762 42112
rect 9723 42044 9912 42072
rect 9723 42041 9735 42044
rect 9677 42035 9735 42041
rect 15378 42032 15384 42084
rect 15436 42072 15442 42084
rect 16482 42072 16488 42084
rect 15436 42044 16488 42072
rect 15436 42032 15442 42044
rect 16482 42032 16488 42044
rect 16540 42032 16546 42084
rect 16942 42032 16948 42084
rect 17000 42032 17006 42084
rect 17310 42032 17316 42084
rect 17368 42032 17374 42084
rect 17678 42032 17684 42084
rect 17736 42032 17742 42084
rect 18046 42032 18052 42084
rect 18104 42032 18110 42084
rect 18616 42072 18644 42112
rect 19168 42112 20208 42140
rect 19168 42081 19196 42112
rect 19153 42075 19211 42081
rect 18616 42044 18828 42072
rect 9766 42004 9772 42016
rect 8956 41976 9772 42004
rect 9766 41964 9772 41976
rect 9824 41964 9830 42016
rect 16298 41964 16304 42016
rect 16356 41964 16362 42016
rect 18322 41964 18328 42016
rect 18380 41964 18386 42016
rect 18506 41964 18512 42016
rect 18564 42004 18570 42016
rect 18693 42007 18751 42013
rect 18693 42004 18705 42007
rect 18564 41976 18705 42004
rect 18564 41964 18570 41976
rect 18693 41973 18705 41976
rect 18739 41973 18751 42007
rect 18800 42004 18828 42044
rect 19153 42041 19165 42075
rect 19199 42041 19211 42075
rect 19153 42035 19211 42041
rect 19518 42032 19524 42084
rect 19576 42032 19582 42084
rect 19886 42032 19892 42084
rect 19944 42032 19950 42084
rect 20180 42072 20208 42112
rect 20254 42100 20260 42152
rect 20312 42140 20318 42152
rect 20732 42140 20760 42171
rect 20990 42168 20996 42220
rect 21048 42168 21054 42220
rect 21266 42168 21272 42220
rect 21324 42168 21330 42220
rect 21652 42217 21680 42248
rect 22738 42236 22744 42248
rect 22796 42236 22802 42288
rect 23032 42276 23060 42316
rect 23109 42313 23121 42347
rect 23155 42344 23167 42347
rect 23198 42344 23204 42356
rect 23155 42316 23204 42344
rect 23155 42313 23167 42316
rect 23109 42307 23167 42313
rect 23198 42304 23204 42316
rect 23256 42304 23262 42356
rect 23661 42347 23719 42353
rect 23661 42313 23673 42347
rect 23707 42344 23719 42347
rect 24486 42344 24492 42356
rect 23707 42316 24492 42344
rect 23707 42313 23719 42316
rect 23661 42307 23719 42313
rect 24486 42304 24492 42316
rect 24544 42304 24550 42356
rect 25590 42304 25596 42356
rect 25648 42304 25654 42356
rect 25608 42276 25636 42304
rect 23032 42248 25636 42276
rect 21637 42211 21695 42217
rect 21637 42177 21649 42211
rect 21683 42177 21695 42211
rect 21637 42171 21695 42177
rect 22005 42211 22063 42217
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 22281 42211 22339 42217
rect 22281 42177 22293 42211
rect 22327 42177 22339 42211
rect 22281 42171 22339 42177
rect 20312 42112 20760 42140
rect 20312 42100 20318 42112
rect 20898 42100 20904 42152
rect 20956 42140 20962 42152
rect 22020 42140 22048 42171
rect 20956 42112 22048 42140
rect 20956 42100 20962 42112
rect 20990 42072 20996 42084
rect 20180 42044 20996 42072
rect 20990 42032 20996 42044
rect 21048 42032 21054 42084
rect 22296 42072 22324 42171
rect 22830 42168 22836 42220
rect 22888 42168 22894 42220
rect 23385 42211 23443 42217
rect 23385 42177 23397 42211
rect 23431 42208 23443 42211
rect 23431 42180 23980 42208
rect 23431 42177 23443 42180
rect 23385 42171 23443 42177
rect 22370 42100 22376 42152
rect 22428 42140 22434 42152
rect 23952 42140 23980 42180
rect 24026 42168 24032 42220
rect 24084 42168 24090 42220
rect 24578 42140 24584 42152
rect 22428 42112 23888 42140
rect 23952 42112 24584 42140
rect 22428 42100 22434 42112
rect 23566 42072 23572 42084
rect 22296 42044 23572 42072
rect 23566 42032 23572 42044
rect 23624 42032 23630 42084
rect 23860 42072 23888 42112
rect 24578 42100 24584 42112
rect 24636 42100 24642 42152
rect 24210 42072 24216 42084
rect 23860 42044 24216 42072
rect 24210 42032 24216 42044
rect 24268 42032 24274 42084
rect 19702 42004 19708 42016
rect 18800 41976 19708 42004
rect 18693 41967 18751 41973
rect 19702 41964 19708 41976
rect 19760 41964 19766 42016
rect 19904 42004 19932 42032
rect 20257 42007 20315 42013
rect 20257 42004 20269 42007
rect 19904 41976 20269 42004
rect 20257 41973 20269 41976
rect 20303 41973 20315 42007
rect 20257 41967 20315 41973
rect 22278 41964 22284 42016
rect 22336 42004 22342 42016
rect 23474 42004 23480 42016
rect 22336 41976 23480 42004
rect 22336 41964 22342 41976
rect 23474 41964 23480 41976
rect 23532 41964 23538 42016
rect 24305 42007 24363 42013
rect 24305 41973 24317 42007
rect 24351 42004 24363 42007
rect 25130 42004 25136 42016
rect 24351 41976 25136 42004
rect 24351 41973 24363 41976
rect 24305 41967 24363 41973
rect 25130 41964 25136 41976
rect 25188 41964 25194 42016
rect 1104 41914 24840 41936
rect 1104 41862 3917 41914
rect 3969 41862 3981 41914
rect 4033 41862 4045 41914
rect 4097 41862 4109 41914
rect 4161 41862 4173 41914
rect 4225 41862 9851 41914
rect 9903 41862 9915 41914
rect 9967 41862 9979 41914
rect 10031 41862 10043 41914
rect 10095 41862 10107 41914
rect 10159 41862 15785 41914
rect 15837 41862 15849 41914
rect 15901 41862 15913 41914
rect 15965 41862 15977 41914
rect 16029 41862 16041 41914
rect 16093 41862 21719 41914
rect 21771 41862 21783 41914
rect 21835 41862 21847 41914
rect 21899 41862 21911 41914
rect 21963 41862 21975 41914
rect 22027 41862 24840 41914
rect 1104 41840 24840 41862
rect 934 41760 940 41812
rect 992 41800 998 41812
rect 1581 41803 1639 41809
rect 1581 41800 1593 41803
rect 992 41772 1593 41800
rect 992 41760 998 41772
rect 1581 41769 1593 41772
rect 1627 41769 1639 41803
rect 1581 41763 1639 41769
rect 1670 41760 1676 41812
rect 1728 41800 1734 41812
rect 2133 41803 2191 41809
rect 2133 41800 2145 41803
rect 1728 41772 2145 41800
rect 1728 41760 1734 41772
rect 2133 41769 2145 41772
rect 2179 41769 2191 41803
rect 2133 41763 2191 41769
rect 2498 41760 2504 41812
rect 2556 41760 2562 41812
rect 2590 41760 2596 41812
rect 2648 41760 2654 41812
rect 2774 41760 2780 41812
rect 2832 41800 2838 41812
rect 3145 41803 3203 41809
rect 3145 41800 3157 41803
rect 2832 41772 3157 41800
rect 2832 41760 2838 41772
rect 3145 41769 3157 41772
rect 3191 41769 3203 41803
rect 3145 41763 3203 41769
rect 3418 41760 3424 41812
rect 3476 41760 3482 41812
rect 3878 41760 3884 41812
rect 3936 41760 3942 41812
rect 4065 41803 4123 41809
rect 4065 41769 4077 41803
rect 4111 41800 4123 41803
rect 4246 41800 4252 41812
rect 4111 41772 4252 41800
rect 4111 41769 4123 41772
rect 4065 41763 4123 41769
rect 4246 41760 4252 41772
rect 4304 41760 4310 41812
rect 4617 41803 4675 41809
rect 4617 41769 4629 41803
rect 4663 41800 4675 41803
rect 4982 41800 4988 41812
rect 4663 41772 4988 41800
rect 4663 41769 4675 41772
rect 4617 41763 4675 41769
rect 4982 41760 4988 41772
rect 5040 41760 5046 41812
rect 5534 41800 5540 41812
rect 5368 41772 5540 41800
rect 2608 41732 2636 41760
rect 3789 41735 3847 41741
rect 3789 41732 3801 41735
rect 2608 41704 3801 41732
rect 3789 41701 3801 41704
rect 3835 41701 3847 41735
rect 3896 41732 3924 41760
rect 4341 41735 4399 41741
rect 3896 41704 4292 41732
rect 3789 41695 3847 41701
rect 1118 41624 1124 41676
rect 1176 41664 1182 41676
rect 1176 41636 2728 41664
rect 1176 41624 1182 41636
rect 2700 41605 2728 41636
rect 2866 41624 2872 41676
rect 2924 41664 2930 41676
rect 4264 41664 4292 41704
rect 4341 41701 4353 41735
rect 4387 41732 4399 41735
rect 4798 41732 4804 41744
rect 4387 41704 4804 41732
rect 4387 41701 4399 41704
rect 4341 41695 4399 41701
rect 4798 41692 4804 41704
rect 4856 41692 4862 41744
rect 4893 41735 4951 41741
rect 4893 41701 4905 41735
rect 4939 41732 4951 41735
rect 5368 41732 5396 41772
rect 5534 41760 5540 41772
rect 5592 41760 5598 41812
rect 5721 41803 5779 41809
rect 5721 41769 5733 41803
rect 5767 41800 5779 41803
rect 5994 41800 6000 41812
rect 5767 41772 6000 41800
rect 5767 41769 5779 41772
rect 5721 41763 5779 41769
rect 5994 41760 6000 41772
rect 6052 41760 6058 41812
rect 6730 41800 6736 41812
rect 6104 41772 6736 41800
rect 4939 41704 5396 41732
rect 5445 41735 5503 41741
rect 4939 41701 4951 41704
rect 4893 41695 4951 41701
rect 5445 41701 5457 41735
rect 5491 41732 5503 41735
rect 6104 41732 6132 41772
rect 6730 41760 6736 41772
rect 6788 41760 6794 41812
rect 7193 41803 7251 41809
rect 7193 41769 7205 41803
rect 7239 41800 7251 41803
rect 7282 41800 7288 41812
rect 7239 41772 7288 41800
rect 7239 41769 7251 41772
rect 7193 41763 7251 41769
rect 7282 41760 7288 41772
rect 7340 41760 7346 41812
rect 7374 41760 7380 41812
rect 7432 41760 7438 41812
rect 7561 41803 7619 41809
rect 7561 41769 7573 41803
rect 7607 41800 7619 41803
rect 7742 41800 7748 41812
rect 7607 41772 7748 41800
rect 7607 41769 7619 41772
rect 7561 41763 7619 41769
rect 7742 41760 7748 41772
rect 7800 41760 7806 41812
rect 7926 41760 7932 41812
rect 7984 41760 7990 41812
rect 8110 41760 8116 41812
rect 8168 41760 8174 41812
rect 8386 41760 8392 41812
rect 8444 41760 8450 41812
rect 8846 41760 8852 41812
rect 8904 41760 8910 41812
rect 8938 41760 8944 41812
rect 8996 41760 9002 41812
rect 9030 41760 9036 41812
rect 9088 41800 9094 41812
rect 12526 41800 12532 41812
rect 9088 41772 12532 41800
rect 9088 41760 9094 41772
rect 12526 41760 12532 41772
rect 12584 41760 12590 41812
rect 17862 41760 17868 41812
rect 17920 41800 17926 41812
rect 17920 41772 18184 41800
rect 17920 41760 17926 41772
rect 5491 41704 6132 41732
rect 6549 41735 6607 41741
rect 5491 41701 5503 41704
rect 5445 41695 5503 41701
rect 6549 41701 6561 41735
rect 6595 41701 6607 41735
rect 6549 41695 6607 41701
rect 6917 41735 6975 41741
rect 6917 41701 6929 41735
rect 6963 41701 6975 41735
rect 7392 41732 7420 41760
rect 7392 41704 7880 41732
rect 6917 41695 6975 41701
rect 2924 41636 4016 41664
rect 4264 41636 5028 41664
rect 2924 41624 2930 41636
rect 2685 41599 2743 41605
rect 1504 41568 2636 41596
rect 1504 41537 1532 41568
rect 1489 41531 1547 41537
rect 1489 41497 1501 41531
rect 1535 41497 1547 41531
rect 1489 41491 1547 41497
rect 1762 41488 1768 41540
rect 1820 41528 1826 41540
rect 2041 41531 2099 41537
rect 2041 41528 2053 41531
rect 1820 41500 2053 41528
rect 1820 41488 1826 41500
rect 2041 41497 2053 41500
rect 2087 41497 2099 41531
rect 2608 41528 2636 41568
rect 2685 41565 2697 41599
rect 2731 41565 2743 41599
rect 2685 41559 2743 41565
rect 3142 41556 3148 41608
rect 3200 41596 3206 41608
rect 3329 41599 3387 41605
rect 3329 41596 3341 41599
rect 3200 41568 3341 41596
rect 3200 41556 3206 41568
rect 3329 41565 3341 41568
rect 3375 41565 3387 41599
rect 3329 41559 3387 41565
rect 3418 41556 3424 41608
rect 3476 41596 3482 41608
rect 3988 41605 4016 41636
rect 3605 41599 3663 41605
rect 3605 41596 3617 41599
rect 3476 41568 3617 41596
rect 3476 41556 3482 41568
rect 3605 41565 3617 41568
rect 3651 41565 3663 41599
rect 3605 41559 3663 41565
rect 3973 41599 4031 41605
rect 3973 41565 3985 41599
rect 4019 41565 4031 41599
rect 3973 41559 4031 41565
rect 4246 41556 4252 41608
rect 4304 41556 4310 41608
rect 4522 41556 4528 41608
rect 4580 41556 4586 41608
rect 4798 41556 4804 41608
rect 4856 41556 4862 41608
rect 4890 41528 4896 41540
rect 2608 41500 3740 41528
rect 2041 41491 2099 41497
rect 566 41420 572 41472
rect 624 41460 630 41472
rect 2682 41460 2688 41472
rect 624 41432 2688 41460
rect 624 41420 630 41432
rect 2682 41420 2688 41432
rect 2740 41420 2746 41472
rect 2866 41420 2872 41472
rect 2924 41460 2930 41472
rect 2961 41463 3019 41469
rect 2961 41460 2973 41463
rect 2924 41432 2973 41460
rect 2924 41420 2930 41432
rect 2961 41429 2973 41432
rect 3007 41460 3019 41463
rect 3142 41460 3148 41472
rect 3007 41432 3148 41460
rect 3007 41429 3019 41432
rect 2961 41423 3019 41429
rect 3142 41420 3148 41432
rect 3200 41420 3206 41472
rect 3712 41460 3740 41500
rect 4632 41500 4896 41528
rect 4632 41460 4660 41500
rect 4890 41488 4896 41500
rect 4948 41488 4954 41540
rect 3712 41432 4660 41460
rect 5000 41460 5028 41636
rect 5166 41624 5172 41676
rect 5224 41664 5230 41676
rect 6564 41664 6592 41695
rect 5224 41636 5948 41664
rect 5224 41624 5230 41636
rect 5077 41599 5135 41605
rect 5077 41565 5089 41599
rect 5123 41565 5135 41599
rect 5077 41559 5135 41565
rect 5092 41528 5120 41559
rect 5350 41556 5356 41608
rect 5408 41556 5414 41608
rect 5629 41599 5687 41605
rect 5629 41565 5641 41599
rect 5675 41596 5687 41599
rect 5810 41596 5816 41608
rect 5675 41568 5816 41596
rect 5675 41565 5687 41568
rect 5629 41559 5687 41565
rect 5810 41556 5816 41568
rect 5868 41556 5874 41608
rect 5920 41605 5948 41636
rect 6012 41636 6592 41664
rect 6932 41664 6960 41695
rect 6932 41636 7420 41664
rect 5905 41599 5963 41605
rect 5905 41565 5917 41599
rect 5951 41565 5963 41599
rect 5905 41559 5963 41565
rect 6012 41528 6040 41636
rect 7392 41605 7420 41636
rect 7558 41624 7564 41676
rect 7616 41664 7622 41676
rect 7616 41636 7788 41664
rect 7616 41624 7622 41636
rect 7760 41605 7788 41636
rect 6733 41599 6791 41605
rect 6733 41596 6745 41599
rect 5092 41500 6040 41528
rect 6196 41568 6745 41596
rect 5169 41463 5227 41469
rect 5169 41460 5181 41463
rect 5000 41432 5181 41460
rect 5169 41429 5181 41432
rect 5215 41429 5227 41463
rect 5169 41423 5227 41429
rect 6086 41420 6092 41472
rect 6144 41460 6150 41472
rect 6196 41469 6224 41568
rect 6733 41565 6745 41568
rect 6779 41565 6791 41599
rect 6733 41559 6791 41565
rect 7101 41599 7159 41605
rect 7101 41565 7113 41599
rect 7147 41565 7159 41599
rect 7101 41559 7159 41565
rect 7377 41599 7435 41605
rect 7377 41565 7389 41599
rect 7423 41565 7435 41599
rect 7377 41559 7435 41565
rect 7745 41599 7803 41605
rect 7745 41565 7757 41599
rect 7791 41565 7803 41599
rect 7852 41596 7880 41704
rect 7944 41664 7972 41760
rect 7944 41636 8340 41664
rect 8312 41605 8340 41636
rect 8021 41599 8079 41605
rect 8021 41596 8033 41599
rect 7852 41568 8033 41596
rect 7745 41559 7803 41565
rect 8021 41565 8033 41568
rect 8067 41565 8079 41599
rect 8021 41559 8079 41565
rect 8297 41599 8355 41605
rect 8297 41565 8309 41599
rect 8343 41565 8355 41599
rect 8297 41559 8355 41565
rect 7116 41528 7144 41559
rect 8570 41556 8576 41608
rect 8628 41556 8634 41608
rect 8864 41596 8892 41760
rect 10689 41735 10747 41741
rect 10689 41701 10701 41735
rect 10735 41701 10747 41735
rect 10689 41695 10747 41701
rect 10502 41624 10508 41676
rect 10560 41664 10566 41676
rect 10704 41664 10732 41695
rect 17954 41692 17960 41744
rect 18012 41692 18018 41744
rect 18156 41732 18184 41772
rect 18230 41760 18236 41812
rect 18288 41800 18294 41812
rect 18785 41803 18843 41809
rect 18785 41800 18797 41803
rect 18288 41772 18797 41800
rect 18288 41760 18294 41772
rect 18785 41769 18797 41772
rect 18831 41769 18843 41803
rect 18785 41763 18843 41769
rect 19150 41760 19156 41812
rect 19208 41760 19214 41812
rect 19426 41760 19432 41812
rect 19484 41800 19490 41812
rect 19613 41803 19671 41809
rect 19613 41800 19625 41803
rect 19484 41772 19625 41800
rect 19484 41760 19490 41772
rect 19613 41769 19625 41772
rect 19659 41769 19671 41803
rect 19613 41763 19671 41769
rect 19702 41760 19708 41812
rect 19760 41800 19766 41812
rect 19760 41772 20668 41800
rect 19760 41760 19766 41772
rect 19168 41732 19196 41760
rect 18156 41704 19196 41732
rect 19337 41735 19395 41741
rect 19337 41701 19349 41735
rect 19383 41732 19395 41735
rect 19383 41704 20208 41732
rect 19383 41701 19395 41704
rect 19337 41695 19395 41701
rect 10560 41636 10732 41664
rect 10796 41636 19564 41664
rect 10560 41624 10566 41636
rect 9125 41599 9183 41605
rect 9125 41596 9137 41599
rect 8864 41568 9137 41596
rect 9125 41565 9137 41568
rect 9171 41565 9183 41599
rect 9125 41559 9183 41565
rect 9674 41556 9680 41608
rect 9732 41556 9738 41608
rect 9858 41556 9864 41608
rect 9916 41596 9922 41608
rect 9951 41599 10009 41605
rect 9951 41596 9963 41599
rect 9916 41568 9963 41596
rect 9916 41556 9922 41568
rect 9951 41565 9963 41568
rect 9997 41596 10009 41599
rect 10796 41596 10824 41636
rect 9997 41568 10824 41596
rect 18141 41599 18199 41605
rect 9997 41565 10009 41568
rect 9951 41559 10009 41565
rect 18141 41565 18153 41599
rect 18187 41596 18199 41599
rect 18230 41596 18236 41608
rect 18187 41568 18236 41596
rect 18187 41565 18199 41568
rect 18141 41559 18199 41565
rect 18230 41556 18236 41568
rect 18288 41556 18294 41608
rect 18325 41599 18383 41605
rect 18325 41565 18337 41599
rect 18371 41596 18383 41599
rect 18414 41596 18420 41608
rect 18371 41568 18420 41596
rect 18371 41565 18383 41568
rect 18325 41559 18383 41565
rect 18414 41556 18420 41568
rect 18472 41556 18478 41608
rect 18966 41556 18972 41608
rect 19024 41556 19030 41608
rect 19536 41605 19564 41636
rect 20180 41605 20208 41704
rect 20438 41692 20444 41744
rect 20496 41692 20502 41744
rect 20530 41692 20536 41744
rect 20588 41692 20594 41744
rect 20456 41605 20484 41692
rect 20548 41605 20576 41692
rect 19521 41599 19579 41605
rect 19521 41565 19533 41599
rect 19567 41565 19579 41599
rect 19521 41559 19579 41565
rect 19797 41599 19855 41605
rect 19797 41565 19809 41599
rect 19843 41565 19855 41599
rect 19797 41559 19855 41565
rect 20165 41599 20223 41605
rect 20165 41565 20177 41599
rect 20211 41565 20223 41599
rect 20165 41559 20223 41565
rect 20441 41599 20499 41605
rect 20441 41565 20453 41599
rect 20487 41565 20499 41599
rect 20441 41559 20499 41565
rect 20533 41599 20591 41605
rect 20533 41565 20545 41599
rect 20579 41565 20591 41599
rect 20640 41596 20668 41772
rect 20714 41760 20720 41812
rect 20772 41760 20778 41812
rect 20806 41760 20812 41812
rect 20864 41800 20870 41812
rect 20864 41772 21036 41800
rect 20864 41760 20870 41772
rect 20901 41735 20959 41741
rect 20901 41701 20913 41735
rect 20947 41701 20959 41735
rect 21008 41732 21036 41772
rect 21082 41760 21088 41812
rect 21140 41800 21146 41812
rect 22922 41800 22928 41812
rect 21140 41772 22928 41800
rect 21140 41760 21146 41772
rect 22922 41760 22928 41772
rect 22980 41760 22986 41812
rect 23017 41803 23075 41809
rect 23017 41769 23029 41803
rect 23063 41800 23075 41803
rect 23658 41800 23664 41812
rect 23063 41772 23664 41800
rect 23063 41769 23075 41772
rect 23017 41763 23075 41769
rect 23658 41760 23664 41772
rect 23716 41760 23722 41812
rect 24121 41803 24179 41809
rect 24121 41769 24133 41803
rect 24167 41800 24179 41803
rect 25314 41800 25320 41812
rect 24167 41772 25320 41800
rect 24167 41769 24179 41772
rect 24121 41763 24179 41769
rect 25314 41760 25320 41772
rect 25372 41760 25378 41812
rect 21634 41732 21640 41744
rect 21008 41704 21640 41732
rect 20901 41695 20959 41701
rect 20916 41664 20944 41695
rect 21634 41692 21640 41704
rect 21692 41692 21698 41744
rect 21818 41692 21824 41744
rect 21876 41732 21882 41744
rect 23569 41735 23627 41741
rect 21876 41704 23336 41732
rect 21876 41692 21882 41704
rect 20916 41636 21956 41664
rect 21085 41599 21143 41605
rect 21085 41596 21097 41599
rect 20640 41568 21097 41596
rect 20533 41559 20591 41565
rect 21085 41565 21097 41568
rect 21131 41565 21143 41599
rect 21361 41599 21419 41605
rect 21361 41596 21373 41599
rect 21085 41559 21143 41565
rect 21192 41568 21373 41596
rect 10594 41528 10600 41540
rect 7116 41500 10600 41528
rect 10594 41488 10600 41500
rect 10652 41488 10658 41540
rect 17954 41488 17960 41540
rect 18012 41528 18018 41540
rect 19426 41528 19432 41540
rect 18012 41500 19432 41528
rect 18012 41488 18018 41500
rect 19426 41488 19432 41500
rect 19484 41488 19490 41540
rect 6181 41463 6239 41469
rect 6181 41460 6193 41463
rect 6144 41432 6193 41460
rect 6144 41420 6150 41432
rect 6181 41429 6193 41432
rect 6227 41429 6239 41463
rect 6181 41423 6239 41429
rect 7190 41420 7196 41472
rect 7248 41460 7254 41472
rect 7837 41463 7895 41469
rect 7837 41460 7849 41463
rect 7248 41432 7849 41460
rect 7248 41420 7254 41432
rect 7837 41429 7849 41432
rect 7883 41429 7895 41463
rect 7837 41423 7895 41429
rect 9950 41420 9956 41472
rect 10008 41460 10014 41472
rect 18138 41460 18144 41472
rect 10008 41432 18144 41460
rect 10008 41420 10014 41432
rect 18138 41420 18144 41432
rect 18196 41420 18202 41472
rect 18414 41420 18420 41472
rect 18472 41420 18478 41472
rect 19334 41420 19340 41472
rect 19392 41460 19398 41472
rect 19812 41460 19840 41559
rect 21192 41528 21220 41568
rect 21361 41565 21373 41568
rect 21407 41565 21419 41599
rect 21361 41559 21419 41565
rect 21634 41556 21640 41608
rect 21692 41556 21698 41608
rect 21928 41605 21956 41636
rect 22278 41624 22284 41676
rect 22336 41664 22342 41676
rect 22465 41667 22523 41673
rect 22465 41664 22477 41667
rect 22336 41636 22477 41664
rect 22336 41624 22342 41636
rect 22465 41633 22477 41636
rect 22511 41633 22523 41667
rect 22465 41627 22523 41633
rect 21913 41599 21971 41605
rect 21913 41565 21925 41599
rect 21959 41565 21971 41599
rect 21913 41559 21971 41565
rect 22066 41568 22508 41596
rect 22066 41528 22094 41568
rect 19996 41500 21220 41528
rect 21376 41500 22094 41528
rect 22189 41531 22247 41537
rect 19996 41469 20024 41500
rect 19392 41432 19840 41460
rect 19981 41463 20039 41469
rect 19392 41420 19398 41432
rect 19981 41429 19993 41463
rect 20027 41429 20039 41463
rect 19981 41423 20039 41429
rect 20254 41420 20260 41472
rect 20312 41420 20318 41472
rect 21177 41463 21235 41469
rect 21177 41429 21189 41463
rect 21223 41460 21235 41463
rect 21376 41460 21404 41500
rect 22189 41497 22201 41531
rect 22235 41528 22247 41531
rect 22370 41528 22376 41540
rect 22235 41500 22376 41528
rect 22235 41497 22247 41500
rect 22189 41491 22247 41497
rect 22370 41488 22376 41500
rect 22428 41488 22434 41540
rect 22480 41528 22508 41568
rect 22646 41528 22652 41540
rect 22480 41500 22652 41528
rect 22646 41488 22652 41500
rect 22704 41488 22710 41540
rect 22741 41531 22799 41537
rect 22741 41497 22753 41531
rect 22787 41528 22799 41531
rect 22922 41528 22928 41540
rect 22787 41500 22928 41528
rect 22787 41497 22799 41500
rect 22741 41491 22799 41497
rect 22922 41488 22928 41500
rect 22980 41488 22986 41540
rect 23308 41537 23336 41704
rect 23569 41701 23581 41735
rect 23615 41732 23627 41735
rect 25222 41732 25228 41744
rect 23615 41704 25228 41732
rect 23615 41701 23627 41704
rect 23569 41695 23627 41701
rect 25222 41692 25228 41704
rect 25280 41692 25286 41744
rect 23293 41531 23351 41537
rect 23293 41497 23305 41531
rect 23339 41497 23351 41531
rect 23293 41491 23351 41497
rect 23842 41488 23848 41540
rect 23900 41488 23906 41540
rect 21223 41432 21404 41460
rect 21223 41429 21235 41432
rect 21177 41423 21235 41429
rect 21450 41420 21456 41472
rect 21508 41420 21514 41472
rect 21729 41463 21787 41469
rect 21729 41429 21741 41463
rect 21775 41460 21787 41463
rect 22002 41460 22008 41472
rect 21775 41432 22008 41460
rect 21775 41429 21787 41432
rect 21729 41423 21787 41429
rect 22002 41420 22008 41432
rect 22060 41420 22066 41472
rect 22554 41420 22560 41472
rect 22612 41460 22618 41472
rect 25498 41460 25504 41472
rect 22612 41432 25504 41460
rect 22612 41420 22618 41432
rect 25498 41420 25504 41432
rect 25556 41420 25562 41472
rect 1104 41370 25000 41392
rect 1104 41318 6884 41370
rect 6936 41318 6948 41370
rect 7000 41318 7012 41370
rect 7064 41318 7076 41370
rect 7128 41318 7140 41370
rect 7192 41318 12818 41370
rect 12870 41318 12882 41370
rect 12934 41318 12946 41370
rect 12998 41318 13010 41370
rect 13062 41318 13074 41370
rect 13126 41318 18752 41370
rect 18804 41318 18816 41370
rect 18868 41318 18880 41370
rect 18932 41318 18944 41370
rect 18996 41318 19008 41370
rect 19060 41318 24686 41370
rect 24738 41318 24750 41370
rect 24802 41318 24814 41370
rect 24866 41318 24878 41370
rect 24930 41318 24942 41370
rect 24994 41318 25000 41370
rect 1104 41296 25000 41318
rect 2406 41216 2412 41268
rect 2464 41256 2470 41268
rect 2685 41259 2743 41265
rect 2685 41256 2697 41259
rect 2464 41228 2697 41256
rect 2464 41216 2470 41228
rect 2685 41225 2697 41228
rect 2731 41225 2743 41259
rect 2685 41219 2743 41225
rect 2774 41216 2780 41268
rect 2832 41256 2838 41268
rect 7558 41256 7564 41268
rect 2832 41228 7564 41256
rect 2832 41216 2838 41228
rect 7558 41216 7564 41228
rect 7616 41216 7622 41268
rect 7745 41259 7803 41265
rect 7745 41225 7757 41259
rect 7791 41256 7803 41259
rect 7834 41256 7840 41268
rect 7791 41228 7840 41256
rect 7791 41225 7803 41228
rect 7745 41219 7803 41225
rect 7834 41216 7840 41228
rect 7892 41216 7898 41268
rect 8018 41216 8024 41268
rect 8076 41256 8082 41268
rect 14642 41256 14648 41268
rect 8076 41228 14648 41256
rect 8076 41216 8082 41228
rect 14642 41216 14648 41228
rect 14700 41256 14706 41268
rect 15102 41256 15108 41268
rect 14700 41228 15108 41256
rect 14700 41216 14706 41228
rect 15102 41216 15108 41228
rect 15160 41216 15166 41268
rect 19521 41259 19579 41265
rect 19521 41225 19533 41259
rect 19567 41225 19579 41259
rect 19521 41219 19579 41225
rect 5534 41188 5540 41200
rect 4908 41160 5540 41188
rect 1210 41080 1216 41132
rect 1268 41120 1274 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 1268 41092 1409 41120
rect 1268 41080 1274 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 1397 41083 1455 41089
rect 2222 41080 2228 41132
rect 2280 41080 2286 41132
rect 2501 41123 2559 41129
rect 2501 41089 2513 41123
rect 2547 41120 2559 41123
rect 2547 41092 2774 41120
rect 2547 41089 2559 41092
rect 2501 41083 2559 41089
rect 2746 40984 2774 41092
rect 3234 41080 3240 41132
rect 3292 41080 3298 41132
rect 3786 41120 3792 41132
rect 3747 41092 3792 41120
rect 3786 41080 3792 41092
rect 3844 41080 3850 41132
rect 4908 41129 4936 41160
rect 5534 41148 5540 41160
rect 5592 41148 5598 41200
rect 12434 41188 12440 41200
rect 9140 41160 12440 41188
rect 4893 41123 4951 41129
rect 4893 41089 4905 41123
rect 4939 41089 4951 41123
rect 4893 41083 4951 41089
rect 5167 41123 5225 41129
rect 5167 41089 5179 41123
rect 5213 41120 5225 41123
rect 5213 41092 7880 41120
rect 5213 41089 5225 41092
rect 5167 41083 5225 41089
rect 3510 41012 3516 41064
rect 3568 41012 3574 41064
rect 3053 40987 3111 40993
rect 3053 40984 3065 40987
rect 2746 40956 3065 40984
rect 3053 40953 3065 40956
rect 3099 40953 3111 40987
rect 3053 40947 3111 40953
rect 4448 40956 5028 40984
rect 2866 40876 2872 40928
rect 2924 40916 2930 40928
rect 4448 40916 4476 40956
rect 2924 40888 4476 40916
rect 2924 40876 2930 40888
rect 4522 40876 4528 40928
rect 4580 40876 4586 40928
rect 5000 40916 5028 40956
rect 5828 40956 6868 40984
rect 5828 40916 5856 40956
rect 5000 40888 5856 40916
rect 5905 40919 5963 40925
rect 5905 40885 5917 40919
rect 5951 40916 5963 40919
rect 5994 40916 6000 40928
rect 5951 40888 6000 40916
rect 5951 40885 5963 40888
rect 5905 40879 5963 40885
rect 5994 40876 6000 40888
rect 6052 40876 6058 40928
rect 6840 40916 6868 40956
rect 6914 40944 6920 40996
rect 6972 40984 6978 40996
rect 6972 40956 7788 40984
rect 6972 40944 6978 40956
rect 7760 40928 7788 40956
rect 7852 40928 7880 41092
rect 7926 41080 7932 41132
rect 7984 41080 7990 41132
rect 9140 41130 9168 41160
rect 12434 41148 12440 41160
rect 12492 41148 12498 41200
rect 8847 41123 8905 41129
rect 8847 41089 8859 41123
rect 8893 41120 8905 41123
rect 9048 41120 9168 41130
rect 8893 41102 9168 41120
rect 8893 41092 9076 41102
rect 8893 41089 8905 41092
rect 8847 41083 8905 41089
rect 9674 41080 9680 41132
rect 9732 41120 9738 41132
rect 10045 41123 10103 41129
rect 10045 41120 10057 41123
rect 9732 41092 10057 41120
rect 9732 41080 9738 41092
rect 10045 41089 10057 41092
rect 10091 41089 10103 41123
rect 10045 41083 10103 41089
rect 10319 41123 10377 41129
rect 10319 41089 10331 41123
rect 10365 41120 10377 41123
rect 10410 41120 10416 41132
rect 10365 41092 10416 41120
rect 10365 41089 10377 41092
rect 10319 41083 10377 41089
rect 10410 41080 10416 41092
rect 10468 41080 10474 41132
rect 19245 41123 19303 41129
rect 19245 41089 19257 41123
rect 19291 41120 19303 41123
rect 19536 41120 19564 41219
rect 19794 41216 19800 41268
rect 19852 41216 19858 41268
rect 20346 41216 20352 41268
rect 20404 41216 20410 41268
rect 20622 41216 20628 41268
rect 20680 41216 20686 41268
rect 20901 41259 20959 41265
rect 20901 41225 20913 41259
rect 20947 41256 20959 41259
rect 21174 41256 21180 41268
rect 20947 41228 21180 41256
rect 20947 41225 20959 41228
rect 20901 41219 20959 41225
rect 21174 41216 21180 41228
rect 21232 41216 21238 41268
rect 21266 41216 21272 41268
rect 21324 41256 21330 41268
rect 21453 41259 21511 41265
rect 21453 41256 21465 41259
rect 21324 41228 21465 41256
rect 21324 41216 21330 41228
rect 21453 41225 21465 41228
rect 21499 41225 21511 41259
rect 21821 41259 21879 41265
rect 21821 41256 21833 41259
rect 21453 41219 21511 41225
rect 21560 41228 21833 41256
rect 19291 41092 19564 41120
rect 19291 41089 19303 41092
rect 19245 41083 19303 41089
rect 19702 41080 19708 41132
rect 19760 41080 19766 41132
rect 19886 41080 19892 41132
rect 19944 41120 19950 41132
rect 19981 41123 20039 41129
rect 19981 41120 19993 41123
rect 19944 41092 19993 41120
rect 19944 41080 19950 41092
rect 19981 41089 19993 41092
rect 20027 41089 20039 41123
rect 19981 41083 20039 41089
rect 20257 41123 20315 41129
rect 20257 41089 20269 41123
rect 20303 41089 20315 41123
rect 20257 41083 20315 41089
rect 8570 41012 8576 41064
rect 8628 41012 8634 41064
rect 9490 41012 9496 41064
rect 9548 41052 9554 41064
rect 11698 41052 11704 41064
rect 9548 41024 9994 41052
rect 9548 41012 9554 41024
rect 9858 40984 9864 40996
rect 9508 40956 9864 40984
rect 7374 40916 7380 40928
rect 6840 40888 7380 40916
rect 7374 40876 7380 40888
rect 7432 40876 7438 40928
rect 7466 40876 7472 40928
rect 7524 40876 7530 40928
rect 7742 40876 7748 40928
rect 7800 40876 7806 40928
rect 7834 40876 7840 40928
rect 7892 40916 7898 40928
rect 9508 40916 9536 40956
rect 9858 40944 9864 40956
rect 9916 40944 9922 40996
rect 7892 40888 9536 40916
rect 7892 40876 7898 40888
rect 9582 40876 9588 40928
rect 9640 40876 9646 40928
rect 9966 40916 9994 41024
rect 10704 41024 11704 41052
rect 10704 40916 10732 41024
rect 11698 41012 11704 41024
rect 11756 41012 11762 41064
rect 16390 41012 16396 41064
rect 16448 41052 16454 41064
rect 20272 41052 20300 41083
rect 20530 41080 20536 41132
rect 20588 41080 20594 41132
rect 20622 41080 20628 41132
rect 20680 41120 20686 41132
rect 20809 41123 20867 41129
rect 20809 41120 20821 41123
rect 20680 41092 20821 41120
rect 20680 41080 20686 41092
rect 20809 41089 20821 41092
rect 20855 41089 20867 41123
rect 20809 41083 20867 41089
rect 21085 41123 21143 41129
rect 21085 41089 21097 41123
rect 21131 41120 21143 41123
rect 21174 41120 21180 41132
rect 21131 41092 21180 41120
rect 21131 41089 21143 41092
rect 21085 41083 21143 41089
rect 21174 41080 21180 41092
rect 21232 41080 21238 41132
rect 21266 41080 21272 41132
rect 21324 41120 21330 41132
rect 21361 41123 21419 41129
rect 21361 41120 21373 41123
rect 21324 41092 21373 41120
rect 21324 41080 21330 41092
rect 21361 41089 21373 41092
rect 21407 41089 21419 41123
rect 21361 41083 21419 41089
rect 16448 41024 20300 41052
rect 16448 41012 16454 41024
rect 20438 41012 20444 41064
rect 20496 41012 20502 41064
rect 20714 41012 20720 41064
rect 20772 41052 20778 41064
rect 21560 41052 21588 41228
rect 21821 41225 21833 41228
rect 21867 41225 21879 41259
rect 21821 41219 21879 41225
rect 22002 41216 22008 41268
rect 22060 41216 22066 41268
rect 22097 41259 22155 41265
rect 22097 41225 22109 41259
rect 22143 41256 22155 41259
rect 22462 41256 22468 41268
rect 22143 41228 22468 41256
rect 22143 41225 22155 41228
rect 22097 41219 22155 41225
rect 22462 41216 22468 41228
rect 22520 41216 22526 41268
rect 23109 41259 23167 41265
rect 23109 41225 23121 41259
rect 23155 41256 23167 41259
rect 23382 41256 23388 41268
rect 23155 41228 23388 41256
rect 23155 41225 23167 41228
rect 23109 41219 23167 41225
rect 23382 41216 23388 41228
rect 23440 41216 23446 41268
rect 24213 41259 24271 41265
rect 24213 41225 24225 41259
rect 24259 41256 24271 41259
rect 25038 41256 25044 41268
rect 24259 41228 25044 41256
rect 24259 41225 24271 41228
rect 24213 41219 24271 41225
rect 25038 41216 25044 41228
rect 25096 41216 25102 41268
rect 22020 41188 22048 41216
rect 22020 41160 22968 41188
rect 21637 41123 21695 41129
rect 21637 41089 21649 41123
rect 21683 41120 21695 41123
rect 21683 41092 21772 41120
rect 21683 41089 21695 41092
rect 21637 41083 21695 41089
rect 20772 41024 21588 41052
rect 21744 41052 21772 41092
rect 21818 41080 21824 41132
rect 21876 41120 21882 41132
rect 22005 41123 22063 41129
rect 22005 41120 22017 41123
rect 21876 41092 22017 41120
rect 21876 41080 21882 41092
rect 22005 41089 22017 41092
rect 22051 41089 22063 41123
rect 22005 41083 22063 41089
rect 22186 41080 22192 41132
rect 22244 41124 22250 41132
rect 22281 41124 22339 41129
rect 22244 41123 22339 41124
rect 22244 41096 22293 41123
rect 22244 41080 22250 41096
rect 22281 41089 22293 41096
rect 22327 41089 22339 41123
rect 22281 41083 22339 41089
rect 22462 41080 22468 41132
rect 22520 41120 22526 41132
rect 22557 41123 22615 41129
rect 22557 41120 22569 41123
rect 22520 41092 22569 41120
rect 22520 41080 22526 41092
rect 22557 41089 22569 41092
rect 22603 41089 22615 41123
rect 22557 41083 22615 41089
rect 22833 41123 22891 41129
rect 22833 41089 22845 41123
rect 22879 41089 22891 41123
rect 22833 41083 22891 41089
rect 22738 41052 22744 41064
rect 21744 41024 22744 41052
rect 20772 41012 20778 41024
rect 22738 41012 22744 41024
rect 22796 41012 22802 41064
rect 20073 40987 20131 40993
rect 20073 40953 20085 40987
rect 20119 40984 20131 40987
rect 20456 40984 20484 41012
rect 20119 40956 20484 40984
rect 20548 40956 21588 40984
rect 20119 40953 20131 40956
rect 20073 40947 20131 40953
rect 9966 40888 10732 40916
rect 11054 40876 11060 40928
rect 11112 40876 11118 40928
rect 19058 40876 19064 40928
rect 19116 40876 19122 40928
rect 20438 40876 20444 40928
rect 20496 40916 20502 40928
rect 20548 40916 20576 40956
rect 20496 40888 20576 40916
rect 21177 40919 21235 40925
rect 20496 40876 20502 40888
rect 21177 40885 21189 40919
rect 21223 40916 21235 40919
rect 21450 40916 21456 40928
rect 21223 40888 21456 40916
rect 21223 40885 21235 40888
rect 21177 40879 21235 40885
rect 21450 40876 21456 40888
rect 21508 40876 21514 40928
rect 21560 40916 21588 40956
rect 21634 40944 21640 40996
rect 21692 40984 21698 40996
rect 22848 40984 22876 41083
rect 22940 41052 22968 41160
rect 23474 41148 23480 41200
rect 23532 41188 23538 41200
rect 23937 41191 23995 41197
rect 23937 41188 23949 41191
rect 23532 41160 23949 41188
rect 23532 41148 23538 41160
rect 23937 41157 23949 41160
rect 23983 41157 23995 41191
rect 23937 41151 23995 41157
rect 23106 41080 23112 41132
rect 23164 41120 23170 41132
rect 23385 41123 23443 41129
rect 23385 41120 23397 41123
rect 23164 41092 23397 41120
rect 23164 41080 23170 41092
rect 23385 41089 23397 41092
rect 23431 41089 23443 41123
rect 23385 41083 23443 41089
rect 23290 41052 23296 41064
rect 22940 41024 23296 41052
rect 23290 41012 23296 41024
rect 23348 41012 23354 41064
rect 21692 40956 22876 40984
rect 21692 40944 21698 40956
rect 21726 40916 21732 40928
rect 21560 40888 21732 40916
rect 21726 40876 21732 40888
rect 21784 40876 21790 40928
rect 22094 40876 22100 40928
rect 22152 40916 22158 40928
rect 22373 40919 22431 40925
rect 22373 40916 22385 40919
rect 22152 40888 22385 40916
rect 22152 40876 22158 40888
rect 22373 40885 22385 40888
rect 22419 40885 22431 40919
rect 22373 40879 22431 40885
rect 23658 40876 23664 40928
rect 23716 40876 23722 40928
rect 1104 40826 24840 40848
rect 1104 40774 3917 40826
rect 3969 40774 3981 40826
rect 4033 40774 4045 40826
rect 4097 40774 4109 40826
rect 4161 40774 4173 40826
rect 4225 40774 9851 40826
rect 9903 40774 9915 40826
rect 9967 40774 9979 40826
rect 10031 40774 10043 40826
rect 10095 40774 10107 40826
rect 10159 40774 15785 40826
rect 15837 40774 15849 40826
rect 15901 40774 15913 40826
rect 15965 40774 15977 40826
rect 16029 40774 16041 40826
rect 16093 40774 21719 40826
rect 21771 40774 21783 40826
rect 21835 40774 21847 40826
rect 21899 40774 21911 40826
rect 21963 40774 21975 40826
rect 22027 40774 24840 40826
rect 1104 40752 24840 40774
rect 2774 40712 2780 40724
rect 2746 40672 2780 40712
rect 2832 40672 2838 40724
rect 3050 40672 3056 40724
rect 3108 40712 3114 40724
rect 3421 40715 3479 40721
rect 3421 40712 3433 40715
rect 3108 40684 3433 40712
rect 3108 40672 3114 40684
rect 3421 40681 3433 40684
rect 3467 40681 3479 40715
rect 3421 40675 3479 40681
rect 3786 40672 3792 40724
rect 3844 40712 3850 40724
rect 8018 40712 8024 40724
rect 3844 40684 8024 40712
rect 3844 40672 3850 40684
rect 2225 40579 2283 40585
rect 2225 40545 2237 40579
rect 2271 40576 2283 40579
rect 2746 40576 2774 40672
rect 4798 40604 4804 40656
rect 4856 40604 4862 40656
rect 2271 40548 2774 40576
rect 2271 40545 2283 40548
rect 2225 40539 2283 40545
rect 3510 40536 3516 40588
rect 3568 40576 3574 40588
rect 3789 40579 3847 40585
rect 3789 40576 3801 40579
rect 3568 40548 3801 40576
rect 3568 40536 3574 40548
rect 3789 40545 3801 40548
rect 3835 40545 3847 40579
rect 3789 40539 3847 40545
rect 1854 40468 1860 40520
rect 1912 40508 1918 40520
rect 3605 40511 3663 40517
rect 3605 40508 3617 40511
rect 1912 40480 3617 40508
rect 1912 40468 1918 40480
rect 3605 40477 3617 40480
rect 3651 40477 3663 40511
rect 3605 40471 3663 40477
rect 1394 40400 1400 40452
rect 1452 40400 1458 40452
rect 2409 40443 2467 40449
rect 2409 40409 2421 40443
rect 2455 40440 2467 40443
rect 2774 40440 2780 40452
rect 2455 40412 2780 40440
rect 2455 40409 2467 40412
rect 2409 40403 2467 40409
rect 2774 40400 2780 40412
rect 2832 40400 2838 40452
rect 3050 40400 3056 40452
rect 3108 40440 3114 40452
rect 3145 40443 3203 40449
rect 3145 40440 3157 40443
rect 3108 40412 3157 40440
rect 3108 40400 3114 40412
rect 3145 40409 3157 40412
rect 3191 40409 3203 40443
rect 3804 40440 3832 40539
rect 5534 40536 5540 40588
rect 5592 40536 5598 40588
rect 3970 40468 3976 40520
rect 4028 40508 4034 40520
rect 4063 40511 4121 40517
rect 4063 40508 4075 40511
rect 4028 40480 4075 40508
rect 4028 40468 4034 40480
rect 4063 40477 4075 40480
rect 4109 40508 4121 40511
rect 5442 40508 5448 40520
rect 4109 40480 5448 40508
rect 4109 40477 4121 40480
rect 4063 40471 4121 40477
rect 5442 40468 5448 40480
rect 5500 40468 5506 40520
rect 5811 40511 5869 40517
rect 5811 40477 5823 40511
rect 5857 40508 5869 40511
rect 6196 40508 6224 40684
rect 8018 40672 8024 40684
rect 8076 40672 8082 40724
rect 10962 40712 10968 40724
rect 9140 40684 10968 40712
rect 5857 40480 6224 40508
rect 6917 40511 6975 40517
rect 5857 40477 5869 40480
rect 5811 40471 5869 40477
rect 6917 40477 6929 40511
rect 6963 40477 6975 40511
rect 6917 40471 6975 40477
rect 7191 40511 7249 40517
rect 7191 40477 7203 40511
rect 7237 40508 7249 40511
rect 7834 40508 7840 40520
rect 7237 40480 7840 40508
rect 7237 40477 7249 40480
rect 7191 40471 7249 40477
rect 6730 40440 6736 40452
rect 3804 40412 6736 40440
rect 3145 40403 3203 40409
rect 6730 40400 6736 40412
rect 6788 40440 6794 40452
rect 6932 40440 6960 40471
rect 7834 40468 7840 40480
rect 7892 40468 7898 40520
rect 6788 40412 6960 40440
rect 6788 40400 6794 40412
rect 7650 40400 7656 40452
rect 7708 40440 7714 40452
rect 9140 40440 9168 40684
rect 10318 40604 10324 40656
rect 10376 40604 10382 40656
rect 10502 40604 10508 40656
rect 10560 40604 10566 40656
rect 10045 40579 10103 40585
rect 10045 40545 10057 40579
rect 10091 40576 10103 40579
rect 10336 40576 10364 40604
rect 10091 40548 10364 40576
rect 10612 40576 10640 40684
rect 10962 40672 10968 40684
rect 11020 40672 11026 40724
rect 16390 40712 16396 40724
rect 11808 40684 16396 40712
rect 10612 40548 10916 40576
rect 10091 40545 10103 40548
rect 10045 40539 10103 40545
rect 9861 40511 9919 40517
rect 9861 40477 9873 40511
rect 9907 40477 9919 40511
rect 9861 40471 9919 40477
rect 7708 40412 9168 40440
rect 7708 40400 7714 40412
rect 9140 40384 9168 40412
rect 3694 40332 3700 40384
rect 3752 40372 3758 40384
rect 5074 40372 5080 40384
rect 3752 40344 5080 40372
rect 3752 40332 3758 40344
rect 5074 40332 5080 40344
rect 5132 40332 5138 40384
rect 6549 40375 6607 40381
rect 6549 40341 6561 40375
rect 6595 40372 6607 40375
rect 6638 40372 6644 40384
rect 6595 40344 6644 40372
rect 6595 40341 6607 40344
rect 6549 40335 6607 40341
rect 6638 40332 6644 40344
rect 6696 40332 6702 40384
rect 7926 40332 7932 40384
rect 7984 40332 7990 40384
rect 8018 40332 8024 40384
rect 8076 40372 8082 40384
rect 8386 40372 8392 40384
rect 8076 40344 8392 40372
rect 8076 40332 8082 40344
rect 8386 40332 8392 40344
rect 8444 40332 8450 40384
rect 8938 40332 8944 40384
rect 8996 40372 9002 40384
rect 9122 40372 9128 40384
rect 8996 40344 9128 40372
rect 8996 40332 9002 40344
rect 9122 40332 9128 40344
rect 9180 40332 9186 40384
rect 9876 40372 9904 40471
rect 10778 40468 10784 40520
rect 10836 40468 10842 40520
rect 10888 40517 10916 40548
rect 11054 40536 11060 40588
rect 11112 40536 11118 40588
rect 11606 40536 11612 40588
rect 11664 40576 11670 40588
rect 11808 40585 11836 40684
rect 16390 40672 16396 40684
rect 16448 40672 16454 40724
rect 19058 40672 19064 40724
rect 19116 40672 19122 40724
rect 20809 40715 20867 40721
rect 20809 40712 20821 40715
rect 20548 40684 20821 40712
rect 11793 40579 11851 40585
rect 11793 40576 11805 40579
rect 11664 40548 11805 40576
rect 11664 40536 11670 40548
rect 11793 40545 11805 40548
rect 11839 40545 11851 40579
rect 11793 40539 11851 40545
rect 10888 40511 10956 40517
rect 10888 40480 10910 40511
rect 10898 40477 10910 40480
rect 10944 40477 10956 40511
rect 10898 40471 10956 40477
rect 12051 40481 12109 40487
rect 12051 40447 12063 40481
rect 12097 40478 12109 40481
rect 12097 40447 12112 40478
rect 12710 40468 12716 40520
rect 12768 40508 12774 40520
rect 13357 40511 13415 40517
rect 13357 40508 13369 40511
rect 12768 40480 13369 40508
rect 12768 40468 12774 40480
rect 13357 40477 13369 40480
rect 13403 40477 13415 40511
rect 19076 40508 19104 40672
rect 19521 40647 19579 40653
rect 19521 40613 19533 40647
rect 19567 40644 19579 40647
rect 19702 40644 19708 40656
rect 19567 40616 19708 40644
rect 19567 40613 19579 40616
rect 19521 40607 19579 40613
rect 19702 40604 19708 40616
rect 19760 40604 19766 40656
rect 20254 40604 20260 40656
rect 20312 40604 20318 40656
rect 20438 40604 20444 40656
rect 20496 40644 20502 40656
rect 20548 40644 20576 40684
rect 20809 40681 20821 40684
rect 20855 40681 20867 40715
rect 20809 40675 20867 40681
rect 21082 40672 21088 40724
rect 21140 40672 21146 40724
rect 21266 40672 21272 40724
rect 21324 40712 21330 40724
rect 21726 40712 21732 40724
rect 21324 40684 21732 40712
rect 21324 40672 21330 40684
rect 21726 40672 21732 40684
rect 21784 40672 21790 40724
rect 22186 40672 22192 40724
rect 22244 40672 22250 40724
rect 22462 40672 22468 40724
rect 22520 40672 22526 40724
rect 22738 40672 22744 40724
rect 22796 40672 22802 40724
rect 23014 40672 23020 40724
rect 23072 40672 23078 40724
rect 23477 40715 23535 40721
rect 23477 40681 23489 40715
rect 23523 40712 23535 40715
rect 24026 40712 24032 40724
rect 23523 40684 24032 40712
rect 23523 40681 23535 40684
rect 23477 40675 23535 40681
rect 24026 40672 24032 40684
rect 24084 40672 24090 40724
rect 22002 40644 22008 40656
rect 20496 40616 20576 40644
rect 20732 40616 22008 40644
rect 20496 40604 20502 40616
rect 19242 40536 19248 40588
rect 19300 40576 19306 40588
rect 20732 40576 20760 40616
rect 22002 40604 22008 40616
rect 22060 40604 22066 40656
rect 21634 40576 21640 40588
rect 19300 40548 20116 40576
rect 19300 40536 19306 40548
rect 19337 40511 19395 40517
rect 19337 40508 19349 40511
rect 19076 40480 19349 40508
rect 13357 40471 13415 40477
rect 19337 40477 19349 40480
rect 19383 40477 19395 40511
rect 19337 40471 19395 40477
rect 19426 40468 19432 40520
rect 19484 40508 19490 40520
rect 19797 40511 19855 40517
rect 19797 40508 19809 40511
rect 19484 40480 19809 40508
rect 19484 40468 19490 40480
rect 19797 40477 19809 40480
rect 19843 40477 19855 40511
rect 19797 40471 19855 40477
rect 12051 40441 12112 40447
rect 12084 40440 12112 40441
rect 12434 40440 12440 40452
rect 12084 40412 12440 40440
rect 12434 40400 12440 40412
rect 12492 40400 12498 40452
rect 17402 40400 17408 40452
rect 17460 40440 17466 40452
rect 20088 40440 20116 40548
rect 20456 40548 20760 40576
rect 21192 40548 21640 40576
rect 20162 40468 20168 40520
rect 20220 40468 20226 40520
rect 20456 40517 20484 40548
rect 20441 40511 20499 40517
rect 20441 40477 20453 40511
rect 20487 40477 20499 40511
rect 20441 40471 20499 40477
rect 20717 40511 20775 40517
rect 20717 40477 20729 40511
rect 20763 40477 20775 40511
rect 20717 40471 20775 40477
rect 20993 40511 21051 40517
rect 20993 40477 21005 40511
rect 21039 40508 21051 40511
rect 21082 40508 21088 40520
rect 21039 40480 21088 40508
rect 21039 40477 21051 40480
rect 20993 40471 21051 40477
rect 20732 40440 20760 40471
rect 21082 40468 21088 40480
rect 21140 40468 21146 40520
rect 17460 40412 20024 40440
rect 20088 40412 20760 40440
rect 21192 40440 21220 40548
rect 21634 40536 21640 40548
rect 21692 40536 21698 40588
rect 21744 40548 22232 40576
rect 21269 40511 21327 40517
rect 21269 40477 21281 40511
rect 21315 40508 21327 40511
rect 21450 40508 21456 40520
rect 21315 40480 21456 40508
rect 21315 40477 21327 40480
rect 21269 40471 21327 40477
rect 21450 40468 21456 40480
rect 21508 40468 21514 40520
rect 21553 40511 21611 40517
rect 21553 40477 21565 40511
rect 21599 40508 21611 40511
rect 21744 40508 21772 40548
rect 21599 40480 21772 40508
rect 21821 40511 21879 40517
rect 21599 40477 21611 40480
rect 21553 40471 21611 40477
rect 21821 40477 21833 40511
rect 21867 40477 21879 40511
rect 21821 40471 21879 40477
rect 21836 40440 21864 40471
rect 22094 40468 22100 40520
rect 22152 40468 22158 40520
rect 21192 40412 21496 40440
rect 21836 40412 21956 40440
rect 17460 40400 17466 40412
rect 11146 40372 11152 40384
rect 9876 40344 11152 40372
rect 11146 40332 11152 40344
rect 11204 40332 11210 40384
rect 11701 40375 11759 40381
rect 11701 40341 11713 40375
rect 11747 40372 11759 40375
rect 12158 40372 12164 40384
rect 11747 40344 12164 40372
rect 11747 40341 11759 40344
rect 11701 40335 11759 40341
rect 12158 40332 12164 40344
rect 12216 40332 12222 40384
rect 12342 40332 12348 40384
rect 12400 40372 12406 40384
rect 12805 40375 12863 40381
rect 12805 40372 12817 40375
rect 12400 40344 12817 40372
rect 12400 40332 12406 40344
rect 12805 40341 12817 40344
rect 12851 40341 12863 40375
rect 12805 40335 12863 40341
rect 19610 40332 19616 40384
rect 19668 40332 19674 40384
rect 19996 40381 20024 40412
rect 19981 40375 20039 40381
rect 19981 40341 19993 40375
rect 20027 40341 20039 40375
rect 19981 40335 20039 40341
rect 20070 40332 20076 40384
rect 20128 40372 20134 40384
rect 20533 40375 20591 40381
rect 20533 40372 20545 40375
rect 20128 40344 20545 40372
rect 20128 40332 20134 40344
rect 20533 40341 20545 40344
rect 20579 40341 20591 40375
rect 20533 40335 20591 40341
rect 21266 40332 21272 40384
rect 21324 40372 21330 40384
rect 21361 40375 21419 40381
rect 21361 40372 21373 40375
rect 21324 40344 21373 40372
rect 21324 40332 21330 40344
rect 21361 40341 21373 40344
rect 21407 40341 21419 40375
rect 21468 40372 21496 40412
rect 21928 40381 21956 40412
rect 21637 40375 21695 40381
rect 21637 40372 21649 40375
rect 21468 40344 21649 40372
rect 21361 40335 21419 40341
rect 21637 40341 21649 40344
rect 21683 40341 21695 40375
rect 21637 40335 21695 40341
rect 21913 40375 21971 40381
rect 21913 40341 21925 40375
rect 21959 40341 21971 40375
rect 22204 40372 22232 40548
rect 22278 40536 22284 40588
rect 22336 40576 22342 40588
rect 23474 40576 23480 40588
rect 22336 40548 23480 40576
rect 22336 40536 22342 40548
rect 23474 40536 23480 40548
rect 23532 40536 23538 40588
rect 22373 40511 22431 40517
rect 22373 40477 22385 40511
rect 22419 40508 22431 40511
rect 22554 40508 22560 40520
rect 22419 40480 22560 40508
rect 22419 40477 22431 40480
rect 22373 40471 22431 40477
rect 22554 40468 22560 40480
rect 22612 40468 22618 40520
rect 22646 40468 22652 40520
rect 22704 40468 22710 40520
rect 22922 40468 22928 40520
rect 22980 40468 22986 40520
rect 23201 40511 23259 40517
rect 23201 40477 23213 40511
rect 23247 40508 23259 40511
rect 23290 40508 23296 40520
rect 23247 40480 23296 40508
rect 23247 40477 23259 40480
rect 23201 40471 23259 40477
rect 23290 40468 23296 40480
rect 23348 40468 23354 40520
rect 23658 40468 23664 40520
rect 23716 40468 23722 40520
rect 23014 40400 23020 40452
rect 23072 40440 23078 40452
rect 23845 40443 23903 40449
rect 23845 40440 23857 40443
rect 23072 40412 23857 40440
rect 23072 40400 23078 40412
rect 23845 40409 23857 40412
rect 23891 40409 23903 40443
rect 23845 40403 23903 40409
rect 24213 40443 24271 40449
rect 24213 40409 24225 40443
rect 24259 40440 24271 40443
rect 25130 40440 25136 40452
rect 24259 40412 25136 40440
rect 24259 40409 24271 40412
rect 24213 40403 24271 40409
rect 25130 40400 25136 40412
rect 25188 40400 25194 40452
rect 22922 40372 22928 40384
rect 22204 40344 22928 40372
rect 21913 40335 21971 40341
rect 22922 40332 22928 40344
rect 22980 40332 22986 40384
rect 23474 40332 23480 40384
rect 23532 40372 23538 40384
rect 25774 40372 25780 40384
rect 23532 40344 25780 40372
rect 23532 40332 23538 40344
rect 25774 40332 25780 40344
rect 25832 40332 25838 40384
rect 1104 40282 25000 40304
rect 1104 40230 6884 40282
rect 6936 40230 6948 40282
rect 7000 40230 7012 40282
rect 7064 40230 7076 40282
rect 7128 40230 7140 40282
rect 7192 40230 12818 40282
rect 12870 40230 12882 40282
rect 12934 40230 12946 40282
rect 12998 40230 13010 40282
rect 13062 40230 13074 40282
rect 13126 40230 18752 40282
rect 18804 40230 18816 40282
rect 18868 40230 18880 40282
rect 18932 40230 18944 40282
rect 18996 40230 19008 40282
rect 19060 40230 24686 40282
rect 24738 40230 24750 40282
rect 24802 40230 24814 40282
rect 24866 40230 24878 40282
rect 24930 40230 24942 40282
rect 24994 40230 25000 40282
rect 1104 40208 25000 40230
rect 2866 40168 2872 40180
rect 1688 40140 2872 40168
rect 1688 40109 1716 40140
rect 2866 40128 2872 40140
rect 2924 40128 2930 40180
rect 2958 40128 2964 40180
rect 3016 40168 3022 40180
rect 4157 40171 4215 40177
rect 4157 40168 4169 40171
rect 3016 40140 4169 40168
rect 3016 40128 3022 40140
rect 4157 40137 4169 40140
rect 4203 40137 4215 40171
rect 5166 40168 5172 40180
rect 4157 40131 4215 40137
rect 4816 40140 5172 40168
rect 1673 40103 1731 40109
rect 1673 40069 1685 40103
rect 1719 40069 1731 40103
rect 2222 40071 2228 40112
rect 1673 40063 1731 40069
rect 2207 40065 2228 40071
rect 1397 40035 1455 40041
rect 1397 40001 1409 40035
rect 1443 40032 1455 40035
rect 1486 40032 1492 40044
rect 1443 40004 1492 40032
rect 1443 40001 1455 40004
rect 1397 39995 1455 40001
rect 1486 39992 1492 40004
rect 1544 39992 1550 40044
rect 2207 40031 2219 40065
rect 2280 40060 2286 40112
rect 3605 40103 3663 40109
rect 3605 40069 3617 40103
rect 3651 40100 3663 40103
rect 4816 40100 4844 40140
rect 5166 40128 5172 40140
rect 5224 40128 5230 40180
rect 5442 40128 5448 40180
rect 5500 40168 5506 40180
rect 7282 40168 7288 40180
rect 5500 40140 7288 40168
rect 5500 40128 5506 40140
rect 5534 40100 5540 40112
rect 3651 40072 4844 40100
rect 4908 40072 5540 40100
rect 3651 40069 3663 40072
rect 3605 40063 3663 40069
rect 2253 40034 2268 40060
rect 2253 40031 2265 40034
rect 2207 40025 2265 40031
rect 2314 39992 2320 40044
rect 2372 40032 2378 40044
rect 3142 40032 3148 40044
rect 2372 40004 3148 40032
rect 2372 39992 2378 40004
rect 3142 39992 3148 40004
rect 3200 39992 3206 40044
rect 3329 40035 3387 40041
rect 3329 40001 3341 40035
rect 3375 40001 3387 40035
rect 3329 39995 3387 40001
rect 1762 39924 1768 39976
rect 1820 39964 1826 39976
rect 1949 39967 2007 39973
rect 1949 39964 1961 39967
rect 1820 39936 1961 39964
rect 1820 39924 1826 39936
rect 1949 39933 1961 39936
rect 1995 39933 2007 39967
rect 1949 39927 2007 39933
rect 3234 39924 3240 39976
rect 3292 39964 3298 39976
rect 3344 39964 3372 39995
rect 4338 39992 4344 40044
rect 4396 39992 4402 40044
rect 4908 40041 4936 40072
rect 5534 40060 5540 40072
rect 5592 40060 5598 40112
rect 4893 40035 4951 40041
rect 4893 40001 4905 40035
rect 4939 40001 4951 40035
rect 4893 39995 4951 40001
rect 5167 40035 5225 40041
rect 5167 40001 5179 40035
rect 5213 40032 5225 40035
rect 5644 40032 5672 40140
rect 7282 40128 7288 40140
rect 7340 40128 7346 40180
rect 7469 40171 7527 40177
rect 7469 40137 7481 40171
rect 7515 40168 7527 40171
rect 7650 40168 7656 40180
rect 7515 40140 7656 40168
rect 7515 40137 7527 40140
rect 7469 40131 7527 40137
rect 7650 40128 7656 40140
rect 7708 40128 7714 40180
rect 8573 40171 8631 40177
rect 7760 40140 8524 40168
rect 7760 40109 7788 40140
rect 7745 40103 7803 40109
rect 7745 40069 7757 40103
rect 7791 40069 7803 40103
rect 7745 40063 7803 40069
rect 7837 40103 7895 40109
rect 7837 40069 7849 40103
rect 7883 40100 7895 40103
rect 8018 40100 8024 40112
rect 7883 40072 8024 40100
rect 7883 40069 7895 40072
rect 7837 40063 7895 40069
rect 8018 40060 8024 40072
rect 8076 40060 8082 40112
rect 8202 40060 8208 40112
rect 8260 40060 8266 40112
rect 8496 40100 8524 40140
rect 8573 40137 8585 40171
rect 8619 40168 8631 40171
rect 8619 40140 10272 40168
rect 8619 40137 8631 40140
rect 8573 40131 8631 40137
rect 8496 40072 9076 40100
rect 5213 40004 5672 40032
rect 5213 40001 5225 40004
rect 5167 39995 5225 40001
rect 6454 39992 6460 40044
rect 6512 40032 6518 40044
rect 9048 40032 9076 40072
rect 9122 40060 9128 40112
rect 9180 40060 9186 40112
rect 9306 40100 9312 40112
rect 9232 40072 9312 40100
rect 9232 40032 9260 40072
rect 9306 40060 9312 40072
rect 9364 40100 9370 40112
rect 9401 40103 9459 40109
rect 9401 40100 9413 40103
rect 9364 40072 9413 40100
rect 9364 40060 9370 40072
rect 9401 40069 9413 40072
rect 9447 40069 9459 40103
rect 9401 40063 9459 40069
rect 9493 40103 9551 40109
rect 9493 40069 9505 40103
rect 9539 40100 9551 40103
rect 9766 40100 9772 40112
rect 9539 40072 9772 40100
rect 9539 40069 9551 40072
rect 9493 40063 9551 40069
rect 9766 40060 9772 40072
rect 9824 40060 9830 40112
rect 10244 40109 10272 40140
rect 19610 40128 19616 40180
rect 19668 40128 19674 40180
rect 20901 40171 20959 40177
rect 20901 40137 20913 40171
rect 20947 40137 20959 40171
rect 20901 40131 20959 40137
rect 21177 40171 21235 40177
rect 21177 40137 21189 40171
rect 21223 40137 21235 40171
rect 21177 40131 21235 40137
rect 9861 40103 9919 40109
rect 9861 40069 9873 40103
rect 9907 40069 9919 40103
rect 9861 40063 9919 40069
rect 10229 40103 10287 40109
rect 10229 40069 10241 40103
rect 10275 40100 10287 40103
rect 10318 40100 10324 40112
rect 10275 40072 10324 40100
rect 10275 40069 10287 40072
rect 10229 40063 10287 40069
rect 6512 40004 8800 40032
rect 9048 40004 9260 40032
rect 6512 39992 6518 40004
rect 3292 39936 3372 39964
rect 3292 39924 3298 39936
rect 7926 39924 7932 39976
rect 7984 39924 7990 39976
rect 2866 39856 2872 39908
rect 2924 39896 2930 39908
rect 3970 39896 3976 39908
rect 2924 39868 3976 39896
rect 2924 39856 2930 39868
rect 3970 39856 3976 39868
rect 4028 39856 4034 39908
rect 8772 39905 8800 40004
rect 9674 39992 9680 40044
rect 9732 40032 9738 40044
rect 9876 40032 9904 40063
rect 10318 40060 10324 40072
rect 10376 40060 10382 40112
rect 19245 40103 19303 40109
rect 19245 40069 19257 40103
rect 19291 40100 19303 40103
rect 19628 40100 19656 40128
rect 20916 40100 20944 40131
rect 19291 40072 19656 40100
rect 20272 40072 20944 40100
rect 21192 40100 21220 40131
rect 21818 40128 21824 40180
rect 21876 40128 21882 40180
rect 21910 40128 21916 40180
rect 21968 40128 21974 40180
rect 22186 40128 22192 40180
rect 22244 40168 22250 40180
rect 22244 40140 23428 40168
rect 22244 40128 22250 40140
rect 21928 40100 21956 40128
rect 21192 40072 21956 40100
rect 19291 40069 19303 40072
rect 19245 40063 19303 40069
rect 9732 40004 9904 40032
rect 9732 39992 9738 40004
rect 10778 39992 10784 40044
rect 10836 40032 10842 40044
rect 11057 40035 11115 40041
rect 11057 40032 11069 40035
rect 10836 40004 11069 40032
rect 10836 39992 10842 40004
rect 11057 40001 11069 40004
rect 11103 40001 11115 40035
rect 11057 39995 11115 40001
rect 12710 39992 12716 40044
rect 12768 39992 12774 40044
rect 19978 39992 19984 40044
rect 20036 39992 20042 40044
rect 20272 40041 20300 40072
rect 22646 40060 22652 40112
rect 22704 40100 22710 40112
rect 22704 40072 23152 40100
rect 22704 40060 22710 40072
rect 20257 40035 20315 40041
rect 20257 40001 20269 40035
rect 20303 40001 20315 40035
rect 20257 39995 20315 40001
rect 20533 40035 20591 40041
rect 20533 40001 20545 40035
rect 20579 40032 20591 40035
rect 20714 40032 20720 40044
rect 20579 40004 20720 40032
rect 20579 40001 20591 40004
rect 20533 39995 20591 40001
rect 20714 39992 20720 40004
rect 20772 39992 20778 40044
rect 20809 40035 20867 40041
rect 20809 40001 20821 40035
rect 20855 40032 20867 40035
rect 20898 40032 20904 40044
rect 20855 40004 20904 40032
rect 20855 40001 20867 40004
rect 20809 39995 20867 40001
rect 20898 39992 20904 40004
rect 20956 39992 20962 40044
rect 21085 40035 21143 40041
rect 21085 40001 21097 40035
rect 21131 40032 21143 40035
rect 21266 40032 21272 40044
rect 21131 40004 21272 40032
rect 21131 40001 21143 40004
rect 21085 39995 21143 40001
rect 21266 39992 21272 40004
rect 21324 39992 21330 40044
rect 21358 39992 21364 40044
rect 21416 39992 21422 40044
rect 21634 39992 21640 40044
rect 21692 39992 21698 40044
rect 22002 39992 22008 40044
rect 22060 39992 22066 40044
rect 22186 39992 22192 40044
rect 22244 40032 22250 40044
rect 22281 40035 22339 40041
rect 22281 40032 22293 40035
rect 22244 40004 22293 40032
rect 22244 39992 22250 40004
rect 22281 40001 22293 40004
rect 22327 40001 22339 40035
rect 22281 39995 22339 40001
rect 22557 40035 22615 40041
rect 22557 40001 22569 40035
rect 22603 40001 22615 40035
rect 22557 39995 22615 40001
rect 9582 39924 9588 39976
rect 9640 39924 9646 39976
rect 11238 39924 11244 39976
rect 11296 39964 11302 39976
rect 11793 39967 11851 39973
rect 11793 39964 11805 39967
rect 11296 39936 11805 39964
rect 11296 39924 11302 39936
rect 11793 39933 11805 39936
rect 11839 39933 11851 39967
rect 11793 39927 11851 39933
rect 11977 39967 12035 39973
rect 11977 39933 11989 39967
rect 12023 39933 12035 39967
rect 11977 39927 12035 39933
rect 8757 39899 8815 39905
rect 8757 39865 8769 39899
rect 8803 39865 8815 39899
rect 8757 39859 8815 39865
rect 2314 39788 2320 39840
rect 2372 39828 2378 39840
rect 2961 39831 3019 39837
rect 2961 39828 2973 39831
rect 2372 39800 2973 39828
rect 2372 39788 2378 39800
rect 2961 39797 2973 39800
rect 3007 39797 3019 39831
rect 2961 39791 3019 39797
rect 3510 39788 3516 39840
rect 3568 39828 3574 39840
rect 4065 39831 4123 39837
rect 4065 39828 4077 39831
rect 3568 39800 4077 39828
rect 3568 39788 3574 39800
rect 4065 39797 4077 39800
rect 4111 39797 4123 39831
rect 4065 39791 4123 39797
rect 4614 39788 4620 39840
rect 4672 39788 4678 39840
rect 5902 39788 5908 39840
rect 5960 39788 5966 39840
rect 10410 39788 10416 39840
rect 10468 39788 10474 39840
rect 11790 39788 11796 39840
rect 11848 39828 11854 39840
rect 11992 39828 12020 39927
rect 12342 39924 12348 39976
rect 12400 39964 12406 39976
rect 12437 39967 12495 39973
rect 12437 39964 12449 39967
rect 12400 39936 12449 39964
rect 12400 39924 12406 39936
rect 12437 39933 12449 39936
rect 12483 39933 12495 39967
rect 12830 39967 12888 39973
rect 12830 39964 12842 39967
rect 12437 39927 12495 39933
rect 12544 39936 12842 39964
rect 11848 39800 12020 39828
rect 11848 39788 11854 39800
rect 12158 39788 12164 39840
rect 12216 39828 12222 39840
rect 12544 39828 12572 39936
rect 12830 39933 12842 39936
rect 12876 39933 12888 39967
rect 12830 39927 12888 39933
rect 12989 39967 13047 39973
rect 12989 39933 13001 39967
rect 13035 39964 13047 39967
rect 13354 39964 13360 39976
rect 13035 39936 13360 39964
rect 13035 39933 13047 39936
rect 12989 39927 13047 39933
rect 13354 39924 13360 39936
rect 13412 39924 13418 39976
rect 22572 39964 22600 39995
rect 22738 39992 22744 40044
rect 22796 40032 22802 40044
rect 23124 40041 23152 40072
rect 23400 40041 23428 40140
rect 23842 40128 23848 40180
rect 23900 40128 23906 40180
rect 23860 40100 23888 40128
rect 23492 40072 23888 40100
rect 22833 40035 22891 40041
rect 22833 40032 22845 40035
rect 22796 40004 22845 40032
rect 22796 39992 22802 40004
rect 22833 40001 22845 40004
rect 22879 40001 22891 40035
rect 22833 39995 22891 40001
rect 23109 40035 23167 40041
rect 23109 40001 23121 40035
rect 23155 40001 23167 40035
rect 23109 39995 23167 40001
rect 23385 40035 23443 40041
rect 23385 40001 23397 40035
rect 23431 40001 23443 40035
rect 23385 39995 23443 40001
rect 20364 39936 22600 39964
rect 19426 39856 19432 39908
rect 19484 39856 19490 39908
rect 19794 39856 19800 39908
rect 19852 39856 19858 39908
rect 20070 39856 20076 39908
rect 20128 39856 20134 39908
rect 20364 39905 20392 39936
rect 20349 39899 20407 39905
rect 20349 39865 20361 39899
rect 20395 39865 20407 39899
rect 20349 39859 20407 39865
rect 20625 39899 20683 39905
rect 20625 39865 20637 39899
rect 20671 39896 20683 39899
rect 21818 39896 21824 39908
rect 20671 39868 21824 39896
rect 20671 39865 20683 39868
rect 20625 39859 20683 39865
rect 21818 39856 21824 39868
rect 21876 39856 21882 39908
rect 22649 39899 22707 39905
rect 22649 39896 22661 39899
rect 21928 39868 22661 39896
rect 12216 39800 12572 39828
rect 13633 39831 13691 39837
rect 12216 39788 12222 39800
rect 13633 39797 13645 39831
rect 13679 39828 13691 39831
rect 20898 39828 20904 39840
rect 13679 39800 20904 39828
rect 13679 39797 13691 39800
rect 13633 39791 13691 39797
rect 20898 39788 20904 39800
rect 20956 39788 20962 39840
rect 21266 39788 21272 39840
rect 21324 39828 21330 39840
rect 21453 39831 21511 39837
rect 21453 39828 21465 39831
rect 21324 39800 21465 39828
rect 21324 39788 21330 39800
rect 21453 39797 21465 39800
rect 21499 39797 21511 39831
rect 21453 39791 21511 39797
rect 21726 39788 21732 39840
rect 21784 39828 21790 39840
rect 21928 39828 21956 39868
rect 22649 39865 22661 39868
rect 22695 39865 22707 39899
rect 22649 39859 22707 39865
rect 22830 39856 22836 39908
rect 22888 39856 22894 39908
rect 23201 39899 23259 39905
rect 23201 39865 23213 39899
rect 23247 39896 23259 39899
rect 23492 39896 23520 40072
rect 23750 39992 23756 40044
rect 23808 40032 23814 40044
rect 23845 40035 23903 40041
rect 23845 40032 23857 40035
rect 23808 40004 23857 40032
rect 23808 39992 23814 40004
rect 23845 40001 23857 40004
rect 23891 40001 23903 40035
rect 23845 39995 23903 40001
rect 24118 39992 24124 40044
rect 24176 39992 24182 40044
rect 23247 39868 23520 39896
rect 23247 39865 23259 39868
rect 23201 39859 23259 39865
rect 21784 39800 21956 39828
rect 22097 39831 22155 39837
rect 21784 39788 21790 39800
rect 22097 39797 22109 39831
rect 22143 39828 22155 39831
rect 22278 39828 22284 39840
rect 22143 39800 22284 39828
rect 22143 39797 22155 39800
rect 22097 39791 22155 39797
rect 22278 39788 22284 39800
rect 22336 39788 22342 39840
rect 22373 39831 22431 39837
rect 22373 39797 22385 39831
rect 22419 39828 22431 39831
rect 22848 39828 22876 39856
rect 22419 39800 22876 39828
rect 22419 39797 22431 39800
rect 22373 39791 22431 39797
rect 22922 39788 22928 39840
rect 22980 39788 22986 39840
rect 23661 39831 23719 39837
rect 23661 39797 23673 39831
rect 23707 39828 23719 39831
rect 23934 39828 23940 39840
rect 23707 39800 23940 39828
rect 23707 39797 23719 39800
rect 23661 39791 23719 39797
rect 23934 39788 23940 39800
rect 23992 39788 23998 39840
rect 24394 39788 24400 39840
rect 24452 39788 24458 39840
rect 1104 39738 24840 39760
rect 1104 39686 3917 39738
rect 3969 39686 3981 39738
rect 4033 39686 4045 39738
rect 4097 39686 4109 39738
rect 4161 39686 4173 39738
rect 4225 39686 9851 39738
rect 9903 39686 9915 39738
rect 9967 39686 9979 39738
rect 10031 39686 10043 39738
rect 10095 39686 10107 39738
rect 10159 39686 15785 39738
rect 15837 39686 15849 39738
rect 15901 39686 15913 39738
rect 15965 39686 15977 39738
rect 16029 39686 16041 39738
rect 16093 39686 21719 39738
rect 21771 39686 21783 39738
rect 21835 39686 21847 39738
rect 21899 39686 21911 39738
rect 21963 39686 21975 39738
rect 22027 39686 24840 39738
rect 1104 39664 24840 39686
rect 3142 39584 3148 39636
rect 3200 39624 3206 39636
rect 3421 39627 3479 39633
rect 3421 39624 3433 39627
rect 3200 39596 3433 39624
rect 3200 39584 3206 39596
rect 3421 39593 3433 39596
rect 3467 39593 3479 39627
rect 3421 39587 3479 39593
rect 3510 39584 3516 39636
rect 3568 39584 3574 39636
rect 5902 39584 5908 39636
rect 5960 39584 5966 39636
rect 6730 39584 6736 39636
rect 6788 39624 6794 39636
rect 7742 39624 7748 39636
rect 6788 39596 7748 39624
rect 6788 39584 6794 39596
rect 2682 39448 2688 39500
rect 2740 39448 2746 39500
rect 3528 39488 3556 39584
rect 5920 39556 5948 39584
rect 6089 39559 6147 39565
rect 6089 39556 6101 39559
rect 5920 39528 6101 39556
rect 6089 39525 6101 39528
rect 6135 39525 6147 39559
rect 6089 39519 6147 39525
rect 3436 39460 3556 39488
rect 2225 39423 2283 39429
rect 2225 39389 2237 39423
rect 2271 39420 2283 39423
rect 3436 39420 3464 39460
rect 4798 39448 4804 39500
rect 4856 39448 4862 39500
rect 5258 39448 5264 39500
rect 5316 39488 5322 39500
rect 7392 39497 7420 39596
rect 7742 39584 7748 39596
rect 7800 39584 7806 39636
rect 8386 39584 8392 39636
rect 8444 39584 8450 39636
rect 9766 39584 9772 39636
rect 9824 39624 9830 39636
rect 10505 39627 10563 39633
rect 10505 39624 10517 39627
rect 9824 39596 10517 39624
rect 9824 39584 9830 39596
rect 10505 39593 10517 39596
rect 10551 39593 10563 39627
rect 10505 39587 10563 39593
rect 13354 39584 13360 39636
rect 13412 39584 13418 39636
rect 19978 39584 19984 39636
rect 20036 39584 20042 39636
rect 20717 39627 20775 39633
rect 20717 39593 20729 39627
rect 20763 39624 20775 39627
rect 20990 39624 20996 39636
rect 20763 39596 20996 39624
rect 20763 39593 20775 39596
rect 20717 39587 20775 39593
rect 20990 39584 20996 39596
rect 21048 39584 21054 39636
rect 21082 39584 21088 39636
rect 21140 39624 21146 39636
rect 21545 39627 21603 39633
rect 21545 39624 21557 39627
rect 21140 39596 21557 39624
rect 21140 39584 21146 39596
rect 21545 39593 21557 39596
rect 21591 39593 21603 39627
rect 21545 39587 21603 39593
rect 21821 39627 21879 39633
rect 21821 39593 21833 39627
rect 21867 39624 21879 39627
rect 22278 39624 22284 39636
rect 21867 39596 22284 39624
rect 21867 39593 21879 39596
rect 21821 39587 21879 39593
rect 22278 39584 22284 39596
rect 22336 39584 22342 39636
rect 22373 39627 22431 39633
rect 22373 39593 22385 39627
rect 22419 39624 22431 39627
rect 22554 39624 22560 39636
rect 22419 39596 22560 39624
rect 22419 39593 22431 39596
rect 22373 39587 22431 39593
rect 22554 39584 22560 39596
rect 22612 39584 22618 39636
rect 5445 39491 5503 39497
rect 5445 39488 5457 39491
rect 5316 39460 5457 39488
rect 5316 39448 5322 39460
rect 5445 39457 5457 39460
rect 5491 39457 5503 39491
rect 5445 39451 5503 39457
rect 6365 39491 6423 39497
rect 6365 39457 6377 39491
rect 6411 39488 6423 39491
rect 7377 39491 7435 39497
rect 6411 39460 7328 39488
rect 6411 39457 6423 39460
rect 6365 39451 6423 39457
rect 2271 39392 3464 39420
rect 2271 39389 2283 39392
rect 2225 39383 2283 39389
rect 3510 39380 3516 39432
rect 3568 39420 3574 39432
rect 3605 39423 3663 39429
rect 3605 39420 3617 39423
rect 3568 39392 3617 39420
rect 3568 39380 3574 39392
rect 3605 39389 3617 39392
rect 3651 39389 3663 39423
rect 3605 39383 3663 39389
rect 4341 39423 4399 39429
rect 4341 39389 4353 39423
rect 4387 39420 4399 39423
rect 4522 39420 4528 39432
rect 4387 39392 4528 39420
rect 4387 39389 4399 39392
rect 4341 39383 4399 39389
rect 4522 39380 4528 39392
rect 4580 39380 4586 39432
rect 5276 39420 5304 39448
rect 4632 39392 5304 39420
rect 5629 39423 5687 39429
rect 1486 39312 1492 39364
rect 1544 39312 1550 39364
rect 1670 39312 1676 39364
rect 1728 39312 1734 39364
rect 2314 39312 2320 39364
rect 2372 39312 2378 39364
rect 2590 39312 2596 39364
rect 2648 39352 2654 39364
rect 2685 39355 2743 39361
rect 2685 39352 2697 39355
rect 2648 39324 2697 39352
rect 2648 39312 2654 39324
rect 2685 39321 2697 39324
rect 2731 39321 2743 39355
rect 2685 39315 2743 39321
rect 3252 39324 4200 39352
rect 1946 39244 1952 39296
rect 2004 39244 2010 39296
rect 2958 39244 2964 39296
rect 3016 39284 3022 39296
rect 3252 39293 3280 39324
rect 3053 39287 3111 39293
rect 3053 39284 3065 39287
rect 3016 39256 3065 39284
rect 3016 39244 3022 39256
rect 3053 39253 3065 39256
rect 3099 39253 3111 39287
rect 3053 39247 3111 39253
rect 3237 39287 3295 39293
rect 3237 39253 3249 39287
rect 3283 39253 3295 39287
rect 3237 39247 3295 39253
rect 3970 39244 3976 39296
rect 4028 39244 4034 39296
rect 4172 39284 4200 39324
rect 4246 39312 4252 39364
rect 4304 39352 4310 39364
rect 4632 39352 4660 39392
rect 5629 39389 5641 39423
rect 5675 39389 5687 39423
rect 5629 39383 5687 39389
rect 4304 39324 4660 39352
rect 4304 39312 4310 39324
rect 4706 39312 4712 39364
rect 4764 39352 4770 39364
rect 5644 39352 5672 39383
rect 6454 39380 6460 39432
rect 6512 39429 6518 39432
rect 6512 39423 6540 39429
rect 6528 39389 6540 39423
rect 6512 39383 6540 39389
rect 6512 39380 6518 39383
rect 6638 39380 6644 39432
rect 6696 39380 6702 39432
rect 4764 39324 5672 39352
rect 7300 39352 7328 39460
rect 7377 39457 7389 39491
rect 7423 39457 7435 39491
rect 7377 39451 7435 39457
rect 11606 39448 11612 39500
rect 11664 39488 11670 39500
rect 12345 39491 12403 39497
rect 12345 39488 12357 39491
rect 11664 39460 12357 39488
rect 11664 39448 11670 39460
rect 12345 39457 12357 39460
rect 12391 39457 12403 39491
rect 19996 39488 20024 39584
rect 22097 39559 22155 39565
rect 22097 39525 22109 39559
rect 22143 39525 22155 39559
rect 22097 39519 22155 39525
rect 19996 39460 21496 39488
rect 12345 39451 12403 39457
rect 7558 39380 7564 39432
rect 7616 39420 7622 39432
rect 7651 39423 7709 39429
rect 7651 39420 7663 39423
rect 7616 39392 7663 39420
rect 7616 39380 7622 39392
rect 7651 39389 7663 39392
rect 7697 39389 7709 39423
rect 7651 39383 7709 39389
rect 8570 39380 8576 39432
rect 8628 39420 8634 39432
rect 9398 39420 9404 39432
rect 8628 39392 9404 39420
rect 8628 39380 8634 39392
rect 9398 39380 9404 39392
rect 9456 39420 9462 39432
rect 9493 39423 9551 39429
rect 9493 39420 9505 39423
rect 9456 39392 9505 39420
rect 9456 39380 9462 39392
rect 9493 39389 9505 39392
rect 9539 39389 9551 39423
rect 9766 39420 9772 39432
rect 9727 39392 9772 39420
rect 9493 39383 9551 39389
rect 9766 39380 9772 39392
rect 9824 39420 9830 39432
rect 12587 39423 12645 39429
rect 12587 39420 12599 39423
rect 9824 39392 12599 39420
rect 9824 39380 9830 39392
rect 12587 39389 12599 39392
rect 12633 39389 12645 39423
rect 12587 39383 12645 39389
rect 20898 39380 20904 39432
rect 20956 39380 20962 39432
rect 21082 39380 21088 39432
rect 21140 39380 21146 39432
rect 21266 39380 21272 39432
rect 21324 39380 21330 39432
rect 10410 39352 10416 39364
rect 7300 39324 10416 39352
rect 4764 39312 4770 39324
rect 10410 39312 10416 39324
rect 10468 39352 10474 39364
rect 11698 39352 11704 39364
rect 10468 39324 11704 39352
rect 10468 39312 10474 39324
rect 11698 39312 11704 39324
rect 11756 39352 11762 39364
rect 12250 39352 12256 39364
rect 11756 39324 12256 39352
rect 11756 39312 11762 39324
rect 12250 39312 12256 39324
rect 12308 39312 12314 39364
rect 4522 39284 4528 39296
rect 4172 39256 4528 39284
rect 4522 39244 4528 39256
rect 4580 39244 4586 39296
rect 4982 39244 4988 39296
rect 5040 39284 5046 39296
rect 5077 39287 5135 39293
rect 5077 39284 5089 39287
rect 5040 39256 5089 39284
rect 5040 39244 5046 39256
rect 5077 39253 5089 39256
rect 5123 39253 5135 39287
rect 5077 39247 5135 39253
rect 5166 39244 5172 39296
rect 5224 39284 5230 39296
rect 5261 39287 5319 39293
rect 5261 39284 5273 39287
rect 5224 39256 5273 39284
rect 5224 39244 5230 39256
rect 5261 39253 5273 39256
rect 5307 39253 5319 39287
rect 5261 39247 5319 39253
rect 7282 39244 7288 39296
rect 7340 39244 7346 39296
rect 7558 39244 7564 39296
rect 7616 39284 7622 39296
rect 10502 39284 10508 39296
rect 7616 39256 10508 39284
rect 7616 39244 7622 39256
rect 10502 39244 10508 39256
rect 10560 39244 10566 39296
rect 21100 39293 21128 39380
rect 21085 39287 21143 39293
rect 21085 39253 21097 39287
rect 21131 39253 21143 39287
rect 21468 39284 21496 39460
rect 21726 39380 21732 39432
rect 21784 39380 21790 39432
rect 22002 39380 22008 39432
rect 22060 39380 22066 39432
rect 22112 39420 22140 39519
rect 22112 39392 22232 39420
rect 22204 39352 22232 39392
rect 22278 39380 22284 39432
rect 22336 39380 22342 39432
rect 22554 39380 22560 39432
rect 22612 39380 22618 39432
rect 23017 39423 23075 39429
rect 23017 39389 23029 39423
rect 23063 39389 23075 39423
rect 23017 39383 23075 39389
rect 23032 39352 23060 39383
rect 23382 39380 23388 39432
rect 23440 39380 23446 39432
rect 23842 39380 23848 39432
rect 23900 39380 23906 39432
rect 23934 39380 23940 39432
rect 23992 39380 23998 39432
rect 22204 39324 23060 39352
rect 22833 39287 22891 39293
rect 22833 39284 22845 39287
rect 21468 39256 22845 39284
rect 21085 39247 21143 39253
rect 22833 39253 22845 39256
rect 22879 39253 22891 39287
rect 22833 39247 22891 39253
rect 23106 39244 23112 39296
rect 23164 39284 23170 39296
rect 23201 39287 23259 39293
rect 23201 39284 23213 39287
rect 23164 39256 23213 39284
rect 23164 39244 23170 39256
rect 23201 39253 23213 39256
rect 23247 39253 23259 39287
rect 23201 39247 23259 39253
rect 23661 39287 23719 39293
rect 23661 39253 23673 39287
rect 23707 39284 23719 39287
rect 23934 39284 23940 39296
rect 23707 39256 23940 39284
rect 23707 39253 23719 39256
rect 23661 39247 23719 39253
rect 23934 39244 23940 39256
rect 23992 39244 23998 39296
rect 24121 39287 24179 39293
rect 24121 39253 24133 39287
rect 24167 39284 24179 39287
rect 25222 39284 25228 39296
rect 24167 39256 25228 39284
rect 24167 39253 24179 39256
rect 24121 39247 24179 39253
rect 25222 39244 25228 39256
rect 25280 39244 25286 39296
rect 1104 39194 25000 39216
rect 1104 39142 6884 39194
rect 6936 39142 6948 39194
rect 7000 39142 7012 39194
rect 7064 39142 7076 39194
rect 7128 39142 7140 39194
rect 7192 39142 12818 39194
rect 12870 39142 12882 39194
rect 12934 39142 12946 39194
rect 12998 39142 13010 39194
rect 13062 39142 13074 39194
rect 13126 39142 18752 39194
rect 18804 39142 18816 39194
rect 18868 39142 18880 39194
rect 18932 39142 18944 39194
rect 18996 39142 19008 39194
rect 19060 39142 24686 39194
rect 24738 39142 24750 39194
rect 24802 39142 24814 39194
rect 24866 39142 24878 39194
rect 24930 39142 24942 39194
rect 24994 39142 25000 39194
rect 1104 39120 25000 39142
rect 1486 39040 1492 39092
rect 1544 39040 1550 39092
rect 1946 39040 1952 39092
rect 2004 39080 2010 39092
rect 3970 39080 3976 39092
rect 2004 39052 3976 39080
rect 2004 39040 2010 39052
rect 3970 39040 3976 39052
rect 4028 39040 4034 39092
rect 7282 39040 7288 39092
rect 7340 39040 7346 39092
rect 7374 39040 7380 39092
rect 7432 39080 7438 39092
rect 7650 39080 7656 39092
rect 7432 39052 7656 39080
rect 7432 39040 7438 39052
rect 7650 39040 7656 39052
rect 7708 39040 7714 39092
rect 8846 39040 8852 39092
rect 8904 39080 8910 39092
rect 13446 39080 13452 39092
rect 8904 39052 13452 39080
rect 8904 39040 8910 39052
rect 13446 39040 13452 39052
rect 13504 39040 13510 39092
rect 20441 39083 20499 39089
rect 20441 39049 20453 39083
rect 20487 39049 20499 39083
rect 20441 39043 20499 39049
rect 20717 39083 20775 39089
rect 20717 39049 20729 39083
rect 20763 39080 20775 39083
rect 20898 39080 20904 39092
rect 20763 39052 20904 39080
rect 20763 39049 20775 39052
rect 20717 39043 20775 39049
rect 1504 39012 1532 39040
rect 7300 39012 7328 39040
rect 1504 38984 7328 39012
rect 7742 38972 7748 39024
rect 7800 39012 7806 39024
rect 8478 39012 8484 39024
rect 7800 38984 8484 39012
rect 7800 38972 7806 38984
rect 8478 38972 8484 38984
rect 8536 39012 8542 39024
rect 11606 39012 11612 39024
rect 8536 38984 11612 39012
rect 8536 38972 8542 38984
rect 11606 38972 11612 38984
rect 11664 38972 11670 39024
rect 12526 38972 12532 39024
rect 12584 39012 12590 39024
rect 19978 39012 19984 39024
rect 12584 38984 19984 39012
rect 12584 38972 12590 38984
rect 19978 38972 19984 38984
rect 20036 38972 20042 39024
rect 20456 39012 20484 39043
rect 20898 39040 20904 39052
rect 20956 39040 20962 39092
rect 21266 39040 21272 39092
rect 21324 39040 21330 39092
rect 21358 39040 21364 39092
rect 21416 39080 21422 39092
rect 22002 39080 22008 39092
rect 21416 39052 22008 39080
rect 21416 39040 21422 39052
rect 22002 39040 22008 39052
rect 22060 39040 22066 39092
rect 23385 39083 23443 39089
rect 23385 39049 23397 39083
rect 23431 39049 23443 39083
rect 23385 39043 23443 39049
rect 23661 39083 23719 39089
rect 23661 39049 23673 39083
rect 23707 39080 23719 39083
rect 23842 39080 23848 39092
rect 23707 39052 23848 39080
rect 23707 39049 23719 39052
rect 23661 39043 23719 39049
rect 21284 39012 21312 39040
rect 20456 38984 21312 39012
rect 21450 38972 21456 39024
rect 21508 39012 21514 39024
rect 23400 39012 23428 39043
rect 23842 39040 23848 39052
rect 23900 39040 23906 39092
rect 24121 39015 24179 39021
rect 24121 39012 24133 39015
rect 21508 38984 23060 39012
rect 23400 38984 24133 39012
rect 21508 38972 21514 38984
rect 1947 38947 2005 38953
rect 1947 38913 1959 38947
rect 1993 38944 2005 38947
rect 2866 38944 2872 38956
rect 1993 38916 2872 38944
rect 1993 38913 2005 38916
rect 1947 38907 2005 38913
rect 2866 38904 2872 38916
rect 2924 38904 2930 38956
rect 3050 38904 3056 38956
rect 3108 38904 3114 38956
rect 3418 38904 3424 38956
rect 3476 38944 3482 38956
rect 4065 38947 4123 38953
rect 4065 38944 4077 38947
rect 3476 38916 4077 38944
rect 3476 38904 3482 38916
rect 4065 38913 4077 38916
rect 4111 38913 4123 38947
rect 4617 38947 4675 38953
rect 4617 38944 4629 38947
rect 4065 38907 4123 38913
rect 4172 38916 4629 38944
rect 1673 38879 1731 38885
rect 1673 38845 1685 38879
rect 1719 38845 1731 38879
rect 1673 38839 1731 38845
rect 1688 38808 1716 38839
rect 2682 38836 2688 38888
rect 2740 38836 2746 38888
rect 3786 38836 3792 38888
rect 3844 38836 3850 38888
rect 3878 38836 3884 38888
rect 3936 38876 3942 38888
rect 4172 38876 4200 38916
rect 4617 38913 4629 38916
rect 4663 38913 4675 38947
rect 6730 38944 6736 38956
rect 4617 38907 4675 38913
rect 4816 38916 6736 38944
rect 3936 38848 4200 38876
rect 4341 38879 4399 38885
rect 3936 38836 3942 38848
rect 4341 38845 4353 38879
rect 4387 38876 4399 38879
rect 4816 38876 4844 38916
rect 6730 38904 6736 38916
rect 6788 38904 6794 38956
rect 7374 38904 7380 38956
rect 7432 38944 7438 38956
rect 8355 38947 8413 38953
rect 8355 38944 8367 38947
rect 7432 38916 8367 38944
rect 7432 38904 7438 38916
rect 8355 38913 8367 38916
rect 8401 38944 8413 38947
rect 11759 38947 11817 38953
rect 11759 38944 11771 38947
rect 8401 38916 11771 38944
rect 8401 38913 8413 38916
rect 8355 38907 8413 38913
rect 11759 38913 11771 38916
rect 11805 38913 11817 38947
rect 11759 38907 11817 38913
rect 20622 38904 20628 38956
rect 20680 38904 20686 38956
rect 20901 38947 20959 38953
rect 20901 38913 20913 38947
rect 20947 38913 20959 38947
rect 20901 38907 20959 38913
rect 4387 38848 4844 38876
rect 4893 38879 4951 38885
rect 4387 38845 4399 38848
rect 4341 38839 4399 38845
rect 4893 38845 4905 38879
rect 4939 38876 4951 38879
rect 7926 38876 7932 38888
rect 4939 38848 7932 38876
rect 4939 38845 4951 38848
rect 4893 38839 4951 38845
rect 7926 38836 7932 38848
rect 7984 38836 7990 38888
rect 8113 38879 8171 38885
rect 8113 38845 8125 38879
rect 8159 38845 8171 38879
rect 8113 38839 8171 38845
rect 1688 38780 1808 38808
rect 1780 38752 1808 38780
rect 1762 38700 1768 38752
rect 1820 38700 1826 38752
rect 2700 38749 2728 38836
rect 2958 38768 2964 38820
rect 3016 38808 3022 38820
rect 4982 38808 4988 38820
rect 3016 38780 4988 38808
rect 3016 38768 3022 38780
rect 4982 38768 4988 38780
rect 5040 38768 5046 38820
rect 7742 38768 7748 38820
rect 7800 38808 7806 38820
rect 8128 38808 8156 38839
rect 11514 38836 11520 38888
rect 11572 38836 11578 38888
rect 7800 38780 8156 38808
rect 7800 38768 7806 38780
rect 16666 38768 16672 38820
rect 16724 38808 16730 38820
rect 20916 38808 20944 38907
rect 20990 38904 20996 38956
rect 21048 38944 21054 38956
rect 21637 38947 21695 38953
rect 21637 38944 21649 38947
rect 21048 38916 21649 38944
rect 21048 38904 21054 38916
rect 21637 38913 21649 38916
rect 21683 38944 21695 38947
rect 22077 38947 22135 38953
rect 22077 38944 22089 38947
rect 21683 38916 22089 38944
rect 21683 38913 21695 38916
rect 21637 38907 21695 38913
rect 22077 38913 22089 38916
rect 22123 38913 22135 38947
rect 23032 38944 23060 38984
rect 24121 38981 24133 38984
rect 24167 38981 24179 39015
rect 24121 38975 24179 38981
rect 23032 38916 23520 38944
rect 22077 38907 22135 38913
rect 21542 38836 21548 38888
rect 21600 38876 21606 38888
rect 21821 38879 21879 38885
rect 21821 38876 21833 38879
rect 21600 38848 21833 38876
rect 21600 38836 21606 38848
rect 21821 38845 21833 38848
rect 21867 38845 21879 38879
rect 23492 38876 23520 38916
rect 23566 38904 23572 38956
rect 23624 38904 23630 38956
rect 23658 38904 23664 38956
rect 23716 38944 23722 38956
rect 23845 38947 23903 38953
rect 23845 38944 23857 38947
rect 23716 38916 23857 38944
rect 23716 38904 23722 38916
rect 23845 38913 23857 38916
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 23492 38848 24072 38876
rect 21821 38839 21879 38845
rect 23842 38808 23848 38820
rect 16724 38780 20944 38808
rect 23124 38780 23848 38808
rect 16724 38768 16730 38780
rect 2685 38743 2743 38749
rect 2685 38709 2697 38743
rect 2731 38709 2743 38743
rect 2685 38703 2743 38709
rect 4338 38700 4344 38752
rect 4396 38740 4402 38752
rect 8570 38740 8576 38752
rect 4396 38712 8576 38740
rect 4396 38700 4402 38712
rect 8570 38700 8576 38712
rect 8628 38700 8634 38752
rect 9122 38700 9128 38752
rect 9180 38700 9186 38752
rect 12526 38700 12532 38752
rect 12584 38700 12590 38752
rect 14458 38700 14464 38752
rect 14516 38740 14522 38752
rect 18598 38740 18604 38752
rect 14516 38712 18604 38740
rect 14516 38700 14522 38712
rect 18598 38700 18604 38712
rect 18656 38700 18662 38752
rect 21453 38743 21511 38749
rect 21453 38709 21465 38743
rect 21499 38740 21511 38743
rect 22094 38740 22100 38752
rect 21499 38712 22100 38740
rect 21499 38709 21511 38712
rect 21453 38703 21511 38709
rect 22094 38700 22100 38712
rect 22152 38700 22158 38752
rect 22186 38700 22192 38752
rect 22244 38740 22250 38752
rect 23124 38740 23152 38780
rect 23842 38768 23848 38780
rect 23900 38768 23906 38820
rect 24044 38752 24072 38848
rect 22244 38712 23152 38740
rect 23201 38743 23259 38749
rect 22244 38700 22250 38712
rect 23201 38709 23213 38743
rect 23247 38740 23259 38743
rect 23290 38740 23296 38752
rect 23247 38712 23296 38740
rect 23247 38709 23259 38712
rect 23201 38703 23259 38709
rect 23290 38700 23296 38712
rect 23348 38700 23354 38752
rect 24026 38700 24032 38752
rect 24084 38700 24090 38752
rect 24394 38700 24400 38752
rect 24452 38700 24458 38752
rect 1104 38650 24840 38672
rect 1104 38598 3917 38650
rect 3969 38598 3981 38650
rect 4033 38598 4045 38650
rect 4097 38598 4109 38650
rect 4161 38598 4173 38650
rect 4225 38598 9851 38650
rect 9903 38598 9915 38650
rect 9967 38598 9979 38650
rect 10031 38598 10043 38650
rect 10095 38598 10107 38650
rect 10159 38598 15785 38650
rect 15837 38598 15849 38650
rect 15901 38598 15913 38650
rect 15965 38598 15977 38650
rect 16029 38598 16041 38650
rect 16093 38598 21719 38650
rect 21771 38598 21783 38650
rect 21835 38598 21847 38650
rect 21899 38598 21911 38650
rect 21963 38598 21975 38650
rect 22027 38598 24840 38650
rect 1104 38576 24840 38598
rect 5350 38496 5356 38548
rect 5408 38536 5414 38548
rect 9214 38536 9220 38548
rect 5408 38508 9220 38536
rect 5408 38496 5414 38508
rect 9214 38496 9220 38508
rect 9272 38496 9278 38548
rect 12526 38536 12532 38548
rect 12084 38508 12532 38536
rect 5994 38428 6000 38480
rect 6052 38428 6058 38480
rect 11606 38468 11612 38480
rect 11440 38440 11612 38468
rect 6390 38403 6448 38409
rect 6390 38400 6402 38403
rect 5184 38372 6402 38400
rect 5184 38344 5212 38372
rect 6390 38369 6402 38372
rect 6436 38369 6448 38403
rect 6390 38363 6448 38369
rect 1762 38292 1768 38344
rect 1820 38332 1826 38344
rect 3789 38335 3847 38341
rect 3789 38332 3801 38335
rect 1820 38304 3801 38332
rect 1820 38292 1826 38304
rect 3789 38301 3801 38304
rect 3835 38301 3847 38335
rect 3789 38295 3847 38301
rect 4047 38305 4105 38311
rect 750 38224 756 38276
rect 808 38264 814 38276
rect 1397 38267 1455 38273
rect 1397 38264 1409 38267
rect 808 38236 1409 38264
rect 808 38224 814 38236
rect 1397 38233 1409 38236
rect 1443 38233 1455 38267
rect 1397 38227 1455 38233
rect 2222 38224 2228 38276
rect 2280 38224 2286 38276
rect 2409 38267 2467 38273
rect 2409 38233 2421 38267
rect 2455 38233 2467 38267
rect 2409 38227 2467 38233
rect 1210 38156 1216 38208
rect 1268 38196 1274 38208
rect 2424 38196 2452 38227
rect 2866 38224 2872 38276
rect 2924 38264 2930 38276
rect 3145 38267 3203 38273
rect 3145 38264 3157 38267
rect 2924 38236 3157 38264
rect 2924 38224 2930 38236
rect 3145 38233 3157 38236
rect 3191 38264 3203 38267
rect 3694 38264 3700 38276
rect 3191 38236 3700 38264
rect 3191 38233 3203 38236
rect 3145 38227 3203 38233
rect 3694 38224 3700 38236
rect 3752 38224 3758 38276
rect 1268 38168 2452 38196
rect 3804 38196 3832 38295
rect 4047 38271 4059 38305
rect 4093 38302 4105 38305
rect 4093 38271 4108 38302
rect 5166 38292 5172 38344
rect 5224 38292 5230 38344
rect 5350 38292 5356 38344
rect 5408 38292 5414 38344
rect 5534 38292 5540 38344
rect 5592 38292 5598 38344
rect 6270 38292 6276 38344
rect 6328 38292 6334 38344
rect 6546 38292 6552 38344
rect 6604 38292 6610 38344
rect 8478 38292 8484 38344
rect 8536 38332 8542 38344
rect 8846 38332 8852 38344
rect 8536 38304 8852 38332
rect 8536 38292 8542 38304
rect 8846 38292 8852 38304
rect 8904 38332 8910 38344
rect 9125 38335 9183 38341
rect 9125 38332 9137 38335
rect 8904 38304 9137 38332
rect 8904 38292 8910 38304
rect 9125 38301 9137 38304
rect 9171 38301 9183 38335
rect 9398 38311 9404 38344
rect 9125 38295 9183 38301
rect 9383 38305 9404 38311
rect 9456 38332 9462 38344
rect 11146 38332 11152 38344
rect 4047 38265 4108 38271
rect 4080 38264 4108 38265
rect 5442 38264 5448 38276
rect 4080 38236 5448 38264
rect 5442 38224 5448 38236
rect 5500 38224 5506 38276
rect 9383 38271 9395 38305
rect 9456 38304 11152 38332
rect 9456 38292 9462 38304
rect 11146 38292 11152 38304
rect 11204 38292 11210 38344
rect 11440 38341 11468 38440
rect 11606 38428 11612 38440
rect 11664 38428 11670 38480
rect 12084 38477 12112 38508
rect 12526 38496 12532 38508
rect 12584 38496 12590 38548
rect 13262 38496 13268 38548
rect 13320 38496 13326 38548
rect 19889 38539 19947 38545
rect 19889 38505 19901 38539
rect 19935 38536 19947 38539
rect 20622 38536 20628 38548
rect 19935 38508 20628 38536
rect 19935 38505 19947 38508
rect 19889 38499 19947 38505
rect 20622 38496 20628 38508
rect 20680 38496 20686 38548
rect 21174 38496 21180 38548
rect 21232 38536 21238 38548
rect 22465 38539 22523 38545
rect 22465 38536 22477 38539
rect 21232 38508 22477 38536
rect 21232 38496 21238 38508
rect 22465 38505 22477 38508
rect 22511 38505 22523 38539
rect 22465 38499 22523 38505
rect 23566 38496 23572 38548
rect 23624 38536 23630 38548
rect 23661 38539 23719 38545
rect 23661 38536 23673 38539
rect 23624 38508 23673 38536
rect 23624 38496 23630 38508
rect 23661 38505 23673 38508
rect 23707 38505 23719 38539
rect 23661 38499 23719 38505
rect 23750 38496 23756 38548
rect 23808 38496 23814 38548
rect 12069 38471 12127 38477
rect 12069 38437 12081 38471
rect 12115 38437 12127 38471
rect 12069 38431 12127 38437
rect 23017 38471 23075 38477
rect 23017 38437 23029 38471
rect 23063 38468 23075 38471
rect 23768 38468 23796 38496
rect 23063 38440 23796 38468
rect 23063 38437 23075 38440
rect 23017 38431 23075 38437
rect 11974 38360 11980 38412
rect 12032 38400 12038 38412
rect 12158 38400 12164 38412
rect 12032 38372 12164 38400
rect 12032 38360 12038 38372
rect 12158 38360 12164 38372
rect 12216 38400 12222 38412
rect 12345 38403 12403 38409
rect 12345 38400 12357 38403
rect 12216 38372 12357 38400
rect 12216 38360 12222 38372
rect 12345 38369 12357 38372
rect 12391 38369 12403 38403
rect 12345 38363 12403 38369
rect 20714 38360 20720 38412
rect 20772 38400 20778 38412
rect 23106 38400 23112 38412
rect 20772 38372 23112 38400
rect 20772 38360 20778 38372
rect 23106 38360 23112 38372
rect 23164 38360 23170 38412
rect 11425 38335 11483 38341
rect 11425 38301 11437 38335
rect 11471 38301 11483 38335
rect 11425 38295 11483 38301
rect 11609 38335 11667 38341
rect 11609 38301 11621 38335
rect 11655 38301 11667 38335
rect 11609 38295 11667 38301
rect 9429 38271 9441 38292
rect 9383 38265 9441 38271
rect 4338 38196 4344 38208
rect 3804 38168 4344 38196
rect 1268 38156 1274 38168
rect 4338 38156 4344 38168
rect 4396 38156 4402 38208
rect 4430 38156 4436 38208
rect 4488 38196 4494 38208
rect 4706 38196 4712 38208
rect 4488 38168 4712 38196
rect 4488 38156 4494 38168
rect 4706 38156 4712 38168
rect 4764 38156 4770 38208
rect 4798 38156 4804 38208
rect 4856 38156 4862 38208
rect 4890 38156 4896 38208
rect 4948 38196 4954 38208
rect 7193 38199 7251 38205
rect 7193 38196 7205 38199
rect 4948 38168 7205 38196
rect 4948 38156 4954 38168
rect 7193 38165 7205 38168
rect 7239 38165 7251 38199
rect 7193 38159 7251 38165
rect 10134 38156 10140 38208
rect 10192 38156 10198 38208
rect 11624 38196 11652 38295
rect 12434 38292 12440 38344
rect 12492 38341 12498 38344
rect 12492 38335 12520 38341
rect 12508 38301 12520 38335
rect 12492 38295 12520 38301
rect 12492 38292 12498 38295
rect 12618 38292 12624 38344
rect 12676 38292 12682 38344
rect 20070 38292 20076 38344
rect 20128 38292 20134 38344
rect 22094 38292 22100 38344
rect 22152 38292 22158 38344
rect 22646 38292 22652 38344
rect 22704 38292 22710 38344
rect 22741 38335 22799 38341
rect 22741 38301 22753 38335
rect 22787 38332 22799 38335
rect 22925 38335 22983 38341
rect 22787 38304 22876 38332
rect 22787 38301 22799 38304
rect 22741 38295 22799 38301
rect 22848 38208 22876 38304
rect 22925 38301 22937 38335
rect 22971 38301 22983 38335
rect 22925 38295 22983 38301
rect 22940 38264 22968 38295
rect 23198 38292 23204 38344
rect 23256 38292 23262 38344
rect 23290 38292 23296 38344
rect 23348 38332 23354 38344
rect 23477 38335 23535 38341
rect 23477 38332 23489 38335
rect 23348 38304 23489 38332
rect 23348 38292 23354 38304
rect 23477 38301 23489 38304
rect 23523 38301 23535 38335
rect 23477 38295 23535 38301
rect 23845 38335 23903 38341
rect 23845 38301 23857 38335
rect 23891 38301 23903 38335
rect 23845 38295 23903 38301
rect 22940 38236 23336 38264
rect 11790 38196 11796 38208
rect 11624 38168 11796 38196
rect 11790 38156 11796 38168
rect 11848 38196 11854 38208
rect 12158 38196 12164 38208
rect 11848 38168 12164 38196
rect 11848 38156 11854 38168
rect 12158 38156 12164 38168
rect 12216 38156 12222 38208
rect 22186 38156 22192 38208
rect 22244 38156 22250 38208
rect 22830 38156 22836 38208
rect 22888 38156 22894 38208
rect 22922 38156 22928 38208
rect 22980 38156 22986 38208
rect 23308 38205 23336 38236
rect 23382 38224 23388 38276
rect 23440 38264 23446 38276
rect 23860 38264 23888 38295
rect 23934 38292 23940 38344
rect 23992 38292 23998 38344
rect 23440 38236 23888 38264
rect 23440 38224 23446 38236
rect 23293 38199 23351 38205
rect 23293 38165 23305 38199
rect 23339 38165 23351 38199
rect 23293 38159 23351 38165
rect 24121 38199 24179 38205
rect 24121 38165 24133 38199
rect 24167 38196 24179 38199
rect 25222 38196 25228 38208
rect 24167 38168 25228 38196
rect 24167 38165 24179 38168
rect 24121 38159 24179 38165
rect 25222 38156 25228 38168
rect 25280 38156 25286 38208
rect 1104 38106 25000 38128
rect 1104 38054 6884 38106
rect 6936 38054 6948 38106
rect 7000 38054 7012 38106
rect 7064 38054 7076 38106
rect 7128 38054 7140 38106
rect 7192 38054 12818 38106
rect 12870 38054 12882 38106
rect 12934 38054 12946 38106
rect 12998 38054 13010 38106
rect 13062 38054 13074 38106
rect 13126 38054 18752 38106
rect 18804 38054 18816 38106
rect 18868 38054 18880 38106
rect 18932 38054 18944 38106
rect 18996 38054 19008 38106
rect 19060 38054 24686 38106
rect 24738 38054 24750 38106
rect 24802 38054 24814 38106
rect 24866 38054 24878 38106
rect 24930 38054 24942 38106
rect 24994 38054 25000 38106
rect 1104 38032 25000 38054
rect 4798 37992 4804 38004
rect 3896 37964 4804 37992
rect 3513 37927 3571 37933
rect 3513 37893 3525 37927
rect 3559 37924 3571 37927
rect 3602 37924 3608 37936
rect 3559 37896 3608 37924
rect 3559 37893 3571 37896
rect 3513 37887 3571 37893
rect 3602 37884 3608 37896
rect 3660 37884 3666 37936
rect 3896 37933 3924 37964
rect 4798 37952 4804 37964
rect 4856 37952 4862 38004
rect 4982 37952 4988 38004
rect 5040 37952 5046 38004
rect 6546 37952 6552 38004
rect 6604 37992 6610 38004
rect 7377 37995 7435 38001
rect 7377 37992 7389 37995
rect 6604 37964 7389 37992
rect 6604 37952 6610 37964
rect 7377 37961 7389 37964
rect 7423 37961 7435 37995
rect 10134 37992 10140 38004
rect 7377 37955 7435 37961
rect 9324 37964 10140 37992
rect 3881 37927 3939 37933
rect 3881 37893 3893 37927
rect 3927 37893 3939 37927
rect 3881 37887 3939 37893
rect 4617 37927 4675 37933
rect 4617 37893 4629 37927
rect 4663 37924 4675 37927
rect 4998 37924 5026 37952
rect 4663 37896 5026 37924
rect 5813 37927 5871 37933
rect 4663 37893 4675 37896
rect 4617 37887 4675 37893
rect 4724 37868 4752 37896
rect 5813 37893 5825 37927
rect 5859 37924 5871 37927
rect 8570 37924 8576 37936
rect 5859 37896 8576 37924
rect 5859 37893 5871 37896
rect 5813 37887 5871 37893
rect 8570 37884 8576 37896
rect 8628 37884 8634 37936
rect 8938 37884 8944 37936
rect 8996 37884 9002 37936
rect 9214 37884 9220 37936
rect 9272 37884 9278 37936
rect 9324 37933 9352 37964
rect 10134 37952 10140 37964
rect 10192 37952 10198 38004
rect 12618 37952 12624 38004
rect 12676 37992 12682 38004
rect 13081 37995 13139 38001
rect 13081 37992 13093 37995
rect 12676 37964 13093 37992
rect 12676 37952 12682 37964
rect 13081 37961 13093 37964
rect 13127 37961 13139 37995
rect 13081 37955 13139 37961
rect 14458 37952 14464 38004
rect 14516 37992 14522 38004
rect 22094 37992 22100 38004
rect 14516 37964 22100 37992
rect 14516 37952 14522 37964
rect 22094 37952 22100 37964
rect 22152 37952 22158 38004
rect 22186 37952 22192 38004
rect 22244 37992 22250 38004
rect 22244 37964 22876 37992
rect 22244 37952 22250 37964
rect 9309 37927 9367 37933
rect 9309 37893 9321 37927
rect 9355 37893 9367 37927
rect 10045 37927 10103 37933
rect 9309 37887 9367 37893
rect 9398 37896 9996 37924
rect 1394 37816 1400 37868
rect 1452 37816 1458 37868
rect 2191 37859 2249 37865
rect 2191 37856 2203 37859
rect 1504 37828 2203 37856
rect 1210 37748 1216 37800
rect 1268 37788 1274 37800
rect 1504 37788 1532 37828
rect 2191 37825 2203 37828
rect 2237 37825 2249 37859
rect 2191 37819 2249 37825
rect 3789 37859 3847 37865
rect 3789 37825 3801 37859
rect 3835 37856 3847 37859
rect 4154 37856 4160 37868
rect 3835 37828 4160 37856
rect 3835 37825 3847 37828
rect 3789 37819 3847 37825
rect 4154 37816 4160 37828
rect 4212 37816 4218 37868
rect 4249 37859 4307 37865
rect 4249 37825 4261 37859
rect 4295 37856 4307 37859
rect 4338 37856 4344 37868
rect 4295 37828 4344 37856
rect 4295 37825 4307 37828
rect 4249 37819 4307 37825
rect 4338 37816 4344 37828
rect 4396 37816 4402 37868
rect 4706 37816 4712 37868
rect 4764 37816 4770 37868
rect 4982 37816 4988 37868
rect 5040 37816 5046 37868
rect 5350 37816 5356 37868
rect 5408 37856 5414 37868
rect 5537 37859 5595 37865
rect 5537 37856 5549 37859
rect 5408 37828 5549 37856
rect 5408 37816 5414 37828
rect 5537 37825 5549 37828
rect 5583 37825 5595 37859
rect 5537 37819 5595 37825
rect 5718 37816 5724 37868
rect 5776 37856 5782 37868
rect 5776 37828 6408 37856
rect 5776 37816 5782 37828
rect 6380 37800 6408 37828
rect 6546 37816 6552 37868
rect 6604 37856 6610 37868
rect 6639 37859 6697 37865
rect 6639 37856 6651 37859
rect 6604 37828 6651 37856
rect 6604 37816 6610 37828
rect 6639 37825 6651 37828
rect 6685 37825 6697 37859
rect 6639 37819 6697 37825
rect 6730 37816 6736 37868
rect 6788 37856 6794 37868
rect 9398 37856 9426 37896
rect 6788 37828 9426 37856
rect 6788 37816 6794 37828
rect 9674 37816 9680 37868
rect 9732 37816 9738 37868
rect 9968 37856 9996 37896
rect 10045 37893 10057 37927
rect 10091 37924 10103 37927
rect 10091 37896 10364 37924
rect 10091 37893 10103 37896
rect 10045 37887 10103 37893
rect 10336 37868 10364 37896
rect 11146 37884 11152 37936
rect 11204 37924 11210 37936
rect 22462 37924 22468 37936
rect 11204 37896 12296 37924
rect 11204 37884 11210 37896
rect 9968 37828 10088 37856
rect 1268 37760 1532 37788
rect 1268 37748 1274 37760
rect 1670 37748 1676 37800
rect 1728 37748 1734 37800
rect 1762 37748 1768 37800
rect 1820 37788 1826 37800
rect 1949 37791 2007 37797
rect 1949 37788 1961 37791
rect 1820 37760 1961 37788
rect 1820 37748 1826 37760
rect 1949 37757 1961 37760
rect 1995 37757 2007 37791
rect 5261 37791 5319 37797
rect 1949 37751 2007 37757
rect 2976 37760 3358 37788
rect 2976 37729 3004 37760
rect 5261 37757 5273 37791
rect 5307 37788 5319 37791
rect 6178 37788 6184 37800
rect 5307 37760 6184 37788
rect 5307 37757 5319 37760
rect 5261 37751 5319 37757
rect 6178 37748 6184 37760
rect 6236 37748 6242 37800
rect 6362 37748 6368 37800
rect 6420 37748 6426 37800
rect 7098 37748 7104 37800
rect 7156 37788 7162 37800
rect 7558 37788 7564 37800
rect 7156 37760 7564 37788
rect 7156 37748 7162 37760
rect 7558 37748 7564 37760
rect 7616 37748 7622 37800
rect 9122 37748 9128 37800
rect 9180 37748 9186 37800
rect 10060 37788 10088 37828
rect 10318 37816 10324 37868
rect 10376 37816 10382 37868
rect 12268 37856 12296 37896
rect 22112 37896 22468 37924
rect 12343 37859 12401 37865
rect 12343 37856 12355 37859
rect 12268 37828 12355 37856
rect 12343 37825 12355 37828
rect 12389 37856 12401 37859
rect 13538 37856 13544 37868
rect 12389 37828 13544 37856
rect 12389 37825 12401 37828
rect 12343 37819 12401 37825
rect 13538 37816 13544 37828
rect 13596 37816 13602 37868
rect 15470 37816 15476 37868
rect 15528 37856 15534 37868
rect 22112 37865 22140 37896
rect 22462 37884 22468 37896
rect 22520 37884 22526 37936
rect 21637 37859 21695 37865
rect 21637 37856 21649 37859
rect 15528 37828 21649 37856
rect 15528 37816 15534 37828
rect 21637 37825 21649 37828
rect 21683 37825 21695 37859
rect 21637 37819 21695 37825
rect 22095 37859 22153 37865
rect 22095 37825 22107 37859
rect 22141 37825 22153 37859
rect 22848 37856 22876 37964
rect 22922 37952 22928 38004
rect 22980 37952 22986 38004
rect 23106 37952 23112 38004
rect 23164 37992 23170 38004
rect 23845 37995 23903 38001
rect 23845 37992 23857 37995
rect 23164 37964 23857 37992
rect 23164 37952 23170 37964
rect 23845 37961 23857 37964
rect 23891 37961 23903 37995
rect 23845 37955 23903 37961
rect 22940 37924 22968 37952
rect 23753 37927 23811 37933
rect 23753 37924 23765 37927
rect 22940 37896 23765 37924
rect 23753 37893 23765 37896
rect 23799 37893 23811 37927
rect 23753 37887 23811 37893
rect 23385 37859 23443 37865
rect 23385 37856 23397 37859
rect 22848 37828 23397 37856
rect 22095 37819 22153 37825
rect 23385 37825 23397 37828
rect 23431 37825 23443 37859
rect 23385 37819 23443 37825
rect 24026 37816 24032 37868
rect 24084 37816 24090 37868
rect 24213 37859 24271 37865
rect 24213 37825 24225 37859
rect 24259 37825 24271 37859
rect 24213 37819 24271 37825
rect 12069 37791 12127 37797
rect 10060 37760 10824 37788
rect 2961 37723 3019 37729
rect 2961 37689 2973 37723
rect 3007 37689 3019 37723
rect 2961 37683 3019 37689
rect 4801 37723 4859 37729
rect 4801 37689 4813 37723
rect 4847 37720 4859 37723
rect 6270 37720 6276 37732
rect 4847 37692 6276 37720
rect 4847 37689 4859 37692
rect 4801 37683 4859 37689
rect 6012 37664 6040 37692
rect 6270 37680 6276 37692
rect 6328 37680 6334 37732
rect 5994 37612 6000 37664
rect 6052 37612 6058 37664
rect 10229 37655 10287 37661
rect 10229 37621 10241 37655
rect 10275 37652 10287 37655
rect 10594 37652 10600 37664
rect 10275 37624 10600 37652
rect 10275 37621 10287 37624
rect 10229 37615 10287 37621
rect 10594 37612 10600 37624
rect 10652 37612 10658 37664
rect 10796 37652 10824 37760
rect 12069 37757 12081 37791
rect 12115 37757 12127 37791
rect 12069 37751 12127 37757
rect 11514 37680 11520 37732
rect 11572 37720 11578 37732
rect 12084 37720 12112 37751
rect 19518 37748 19524 37800
rect 19576 37788 19582 37800
rect 21821 37791 21879 37797
rect 21821 37788 21833 37791
rect 19576 37760 21833 37788
rect 19576 37748 19582 37760
rect 21821 37757 21833 37760
rect 21867 37757 21879 37791
rect 21821 37751 21879 37757
rect 23201 37791 23259 37797
rect 23201 37757 23213 37791
rect 23247 37757 23259 37791
rect 24228 37788 24256 37819
rect 23201 37751 23259 37757
rect 23308 37760 24256 37788
rect 11572 37692 12112 37720
rect 11572 37680 11578 37692
rect 10962 37652 10968 37664
rect 10796 37624 10968 37652
rect 10962 37612 10968 37624
rect 11020 37652 11026 37664
rect 11790 37652 11796 37664
rect 11020 37624 11796 37652
rect 11020 37612 11026 37624
rect 11790 37612 11796 37624
rect 11848 37612 11854 37664
rect 12084 37652 12112 37692
rect 20162 37680 20168 37732
rect 20220 37720 20226 37732
rect 21453 37723 21511 37729
rect 21453 37720 21465 37723
rect 20220 37692 21465 37720
rect 20220 37680 20226 37692
rect 21453 37689 21465 37692
rect 21499 37689 21511 37723
rect 21453 37683 21511 37689
rect 13906 37652 13912 37664
rect 12084 37624 13912 37652
rect 13906 37612 13912 37624
rect 13964 37612 13970 37664
rect 21836 37652 21864 37751
rect 22830 37680 22836 37732
rect 22888 37720 22894 37732
rect 23216 37720 23244 37751
rect 22888 37692 23244 37720
rect 22888 37680 22894 37692
rect 22554 37652 22560 37664
rect 21836 37624 22560 37652
rect 22554 37612 22560 37624
rect 22612 37612 22618 37664
rect 22922 37612 22928 37664
rect 22980 37652 22986 37664
rect 23308 37652 23336 37760
rect 23661 37723 23719 37729
rect 23661 37689 23673 37723
rect 23707 37720 23719 37723
rect 23707 37692 25084 37720
rect 23707 37689 23719 37692
rect 23661 37683 23719 37689
rect 25056 37664 25084 37692
rect 22980 37624 23336 37652
rect 22980 37612 22986 37624
rect 24394 37612 24400 37664
rect 24452 37612 24458 37664
rect 25038 37612 25044 37664
rect 25096 37612 25102 37664
rect 1104 37562 24840 37584
rect 1104 37510 3917 37562
rect 3969 37510 3981 37562
rect 4033 37510 4045 37562
rect 4097 37510 4109 37562
rect 4161 37510 4173 37562
rect 4225 37510 9851 37562
rect 9903 37510 9915 37562
rect 9967 37510 9979 37562
rect 10031 37510 10043 37562
rect 10095 37510 10107 37562
rect 10159 37510 15785 37562
rect 15837 37510 15849 37562
rect 15901 37510 15913 37562
rect 15965 37510 15977 37562
rect 16029 37510 16041 37562
rect 16093 37510 21719 37562
rect 21771 37510 21783 37562
rect 21835 37510 21847 37562
rect 21899 37510 21911 37562
rect 21963 37510 21975 37562
rect 22027 37510 24840 37562
rect 1104 37488 24840 37510
rect 3418 37408 3424 37460
rect 3476 37408 3482 37460
rect 3878 37408 3884 37460
rect 3936 37448 3942 37460
rect 4982 37448 4988 37460
rect 3936 37420 4988 37448
rect 3936 37408 3942 37420
rect 4982 37408 4988 37420
rect 5040 37408 5046 37460
rect 6178 37408 6184 37460
rect 6236 37448 6242 37460
rect 6236 37420 7420 37448
rect 6236 37408 6242 37420
rect 7392 37380 7420 37420
rect 7466 37408 7472 37460
rect 7524 37448 7530 37460
rect 7524 37420 10732 37448
rect 7524 37408 7530 37420
rect 7558 37380 7564 37392
rect 7392 37352 7564 37380
rect 7558 37340 7564 37352
rect 7616 37380 7622 37392
rect 7616 37352 8616 37380
rect 7616 37340 7622 37352
rect 842 37272 848 37324
rect 900 37312 906 37324
rect 2130 37312 2136 37324
rect 900 37284 2136 37312
rect 900 37272 906 37284
rect 2130 37272 2136 37284
rect 2188 37272 2194 37324
rect 2424 37284 3004 37312
rect 1026 37204 1032 37256
rect 1084 37244 1090 37256
rect 2424 37244 2452 37284
rect 1084 37216 2452 37244
rect 2501 37247 2559 37253
rect 1084 37204 1090 37216
rect 2501 37213 2513 37247
rect 2547 37244 2559 37247
rect 2976 37244 3004 37284
rect 3418 37272 3424 37324
rect 3476 37312 3482 37324
rect 3476 37284 4384 37312
rect 3476 37272 3482 37284
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 2547 37216 2912 37244
rect 2976 37216 3801 37244
rect 2547 37213 2559 37216
rect 2501 37207 2559 37213
rect 2884 37188 2912 37216
rect 3789 37213 3801 37216
rect 3835 37213 3847 37247
rect 3789 37207 3847 37213
rect 1397 37179 1455 37185
rect 1397 37145 1409 37179
rect 1443 37176 1455 37179
rect 1486 37176 1492 37188
rect 1443 37148 1492 37176
rect 1443 37145 1455 37148
rect 1397 37139 1455 37145
rect 1486 37136 1492 37148
rect 1544 37136 1550 37188
rect 2222 37136 2228 37188
rect 2280 37136 2286 37188
rect 2774 37136 2780 37188
rect 2832 37136 2838 37188
rect 2866 37136 2872 37188
rect 2924 37136 2930 37188
rect 3145 37179 3203 37185
rect 3145 37145 3157 37179
rect 3191 37145 3203 37179
rect 3145 37139 3203 37145
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 3160 37108 3188 37139
rect 4062 37136 4068 37188
rect 4120 37136 4126 37188
rect 4356 37176 4384 37284
rect 7282 37272 7288 37324
rect 7340 37312 7346 37324
rect 8205 37315 8263 37321
rect 7340 37284 8064 37312
rect 7340 37272 7346 37284
rect 4709 37247 4767 37253
rect 4709 37213 4721 37247
rect 4755 37244 4767 37247
rect 4755 37216 4936 37244
rect 4755 37213 4767 37216
rect 4709 37207 4767 37213
rect 4798 37176 4804 37188
rect 4356 37148 4804 37176
rect 4798 37136 4804 37148
rect 4856 37136 4862 37188
rect 4908 37176 4936 37216
rect 4982 37204 4988 37256
rect 5040 37244 5046 37256
rect 5442 37244 5448 37256
rect 5040 37216 5448 37244
rect 5040 37204 5046 37216
rect 5442 37204 5448 37216
rect 5500 37204 5506 37256
rect 8036 37253 8064 37284
rect 8205 37281 8217 37315
rect 8251 37312 8263 37315
rect 8389 37315 8447 37321
rect 8389 37312 8401 37315
rect 8251 37284 8401 37312
rect 8251 37281 8263 37284
rect 8205 37275 8263 37281
rect 8389 37281 8401 37284
rect 8435 37281 8447 37315
rect 8389 37275 8447 37281
rect 6549 37247 6607 37253
rect 6549 37213 6561 37247
rect 6595 37213 6607 37247
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 6549 37207 6607 37213
rect 6807 37217 6865 37223
rect 5534 37176 5540 37188
rect 4908 37148 5540 37176
rect 5534 37136 5540 37148
rect 5592 37176 5598 37188
rect 6564 37176 6592 37207
rect 6807 37183 6819 37217
rect 6853 37214 6865 37217
rect 7576 37216 7941 37244
rect 6853 37183 6868 37214
rect 6807 37177 6868 37183
rect 5592 37148 6592 37176
rect 5592 37136 5598 37148
rect 1360 37080 3188 37108
rect 1360 37068 1366 37080
rect 3694 37068 3700 37120
rect 3752 37108 3758 37120
rect 4890 37108 4896 37120
rect 3752 37080 4896 37108
rect 3752 37068 3758 37080
rect 4890 37068 4896 37080
rect 4948 37068 4954 37120
rect 5718 37068 5724 37120
rect 5776 37068 5782 37120
rect 6730 37068 6736 37120
rect 6788 37108 6794 37120
rect 6840 37108 6868 37177
rect 7576 37117 7604 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 7929 37207 7987 37213
rect 8021 37247 8079 37253
rect 8021 37213 8033 37247
rect 8067 37213 8079 37247
rect 8021 37207 8079 37213
rect 8297 37247 8355 37253
rect 8297 37213 8309 37247
rect 8343 37213 8355 37247
rect 8297 37207 8355 37213
rect 7944 37176 7972 37207
rect 8312 37176 8340 37207
rect 8478 37204 8484 37256
rect 8536 37204 8542 37256
rect 7944 37148 8340 37176
rect 8588 37176 8616 37352
rect 10042 37272 10048 37324
rect 10100 37272 10106 37324
rect 10704 37312 10732 37420
rect 20070 37408 20076 37460
rect 20128 37408 20134 37460
rect 22557 37451 22615 37457
rect 22557 37417 22569 37451
rect 22603 37448 22615 37451
rect 22646 37448 22652 37460
rect 22603 37420 22652 37448
rect 22603 37417 22615 37420
rect 22557 37411 22615 37417
rect 22646 37408 22652 37420
rect 22704 37408 22710 37460
rect 22833 37451 22891 37457
rect 22833 37417 22845 37451
rect 22879 37448 22891 37451
rect 23382 37448 23388 37460
rect 22879 37420 23388 37448
rect 22879 37417 22891 37420
rect 22833 37411 22891 37417
rect 23382 37408 23388 37420
rect 23440 37408 23446 37460
rect 11790 37340 11796 37392
rect 11848 37380 11854 37392
rect 20088 37380 20116 37408
rect 11848 37352 20116 37380
rect 21913 37383 21971 37389
rect 11848 37340 11854 37352
rect 21913 37349 21925 37383
rect 21959 37380 21971 37383
rect 23198 37380 23204 37392
rect 21959 37352 23204 37380
rect 21959 37349 21971 37352
rect 21913 37343 21971 37349
rect 23198 37340 23204 37352
rect 23256 37340 23262 37392
rect 13722 37312 13728 37324
rect 10704 37284 13728 37312
rect 13722 37272 13728 37284
rect 13780 37272 13786 37324
rect 20456 37284 20852 37312
rect 8662 37204 8668 37256
rect 8720 37244 8726 37256
rect 10319 37247 10377 37253
rect 10319 37244 10331 37247
rect 8720 37216 10331 37244
rect 8720 37204 8726 37216
rect 10319 37213 10331 37216
rect 10365 37244 10377 37247
rect 20254 37244 20260 37256
rect 10365 37216 20260 37244
rect 10365 37213 10377 37216
rect 10319 37207 10377 37213
rect 20254 37204 20260 37216
rect 20312 37204 20318 37256
rect 20456 37176 20484 37284
rect 20530 37204 20536 37256
rect 20588 37204 20594 37256
rect 20714 37204 20720 37256
rect 20772 37204 20778 37256
rect 20824 37244 20852 37284
rect 21744 37284 22232 37312
rect 21744 37244 21772 37284
rect 20824 37216 21772 37244
rect 21818 37204 21824 37256
rect 21876 37204 21882 37256
rect 22097 37247 22155 37253
rect 22097 37213 22109 37247
rect 22143 37213 22155 37247
rect 22097 37207 22155 37213
rect 8588 37148 20484 37176
rect 6788 37080 6868 37108
rect 7561 37111 7619 37117
rect 6788 37068 6794 37080
rect 7561 37077 7573 37111
rect 7607 37077 7619 37111
rect 7561 37071 7619 37077
rect 8110 37068 8116 37120
rect 8168 37108 8174 37120
rect 8205 37111 8263 37117
rect 8205 37108 8217 37111
rect 8168 37080 8217 37108
rect 8168 37068 8174 37080
rect 8205 37077 8217 37080
rect 8251 37077 8263 37111
rect 8205 37071 8263 37077
rect 11054 37068 11060 37120
rect 11112 37068 11118 37120
rect 20548 37117 20576 37204
rect 21910 37136 21916 37188
rect 21968 37176 21974 37188
rect 22112 37176 22140 37207
rect 22204 37188 22232 37284
rect 24118 37272 24124 37324
rect 24176 37272 24182 37324
rect 22738 37204 22744 37256
rect 22796 37204 22802 37256
rect 23017 37247 23075 37253
rect 23017 37213 23029 37247
rect 23063 37213 23075 37247
rect 23017 37207 23075 37213
rect 21968 37148 22140 37176
rect 21968 37136 21974 37148
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 23032 37176 23060 37207
rect 23106 37204 23112 37256
rect 23164 37244 23170 37256
rect 23293 37247 23351 37253
rect 23293 37244 23305 37247
rect 23164 37216 23305 37244
rect 23164 37204 23170 37216
rect 23293 37213 23305 37216
rect 23339 37213 23351 37247
rect 23293 37207 23351 37213
rect 23566 37204 23572 37256
rect 23624 37204 23630 37256
rect 23658 37204 23664 37256
rect 23716 37204 23722 37256
rect 24210 37204 24216 37256
rect 24268 37204 24274 37256
rect 23676 37176 23704 37204
rect 22244 37148 23060 37176
rect 23124 37148 23704 37176
rect 22244 37136 22250 37148
rect 20533 37111 20591 37117
rect 20533 37077 20545 37111
rect 20579 37077 20591 37111
rect 20533 37071 20591 37077
rect 21637 37111 21695 37117
rect 21637 37077 21649 37111
rect 21683 37108 21695 37111
rect 22922 37108 22928 37120
rect 21683 37080 22928 37108
rect 21683 37077 21695 37080
rect 21637 37071 21695 37077
rect 22922 37068 22928 37080
rect 22980 37068 22986 37120
rect 23124 37117 23152 37148
rect 23842 37136 23848 37188
rect 23900 37136 23906 37188
rect 23109 37111 23167 37117
rect 23109 37077 23121 37111
rect 23155 37077 23167 37111
rect 23109 37071 23167 37077
rect 23385 37111 23443 37117
rect 23385 37077 23397 37111
rect 23431 37108 23443 37111
rect 24228 37108 24256 37204
rect 23431 37080 24256 37108
rect 23431 37077 23443 37080
rect 23385 37071 23443 37077
rect 1104 37018 25000 37040
rect 1104 36966 6884 37018
rect 6936 36966 6948 37018
rect 7000 36966 7012 37018
rect 7064 36966 7076 37018
rect 7128 36966 7140 37018
rect 7192 36966 12818 37018
rect 12870 36966 12882 37018
rect 12934 36966 12946 37018
rect 12998 36966 13010 37018
rect 13062 36966 13074 37018
rect 13126 36966 18752 37018
rect 18804 36966 18816 37018
rect 18868 36966 18880 37018
rect 18932 36966 18944 37018
rect 18996 36966 19008 37018
rect 19060 36966 24686 37018
rect 24738 36966 24750 37018
rect 24802 36966 24814 37018
rect 24866 36966 24878 37018
rect 24930 36966 24942 37018
rect 24994 36966 25000 37018
rect 1104 36944 25000 36966
rect 474 36864 480 36916
rect 532 36864 538 36916
rect 3694 36904 3700 36916
rect 1596 36876 3700 36904
rect 492 36712 520 36864
rect 1596 36845 1624 36876
rect 3694 36864 3700 36876
rect 3752 36864 3758 36916
rect 5905 36907 5963 36913
rect 5905 36904 5917 36907
rect 3804 36876 5917 36904
rect 1581 36839 1639 36845
rect 1581 36805 1593 36839
rect 1627 36805 1639 36839
rect 1581 36799 1639 36805
rect 3418 36796 3424 36848
rect 3476 36836 3482 36848
rect 3602 36836 3608 36848
rect 3476 36808 3608 36836
rect 3476 36796 3482 36808
rect 3602 36796 3608 36808
rect 3660 36796 3666 36848
rect 3804 36845 3832 36876
rect 5905 36873 5917 36876
rect 5951 36873 5963 36907
rect 5905 36867 5963 36873
rect 7193 36907 7251 36913
rect 7193 36873 7205 36907
rect 7239 36873 7251 36907
rect 7193 36867 7251 36873
rect 3789 36839 3847 36845
rect 3789 36805 3801 36839
rect 3835 36805 3847 36839
rect 4246 36836 4252 36848
rect 3789 36799 3847 36805
rect 3988 36808 4252 36836
rect 2131 36771 2189 36777
rect 2131 36737 2143 36771
rect 2177 36768 2189 36771
rect 2774 36768 2780 36780
rect 2177 36740 2780 36768
rect 2177 36737 2189 36740
rect 2131 36731 2189 36737
rect 2774 36728 2780 36740
rect 2832 36728 2838 36780
rect 3697 36771 3755 36777
rect 3697 36737 3709 36771
rect 3743 36768 3755 36771
rect 3988 36768 4016 36808
rect 4246 36796 4252 36808
rect 4304 36796 4310 36848
rect 4525 36839 4583 36845
rect 4525 36805 4537 36839
rect 4571 36836 4583 36839
rect 4571 36808 4752 36836
rect 4571 36805 4583 36808
rect 4525 36799 4583 36805
rect 4724 36780 4752 36808
rect 4798 36796 4804 36848
rect 4856 36836 4862 36848
rect 5810 36836 5816 36848
rect 4856 36808 5816 36836
rect 4856 36796 4862 36808
rect 3743 36740 4016 36768
rect 4157 36771 4215 36777
rect 3743 36737 3755 36740
rect 3697 36731 3755 36737
rect 4157 36737 4169 36771
rect 4203 36768 4215 36771
rect 4338 36768 4344 36780
rect 4203 36740 4344 36768
rect 4203 36737 4215 36740
rect 4157 36731 4215 36737
rect 4338 36728 4344 36740
rect 4396 36768 4402 36780
rect 4614 36768 4620 36780
rect 4396 36740 4620 36768
rect 4396 36728 4402 36740
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 4706 36728 4712 36780
rect 4764 36728 4770 36780
rect 5166 36777 5194 36808
rect 5810 36796 5816 36808
rect 5868 36796 5874 36848
rect 7208 36836 7236 36867
rect 8478 36864 8484 36916
rect 8536 36864 8542 36916
rect 8570 36864 8576 36916
rect 8628 36904 8634 36916
rect 20349 36907 20407 36913
rect 8628 36876 17264 36904
rect 8628 36864 8634 36876
rect 8496 36836 8524 36864
rect 17236 36836 17264 36876
rect 20349 36873 20361 36907
rect 20395 36904 20407 36907
rect 20714 36904 20720 36916
rect 20395 36876 20720 36904
rect 20395 36873 20407 36876
rect 20349 36867 20407 36873
rect 20714 36864 20720 36876
rect 20772 36864 20778 36916
rect 20901 36907 20959 36913
rect 20901 36873 20913 36907
rect 20947 36904 20959 36907
rect 21818 36904 21824 36916
rect 20947 36876 21824 36904
rect 20947 36873 20959 36876
rect 20901 36867 20959 36873
rect 21818 36864 21824 36876
rect 21876 36864 21882 36916
rect 21910 36864 21916 36916
rect 21968 36864 21974 36916
rect 23842 36904 23848 36916
rect 22066 36876 23848 36904
rect 21928 36836 21956 36864
rect 7208 36808 8524 36836
rect 12406 36808 17172 36836
rect 17236 36808 21956 36836
rect 5151 36771 5209 36777
rect 5151 36737 5163 36771
rect 5197 36737 5209 36771
rect 5151 36731 5209 36737
rect 6914 36728 6920 36780
rect 6972 36728 6978 36780
rect 7009 36771 7067 36777
rect 7009 36737 7021 36771
rect 7055 36768 7067 36771
rect 7282 36768 7288 36780
rect 7055 36740 7288 36768
rect 7055 36737 7067 36740
rect 7009 36731 7067 36737
rect 7282 36728 7288 36740
rect 7340 36728 7346 36780
rect 7374 36728 7380 36780
rect 7432 36728 7438 36780
rect 7650 36728 7656 36780
rect 7708 36768 7714 36780
rect 7743 36771 7801 36777
rect 7743 36768 7755 36771
rect 7708 36740 7755 36768
rect 7708 36728 7714 36740
rect 7743 36737 7755 36740
rect 7789 36768 7801 36771
rect 7789 36740 8156 36768
rect 7789 36737 7801 36740
rect 7743 36731 7801 36737
rect 474 36660 480 36712
rect 532 36660 538 36712
rect 1857 36703 1915 36709
rect 1857 36669 1869 36703
rect 1903 36669 1915 36703
rect 1857 36663 1915 36669
rect 934 36524 940 36576
rect 992 36564 998 36576
rect 1673 36567 1731 36573
rect 1673 36564 1685 36567
rect 992 36536 1685 36564
rect 992 36524 998 36536
rect 1673 36533 1685 36536
rect 1719 36533 1731 36567
rect 1872 36564 1900 36663
rect 2869 36635 2927 36641
rect 2869 36601 2881 36635
rect 2915 36632 2927 36635
rect 3252 36632 3280 36686
rect 4890 36660 4896 36712
rect 4948 36660 4954 36712
rect 7469 36703 7527 36709
rect 7469 36700 7481 36703
rect 7300 36672 7481 36700
rect 7300 36644 7328 36672
rect 7469 36669 7481 36672
rect 7515 36669 7527 36703
rect 8128 36700 8156 36740
rect 9122 36728 9128 36780
rect 9180 36768 9186 36780
rect 11759 36771 11817 36777
rect 11759 36768 11771 36771
rect 9180 36740 11771 36768
rect 9180 36728 9186 36740
rect 11759 36737 11771 36740
rect 11805 36768 11817 36771
rect 12406 36768 12434 36808
rect 11805 36740 12434 36768
rect 11805 36737 11817 36740
rect 11759 36731 11817 36737
rect 16666 36728 16672 36780
rect 16724 36728 16730 36780
rect 8478 36700 8484 36712
rect 8128 36672 8484 36700
rect 7469 36663 7527 36669
rect 8478 36660 8484 36672
rect 8536 36700 8542 36712
rect 8662 36700 8668 36712
rect 8536 36672 8668 36700
rect 8536 36660 8542 36672
rect 8662 36660 8668 36672
rect 8720 36660 8726 36712
rect 10042 36660 10048 36712
rect 10100 36700 10106 36712
rect 10410 36700 10416 36712
rect 10100 36672 10416 36700
rect 10100 36660 10106 36672
rect 10410 36660 10416 36672
rect 10468 36700 10474 36712
rect 11517 36703 11575 36709
rect 11517 36700 11529 36703
rect 10468 36672 11529 36700
rect 10468 36660 10474 36672
rect 11517 36669 11529 36672
rect 11563 36669 11575 36703
rect 11517 36663 11575 36669
rect 2915 36604 3280 36632
rect 2915 36601 2927 36604
rect 2869 36595 2927 36601
rect 7282 36592 7288 36644
rect 7340 36592 7346 36644
rect 9766 36632 9772 36644
rect 8312 36604 9772 36632
rect 2314 36564 2320 36576
rect 1872 36536 2320 36564
rect 1673 36527 1731 36533
rect 2314 36524 2320 36536
rect 2372 36524 2378 36576
rect 4709 36567 4767 36573
rect 4709 36533 4721 36567
rect 4755 36564 4767 36567
rect 5626 36564 5632 36576
rect 4755 36536 5632 36564
rect 4755 36533 4767 36536
rect 4709 36527 4767 36533
rect 5626 36524 5632 36536
rect 5684 36524 5690 36576
rect 6730 36524 6736 36576
rect 6788 36564 6794 36576
rect 8312 36564 8340 36604
rect 9766 36592 9772 36604
rect 9824 36632 9830 36644
rect 10778 36632 10784 36644
rect 9824 36604 10784 36632
rect 9824 36592 9830 36604
rect 10778 36592 10784 36604
rect 10836 36592 10842 36644
rect 11532 36632 11560 36663
rect 16684 36632 16712 36728
rect 11532 36604 11585 36632
rect 6788 36536 8340 36564
rect 6788 36524 6794 36536
rect 8386 36524 8392 36576
rect 8444 36564 8450 36576
rect 8481 36567 8539 36573
rect 8481 36564 8493 36567
rect 8444 36536 8493 36564
rect 8444 36524 8450 36536
rect 8481 36533 8493 36536
rect 8527 36533 8539 36567
rect 11557 36564 11585 36604
rect 12176 36604 16712 36632
rect 12176 36564 12204 36604
rect 17144 36576 17172 36808
rect 17773 36771 17831 36777
rect 17773 36768 17785 36771
rect 17420 36740 17785 36768
rect 17420 36576 17448 36740
rect 17773 36737 17785 36740
rect 17819 36737 17831 36771
rect 17773 36731 17831 36737
rect 19153 36771 19211 36777
rect 19153 36737 19165 36771
rect 19199 36768 19211 36771
rect 19242 36768 19248 36780
rect 19199 36740 19248 36768
rect 19199 36737 19211 36740
rect 19153 36731 19211 36737
rect 19242 36728 19248 36740
rect 19300 36728 19306 36780
rect 19797 36771 19855 36777
rect 19797 36737 19809 36771
rect 19843 36737 19855 36771
rect 19797 36731 19855 36737
rect 19812 36700 19840 36731
rect 20254 36728 20260 36780
rect 20312 36728 20318 36780
rect 20530 36728 20536 36780
rect 20588 36728 20594 36780
rect 20714 36728 20720 36780
rect 20772 36768 20778 36780
rect 20809 36771 20867 36777
rect 20809 36768 20821 36771
rect 20772 36740 20821 36768
rect 20772 36728 20778 36740
rect 20809 36737 20821 36740
rect 20855 36737 20867 36771
rect 20809 36731 20867 36737
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36737 21143 36771
rect 21085 36731 21143 36737
rect 21100 36700 21128 36731
rect 18984 36672 19840 36700
rect 20088 36672 21128 36700
rect 18984 36641 19012 36672
rect 20088 36641 20116 36672
rect 18969 36635 19027 36641
rect 18969 36601 18981 36635
rect 19015 36601 19027 36635
rect 18969 36595 19027 36601
rect 20073 36635 20131 36641
rect 20073 36601 20085 36635
rect 20119 36601 20131 36635
rect 20073 36595 20131 36601
rect 20625 36635 20683 36641
rect 20625 36601 20637 36635
rect 20671 36632 20683 36635
rect 22066 36632 22094 36876
rect 23842 36864 23848 36876
rect 23900 36864 23906 36916
rect 23937 36907 23995 36913
rect 23937 36873 23949 36907
rect 23983 36904 23995 36907
rect 24026 36904 24032 36916
rect 23983 36876 24032 36904
rect 23983 36873 23995 36876
rect 23937 36867 23995 36873
rect 24026 36864 24032 36876
rect 24084 36864 24090 36916
rect 23106 36836 23112 36848
rect 20671 36604 22094 36632
rect 22296 36808 23112 36836
rect 20671 36601 20683 36604
rect 20625 36595 20683 36601
rect 11557 36536 12204 36564
rect 8481 36527 8539 36533
rect 12526 36524 12532 36576
rect 12584 36524 12590 36576
rect 17126 36524 17132 36576
rect 17184 36524 17190 36576
rect 17402 36524 17408 36576
rect 17460 36524 17466 36576
rect 17589 36567 17647 36573
rect 17589 36533 17601 36567
rect 17635 36564 17647 36567
rect 17954 36564 17960 36576
rect 17635 36536 17960 36564
rect 17635 36533 17647 36536
rect 17589 36527 17647 36533
rect 17954 36524 17960 36536
rect 18012 36524 18018 36576
rect 19613 36567 19671 36573
rect 19613 36533 19625 36567
rect 19659 36564 19671 36567
rect 20714 36564 20720 36576
rect 19659 36536 20720 36564
rect 19659 36533 19671 36536
rect 19613 36527 19671 36533
rect 20714 36524 20720 36536
rect 20772 36524 20778 36576
rect 21082 36524 21088 36576
rect 21140 36564 21146 36576
rect 22296 36564 22324 36808
rect 23106 36796 23112 36808
rect 23164 36796 23170 36848
rect 23661 36839 23719 36845
rect 23661 36805 23673 36839
rect 23707 36836 23719 36839
rect 23707 36808 24532 36836
rect 23707 36805 23719 36808
rect 23661 36799 23719 36805
rect 23014 36728 23020 36780
rect 23072 36728 23078 36780
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 24026 36768 24032 36780
rect 23339 36740 24032 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 24026 36728 24032 36740
rect 24084 36728 24090 36780
rect 24136 36777 24164 36808
rect 24504 36780 24532 36808
rect 24121 36771 24179 36777
rect 24121 36737 24133 36771
rect 24167 36737 24179 36771
rect 24121 36731 24179 36737
rect 24213 36771 24271 36777
rect 24213 36737 24225 36771
rect 24259 36737 24271 36771
rect 24213 36731 24271 36737
rect 22370 36660 22376 36712
rect 22428 36700 22434 36712
rect 24228 36700 24256 36731
rect 24486 36728 24492 36780
rect 24544 36728 24550 36780
rect 22428 36672 24256 36700
rect 22428 36660 22434 36672
rect 23109 36635 23167 36641
rect 23109 36601 23121 36635
rect 23155 36632 23167 36635
rect 23474 36632 23480 36644
rect 23155 36604 23480 36632
rect 23155 36601 23167 36604
rect 23109 36595 23167 36601
rect 23474 36592 23480 36604
rect 23532 36592 23538 36644
rect 21140 36536 22324 36564
rect 21140 36524 21146 36536
rect 22830 36524 22836 36576
rect 22888 36524 22894 36576
rect 24394 36524 24400 36576
rect 24452 36524 24458 36576
rect 1104 36474 24840 36496
rect 1104 36422 3917 36474
rect 3969 36422 3981 36474
rect 4033 36422 4045 36474
rect 4097 36422 4109 36474
rect 4161 36422 4173 36474
rect 4225 36422 9851 36474
rect 9903 36422 9915 36474
rect 9967 36422 9979 36474
rect 10031 36422 10043 36474
rect 10095 36422 10107 36474
rect 10159 36422 15785 36474
rect 15837 36422 15849 36474
rect 15901 36422 15913 36474
rect 15965 36422 15977 36474
rect 16029 36422 16041 36474
rect 16093 36422 21719 36474
rect 21771 36422 21783 36474
rect 21835 36422 21847 36474
rect 21899 36422 21911 36474
rect 21963 36422 21975 36474
rect 22027 36422 24840 36474
rect 1104 36400 24840 36422
rect 6914 36320 6920 36372
rect 6972 36360 6978 36372
rect 7009 36363 7067 36369
rect 7009 36360 7021 36363
rect 6972 36332 7021 36360
rect 6972 36320 6978 36332
rect 7009 36329 7021 36332
rect 7055 36329 7067 36363
rect 7009 36323 7067 36329
rect 11054 36320 11060 36372
rect 11112 36320 11118 36372
rect 17126 36320 17132 36372
rect 17184 36360 17190 36372
rect 21082 36360 21088 36372
rect 17184 36332 21088 36360
rect 17184 36320 17190 36332
rect 21082 36320 21088 36332
rect 21140 36320 21146 36372
rect 22370 36320 22376 36372
rect 22428 36320 22434 36372
rect 22830 36320 22836 36372
rect 22888 36320 22894 36372
rect 23385 36363 23443 36369
rect 23385 36329 23397 36363
rect 23431 36360 23443 36363
rect 23566 36360 23572 36372
rect 23431 36332 23572 36360
rect 23431 36329 23443 36332
rect 23385 36323 23443 36329
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 3878 36292 3884 36304
rect 2700 36264 3884 36292
rect 1302 36116 1308 36168
rect 1360 36156 1366 36168
rect 1489 36159 1547 36165
rect 1489 36156 1501 36159
rect 1360 36128 1501 36156
rect 1360 36116 1366 36128
rect 1489 36125 1501 36128
rect 1535 36125 1547 36159
rect 1489 36119 1547 36125
rect 1763 36159 1821 36165
rect 1763 36125 1775 36159
rect 1809 36156 1821 36159
rect 2700 36156 2728 36264
rect 3878 36252 3884 36264
rect 3936 36252 3942 36304
rect 4890 36252 4896 36304
rect 4948 36292 4954 36304
rect 4948 36264 5488 36292
rect 4948 36252 4954 36264
rect 2774 36184 2780 36236
rect 2832 36224 2838 36236
rect 4709 36227 4767 36233
rect 4709 36224 4721 36227
rect 2832 36196 4721 36224
rect 2832 36184 2838 36196
rect 4709 36193 4721 36196
rect 4755 36224 4767 36227
rect 5460 36224 5488 36264
rect 5718 36252 5724 36304
rect 5776 36252 5782 36304
rect 7282 36292 7288 36304
rect 6654 36264 7288 36292
rect 6654 36224 6682 36264
rect 7282 36252 7288 36264
rect 7340 36292 7346 36304
rect 10965 36295 11023 36301
rect 7340 36264 8340 36292
rect 7340 36252 7346 36264
rect 4755 36196 5396 36224
rect 5460 36196 6682 36224
rect 6917 36227 6975 36233
rect 4755 36193 4767 36196
rect 4709 36187 4767 36193
rect 1809 36128 2728 36156
rect 2869 36159 2927 36165
rect 1809 36125 1821 36128
rect 1763 36119 1821 36125
rect 2869 36125 2881 36159
rect 2915 36156 2927 36159
rect 2958 36156 2964 36168
rect 2915 36128 2964 36156
rect 2915 36125 2927 36128
rect 2869 36119 2927 36125
rect 2958 36116 2964 36128
rect 3016 36116 3022 36168
rect 3786 36116 3792 36168
rect 3844 36116 3850 36168
rect 4798 36116 4804 36168
rect 4856 36156 4862 36168
rect 5077 36159 5135 36165
rect 5077 36156 5089 36159
rect 4856 36128 5089 36156
rect 4856 36116 4862 36128
rect 5077 36125 5089 36128
rect 5123 36156 5135 36159
rect 5166 36156 5172 36168
rect 5123 36128 5172 36156
rect 5123 36125 5135 36128
rect 5077 36119 5135 36125
rect 5166 36116 5172 36128
rect 5224 36116 5230 36168
rect 5261 36159 5319 36165
rect 5261 36125 5273 36159
rect 5307 36125 5319 36159
rect 5368 36156 5396 36196
rect 6917 36193 6929 36227
rect 6963 36224 6975 36227
rect 7374 36224 7380 36236
rect 6963 36196 7380 36224
rect 6963 36193 6975 36196
rect 6917 36187 6975 36193
rect 7374 36184 7380 36196
rect 7432 36184 7438 36236
rect 8312 36168 8340 36264
rect 10965 36261 10977 36295
rect 11011 36292 11023 36295
rect 11072 36292 11100 36320
rect 11011 36264 11100 36292
rect 18509 36295 18567 36301
rect 11011 36261 11023 36264
rect 10965 36255 11023 36261
rect 18509 36261 18521 36295
rect 18555 36261 18567 36295
rect 18509 36255 18567 36261
rect 11238 36184 11244 36236
rect 11296 36184 11302 36236
rect 12526 36224 12532 36236
rect 11557 36196 12532 36224
rect 5442 36156 5448 36168
rect 5368 36128 5448 36156
rect 5261 36119 5319 36125
rect 382 36048 388 36100
rect 440 36088 446 36100
rect 1854 36088 1860 36100
rect 440 36060 1860 36088
rect 440 36048 446 36060
rect 1854 36048 1860 36060
rect 1912 36048 1918 36100
rect 2406 36048 2412 36100
rect 2464 36088 2470 36100
rect 3145 36091 3203 36097
rect 3145 36088 3157 36091
rect 2464 36060 3157 36088
rect 2464 36048 2470 36060
rect 3145 36057 3157 36060
rect 3191 36057 3203 36091
rect 3145 36051 3203 36057
rect 4062 36048 4068 36100
rect 4120 36048 4126 36100
rect 4433 36091 4491 36097
rect 4433 36057 4445 36091
rect 4479 36057 4491 36091
rect 4433 36051 4491 36057
rect 2501 36023 2559 36029
rect 2501 35989 2513 36023
rect 2547 36020 2559 36023
rect 2682 36020 2688 36032
rect 2547 35992 2688 36020
rect 2547 35989 2559 35992
rect 2501 35983 2559 35989
rect 2682 35980 2688 35992
rect 2740 35980 2746 36032
rect 3418 35980 3424 36032
rect 3476 36020 3482 36032
rect 4448 36020 4476 36051
rect 3476 35992 4476 36020
rect 3476 35980 3482 35992
rect 4706 35980 4712 36032
rect 4764 36020 4770 36032
rect 5166 36020 5172 36032
rect 4764 35992 5172 36020
rect 4764 35980 4770 35992
rect 5166 35980 5172 35992
rect 5224 35980 5230 36032
rect 5276 36020 5304 36119
rect 5442 36116 5448 36128
rect 5500 36116 5506 36168
rect 5994 36116 6000 36168
rect 6052 36116 6058 36168
rect 6086 36116 6092 36168
rect 6144 36165 6150 36168
rect 6144 36159 6172 36165
rect 6160 36125 6172 36159
rect 6144 36119 6172 36125
rect 6144 36116 6150 36119
rect 6270 36116 6276 36168
rect 6328 36116 6334 36168
rect 7193 36159 7251 36165
rect 7193 36125 7205 36159
rect 7239 36156 7251 36159
rect 7282 36156 7288 36168
rect 7239 36128 7288 36156
rect 7239 36125 7251 36128
rect 7193 36119 7251 36125
rect 7282 36116 7288 36128
rect 7340 36116 7346 36168
rect 8294 36116 8300 36168
rect 8352 36156 8358 36168
rect 8846 36156 8852 36168
rect 8352 36128 8852 36156
rect 8352 36116 8358 36128
rect 8846 36116 8852 36128
rect 8904 36156 8910 36168
rect 8941 36159 8999 36165
rect 8941 36156 8953 36159
rect 8904 36128 8953 36156
rect 8904 36116 8910 36128
rect 8941 36125 8953 36128
rect 8987 36125 8999 36159
rect 8941 36119 8999 36125
rect 9122 36116 9128 36168
rect 9180 36156 9186 36168
rect 9215 36159 9273 36165
rect 9215 36156 9227 36159
rect 9180 36128 9227 36156
rect 9180 36116 9186 36128
rect 9215 36125 9227 36128
rect 9261 36125 9273 36159
rect 9215 36119 9273 36125
rect 9766 36116 9772 36168
rect 9824 36156 9830 36168
rect 10321 36159 10379 36165
rect 10321 36156 10333 36159
rect 9824 36128 10333 36156
rect 9824 36116 9830 36128
rect 10321 36125 10333 36128
rect 10367 36125 10379 36159
rect 10321 36119 10379 36125
rect 10502 36116 10508 36168
rect 10560 36116 10566 36168
rect 11330 36116 11336 36168
rect 11388 36165 11394 36168
rect 11557 36165 11585 36196
rect 12526 36184 12532 36196
rect 12584 36184 12590 36236
rect 11388 36159 11416 36165
rect 11404 36125 11416 36159
rect 11388 36119 11416 36125
rect 11527 36159 11585 36165
rect 11527 36125 11539 36159
rect 11573 36125 11585 36159
rect 11527 36119 11585 36125
rect 17129 36159 17187 36165
rect 17129 36125 17141 36159
rect 17175 36156 17187 36159
rect 17218 36156 17224 36168
rect 17175 36128 17224 36156
rect 17175 36125 17187 36128
rect 17129 36119 17187 36125
rect 11388 36116 11394 36119
rect 17218 36116 17224 36128
rect 17276 36156 17282 36168
rect 17862 36156 17868 36168
rect 17276 36128 17868 36156
rect 17276 36116 17282 36128
rect 17862 36116 17868 36128
rect 17920 36116 17926 36168
rect 18524 36156 18552 36255
rect 20254 36252 20260 36304
rect 20312 36292 20318 36304
rect 20806 36292 20812 36304
rect 20312 36264 20812 36292
rect 20312 36252 20318 36264
rect 20806 36252 20812 36264
rect 20864 36252 20870 36304
rect 20993 36295 21051 36301
rect 20993 36261 21005 36295
rect 21039 36261 21051 36295
rect 20993 36255 21051 36261
rect 20530 36224 20536 36236
rect 19306 36196 20536 36224
rect 18785 36159 18843 36165
rect 18785 36156 18797 36159
rect 18524 36128 18797 36156
rect 18785 36125 18797 36128
rect 18831 36125 18843 36159
rect 18785 36119 18843 36125
rect 17402 36097 17408 36100
rect 12161 36091 12219 36097
rect 12161 36057 12173 36091
rect 12207 36088 12219 36091
rect 17374 36091 17408 36097
rect 17374 36088 17386 36091
rect 12207 36060 17386 36088
rect 12207 36057 12219 36060
rect 12161 36051 12219 36057
rect 17374 36057 17386 36060
rect 17374 36051 17408 36057
rect 17402 36048 17408 36051
rect 17460 36048 17466 36100
rect 17770 36048 17776 36100
rect 17828 36088 17834 36100
rect 19306 36088 19334 36196
rect 20530 36184 20536 36196
rect 20588 36184 20594 36236
rect 21008 36224 21036 36255
rect 22848 36224 22876 36320
rect 21008 36196 21864 36224
rect 22848 36196 23888 36224
rect 21836 36165 21864 36196
rect 21177 36159 21235 36165
rect 21177 36156 21189 36159
rect 17828 36060 19334 36088
rect 19812 36128 21189 36156
rect 17828 36048 17834 36060
rect 19812 36032 19840 36128
rect 21177 36125 21189 36128
rect 21223 36125 21235 36159
rect 21177 36119 21235 36125
rect 21821 36159 21879 36165
rect 21821 36125 21833 36159
rect 21867 36125 21879 36159
rect 22557 36159 22615 36165
rect 22557 36156 22569 36159
rect 21821 36119 21879 36125
rect 22066 36128 22569 36156
rect 5626 36020 5632 36032
rect 5276 35992 5632 36020
rect 5626 35980 5632 35992
rect 5684 35980 5690 36032
rect 7558 35980 7564 36032
rect 7616 36020 7622 36032
rect 8110 36020 8116 36032
rect 7616 35992 8116 36020
rect 7616 35980 7622 35992
rect 8110 35980 8116 35992
rect 8168 35980 8174 36032
rect 8570 35980 8576 36032
rect 8628 36020 8634 36032
rect 9953 36023 10011 36029
rect 9953 36020 9965 36023
rect 8628 35992 9965 36020
rect 8628 35980 8634 35992
rect 9953 35989 9965 35992
rect 9999 35989 10011 36023
rect 9953 35983 10011 35989
rect 11330 35980 11336 36032
rect 11388 36020 11394 36032
rect 11606 36020 11612 36032
rect 11388 35992 11612 36020
rect 11388 35980 11394 35992
rect 11606 35980 11612 35992
rect 11664 35980 11670 36032
rect 12250 35980 12256 36032
rect 12308 36020 12314 36032
rect 12618 36020 12624 36032
rect 12308 35992 12624 36020
rect 12308 35980 12314 35992
rect 12618 35980 12624 35992
rect 12676 35980 12682 36032
rect 18601 36023 18659 36029
rect 18601 35989 18613 36023
rect 18647 36020 18659 36023
rect 19334 36020 19340 36032
rect 18647 35992 19340 36020
rect 18647 35989 18659 35992
rect 18601 35983 18659 35989
rect 19334 35980 19340 35992
rect 19392 35980 19398 36032
rect 19794 35980 19800 36032
rect 19852 35980 19858 36032
rect 21637 36023 21695 36029
rect 21637 35989 21649 36023
rect 21683 36020 21695 36023
rect 22066 36020 22094 36128
rect 22557 36125 22569 36128
rect 22603 36125 22615 36159
rect 22557 36119 22615 36125
rect 23566 36116 23572 36168
rect 23624 36116 23630 36168
rect 23860 36165 23888 36196
rect 23845 36159 23903 36165
rect 23845 36125 23857 36159
rect 23891 36125 23903 36159
rect 23845 36119 23903 36125
rect 24213 36091 24271 36097
rect 24213 36057 24225 36091
rect 24259 36088 24271 36091
rect 25130 36088 25136 36100
rect 24259 36060 25136 36088
rect 24259 36057 24271 36060
rect 24213 36051 24271 36057
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 21683 35992 22094 36020
rect 21683 35989 21695 35992
rect 21637 35983 21695 35989
rect 1104 35930 25000 35952
rect 1104 35878 6884 35930
rect 6936 35878 6948 35930
rect 7000 35878 7012 35930
rect 7064 35878 7076 35930
rect 7128 35878 7140 35930
rect 7192 35878 12818 35930
rect 12870 35878 12882 35930
rect 12934 35878 12946 35930
rect 12998 35878 13010 35930
rect 13062 35878 13074 35930
rect 13126 35878 18752 35930
rect 18804 35878 18816 35930
rect 18868 35878 18880 35930
rect 18932 35878 18944 35930
rect 18996 35878 19008 35930
rect 19060 35878 24686 35930
rect 24738 35878 24750 35930
rect 24802 35878 24814 35930
rect 24866 35878 24878 35930
rect 24930 35878 24942 35930
rect 24994 35878 25000 35930
rect 1104 35856 25000 35878
rect 3329 35819 3387 35825
rect 3329 35785 3341 35819
rect 3375 35816 3387 35819
rect 3510 35816 3516 35828
rect 3375 35788 3516 35816
rect 3375 35785 3387 35788
rect 3329 35779 3387 35785
rect 3510 35776 3516 35788
rect 3568 35776 3574 35828
rect 6181 35819 6239 35825
rect 4080 35788 6132 35816
rect 1489 35683 1547 35689
rect 1489 35649 1501 35683
rect 1535 35680 1547 35683
rect 1854 35680 1860 35692
rect 1535 35652 1860 35680
rect 1535 35649 1547 35652
rect 1489 35643 1547 35649
rect 1854 35640 1860 35652
rect 1912 35640 1918 35692
rect 2682 35640 2688 35692
rect 2740 35640 2746 35692
rect 3418 35640 3424 35692
rect 3476 35640 3482 35692
rect 4080 35680 4108 35788
rect 6104 35760 6132 35788
rect 6181 35785 6193 35819
rect 6227 35816 6239 35819
rect 7282 35816 7288 35828
rect 6227 35788 7288 35816
rect 6227 35785 6239 35788
rect 6181 35779 6239 35785
rect 7282 35776 7288 35788
rect 7340 35776 7346 35828
rect 8205 35819 8263 35825
rect 8205 35785 8217 35819
rect 8251 35816 8263 35819
rect 8938 35816 8944 35828
rect 8251 35788 8944 35816
rect 8251 35785 8263 35788
rect 8205 35779 8263 35785
rect 8938 35776 8944 35788
rect 8996 35776 9002 35828
rect 9214 35776 9220 35828
rect 9272 35776 9278 35828
rect 9582 35776 9588 35828
rect 9640 35816 9646 35828
rect 11882 35816 11888 35828
rect 9640 35788 11888 35816
rect 9640 35776 9646 35788
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 14185 35819 14243 35825
rect 14185 35816 14197 35819
rect 12084 35788 14197 35816
rect 4522 35708 4528 35760
rect 4580 35708 4586 35760
rect 6086 35708 6092 35760
rect 6144 35708 6150 35760
rect 8570 35708 8576 35760
rect 8628 35708 8634 35760
rect 9232 35748 9260 35776
rect 8680 35720 9260 35748
rect 9309 35751 9367 35757
rect 4540 35680 4568 35708
rect 3528 35652 4108 35680
rect 4172 35652 4568 35680
rect 8481 35683 8539 35689
rect 1673 35615 1731 35621
rect 1673 35581 1685 35615
rect 1719 35612 1731 35615
rect 2038 35612 2044 35624
rect 1719 35584 2044 35612
rect 1719 35581 1731 35584
rect 1673 35575 1731 35581
rect 2038 35572 2044 35584
rect 2096 35572 2102 35624
rect 2409 35615 2467 35621
rect 2409 35612 2421 35615
rect 2240 35584 2421 35612
rect 2130 35504 2136 35556
rect 2188 35504 2194 35556
rect 1762 35436 1768 35488
rect 1820 35476 1826 35488
rect 2038 35476 2044 35488
rect 1820 35448 2044 35476
rect 1820 35436 1826 35448
rect 2038 35436 2044 35448
rect 2096 35436 2102 35488
rect 2240 35476 2268 35584
rect 2409 35581 2421 35584
rect 2455 35581 2467 35615
rect 2409 35575 2467 35581
rect 2547 35615 2605 35621
rect 2547 35581 2559 35615
rect 2593 35612 2605 35615
rect 3528 35612 3556 35652
rect 2593 35584 3556 35612
rect 2593 35581 2605 35584
rect 2547 35575 2605 35581
rect 3602 35572 3608 35624
rect 3660 35612 3666 35624
rect 3878 35612 3884 35624
rect 3660 35584 3884 35612
rect 3660 35572 3666 35584
rect 3878 35572 3884 35584
rect 3936 35572 3942 35624
rect 3050 35476 3056 35488
rect 2240 35448 3056 35476
rect 3050 35436 3056 35448
rect 3108 35476 3114 35488
rect 4172 35476 4200 35652
rect 8481 35649 8493 35683
rect 8527 35680 8539 35683
rect 8680 35680 8708 35720
rect 9309 35717 9321 35751
rect 9355 35748 9367 35751
rect 9398 35748 9404 35760
rect 9355 35720 9404 35748
rect 9355 35717 9367 35720
rect 9309 35711 9367 35717
rect 9398 35708 9404 35720
rect 9456 35708 9462 35760
rect 9674 35748 9680 35760
rect 9600 35720 9680 35748
rect 8527 35652 8708 35680
rect 8527 35649 8539 35652
rect 8481 35643 8539 35649
rect 8846 35640 8852 35692
rect 8904 35680 8910 35692
rect 8941 35683 8999 35689
rect 8941 35680 8953 35683
rect 8904 35652 8953 35680
rect 8904 35640 8910 35652
rect 8941 35649 8953 35652
rect 8987 35680 8999 35683
rect 9600 35680 9628 35720
rect 9674 35708 9680 35720
rect 9732 35708 9738 35760
rect 11514 35748 11520 35760
rect 9966 35720 11520 35748
rect 9966 35719 9994 35720
rect 9935 35713 9994 35719
rect 8987 35652 9628 35680
rect 9935 35679 9947 35713
rect 9981 35682 9994 35713
rect 9981 35679 9993 35682
rect 9935 35673 9993 35679
rect 8987 35649 8999 35652
rect 8941 35643 8999 35649
rect 4341 35615 4399 35621
rect 4341 35581 4353 35615
rect 4387 35581 4399 35615
rect 4341 35575 4399 35581
rect 4356 35544 4384 35575
rect 4522 35572 4528 35624
rect 4580 35572 4586 35624
rect 5258 35572 5264 35624
rect 5316 35572 5322 35624
rect 5442 35621 5448 35624
rect 5399 35615 5448 35621
rect 5399 35581 5411 35615
rect 5445 35581 5448 35615
rect 5399 35575 5448 35581
rect 5442 35572 5448 35575
rect 5500 35572 5506 35624
rect 5537 35615 5595 35621
rect 5537 35581 5549 35615
rect 5583 35612 5595 35615
rect 6270 35612 6276 35624
rect 5583 35584 6276 35612
rect 5583 35581 5595 35584
rect 5537 35575 5595 35581
rect 6270 35572 6276 35584
rect 6328 35572 6334 35624
rect 8386 35572 8392 35624
rect 8444 35572 8450 35624
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 4706 35544 4712 35556
rect 4356 35516 4712 35544
rect 4706 35504 4712 35516
rect 4764 35504 4770 35556
rect 4985 35547 5043 35553
rect 4985 35513 4997 35547
rect 5031 35513 5043 35547
rect 4985 35507 5043 35513
rect 3108 35448 4200 35476
rect 5000 35476 5028 35507
rect 5718 35476 5724 35488
rect 5000 35448 5724 35476
rect 3108 35436 3114 35448
rect 5718 35436 5724 35448
rect 5776 35436 5782 35488
rect 5902 35436 5908 35488
rect 5960 35476 5966 35488
rect 7466 35476 7472 35488
rect 5960 35448 7472 35476
rect 5960 35436 5966 35448
rect 7466 35436 7472 35448
rect 7524 35436 7530 35488
rect 9398 35436 9404 35488
rect 9456 35476 9462 35488
rect 9493 35479 9551 35485
rect 9493 35476 9505 35479
rect 9456 35448 9505 35476
rect 9456 35436 9462 35448
rect 9493 35445 9505 35448
rect 9539 35445 9551 35479
rect 9493 35439 9551 35445
rect 9582 35436 9588 35488
rect 9640 35476 9646 35488
rect 10334 35476 10362 35720
rect 11514 35708 11520 35720
rect 11572 35708 11578 35760
rect 11698 35708 11704 35760
rect 11756 35708 11762 35760
rect 11974 35708 11980 35760
rect 12032 35708 12038 35760
rect 12084 35757 12112 35788
rect 14185 35785 14197 35788
rect 14231 35785 14243 35819
rect 14185 35779 14243 35785
rect 19334 35776 19340 35828
rect 19392 35776 19398 35828
rect 21085 35819 21143 35825
rect 21085 35785 21097 35819
rect 21131 35785 21143 35819
rect 21085 35779 21143 35785
rect 21821 35819 21879 35825
rect 21821 35785 21833 35819
rect 21867 35816 21879 35819
rect 21867 35788 22324 35816
rect 21867 35785 21879 35788
rect 21821 35779 21879 35785
rect 12069 35751 12127 35757
rect 12069 35717 12081 35751
rect 12115 35717 12127 35751
rect 12069 35711 12127 35717
rect 12158 35708 12164 35760
rect 12216 35748 12222 35760
rect 12805 35751 12863 35757
rect 12805 35748 12817 35751
rect 12216 35720 12817 35748
rect 12216 35708 12222 35720
rect 12805 35717 12817 35720
rect 12851 35717 12863 35751
rect 12805 35711 12863 35717
rect 13814 35708 13820 35760
rect 13872 35748 13878 35760
rect 18230 35748 18236 35760
rect 13872 35720 18236 35748
rect 13872 35708 13878 35720
rect 18230 35708 18236 35720
rect 18288 35708 18294 35760
rect 19352 35748 19380 35776
rect 21100 35748 21128 35779
rect 19352 35720 19564 35748
rect 21100 35720 21772 35748
rect 11606 35680 11612 35692
rect 10520 35652 11612 35680
rect 9640 35448 10362 35476
rect 9640 35436 9646 35448
rect 10410 35436 10416 35488
rect 10468 35476 10474 35488
rect 10520 35476 10548 35652
rect 11606 35640 11612 35652
rect 11664 35680 11670 35692
rect 12437 35683 12495 35689
rect 12437 35680 12449 35683
rect 11664 35652 12449 35680
rect 11664 35640 11670 35652
rect 12437 35649 12449 35652
rect 12483 35649 12495 35683
rect 12437 35643 12495 35649
rect 12618 35640 12624 35692
rect 12676 35680 12682 35692
rect 13447 35683 13505 35689
rect 13447 35680 13459 35683
rect 12676 35652 13459 35680
rect 12676 35640 12682 35652
rect 13447 35649 13459 35652
rect 13493 35680 13505 35683
rect 13493 35652 15976 35680
rect 13493 35649 13505 35652
rect 13447 35643 13505 35649
rect 12802 35612 12808 35624
rect 12742 35584 12808 35612
rect 12802 35572 12808 35584
rect 12860 35572 12866 35624
rect 13173 35615 13231 35621
rect 13173 35581 13185 35615
rect 13219 35581 13231 35615
rect 13173 35575 13231 35581
rect 12986 35504 12992 35556
rect 13044 35504 13050 35556
rect 13188 35544 13216 35575
rect 13188 35516 13308 35544
rect 10468 35448 10548 35476
rect 10689 35479 10747 35485
rect 10468 35436 10474 35448
rect 10689 35445 10701 35479
rect 10735 35476 10747 35479
rect 11054 35476 11060 35488
rect 10735 35448 11060 35476
rect 10735 35445 10747 35448
rect 10689 35439 10747 35445
rect 11054 35436 11060 35448
rect 11112 35436 11118 35488
rect 13280 35476 13308 35516
rect 14182 35476 14188 35488
rect 13280 35448 14188 35476
rect 14182 35436 14188 35448
rect 14240 35476 14246 35488
rect 15470 35476 15476 35488
rect 14240 35448 15476 35476
rect 14240 35436 14246 35448
rect 15470 35436 15476 35448
rect 15528 35436 15534 35488
rect 15948 35476 15976 35652
rect 16850 35640 16856 35692
rect 16908 35680 16914 35692
rect 19536 35689 19564 35720
rect 17831 35683 17889 35689
rect 17831 35680 17843 35683
rect 16908 35652 17843 35680
rect 16908 35640 16914 35652
rect 17831 35649 17843 35652
rect 17877 35649 17889 35683
rect 18969 35683 19027 35689
rect 18969 35680 18981 35683
rect 17831 35643 17889 35649
rect 18616 35652 18981 35680
rect 17586 35572 17592 35624
rect 17644 35572 17650 35624
rect 18616 35553 18644 35652
rect 18969 35649 18981 35652
rect 19015 35680 19027 35683
rect 19337 35683 19395 35689
rect 19337 35680 19349 35683
rect 19015 35652 19349 35680
rect 19015 35649 19027 35652
rect 18969 35643 19027 35649
rect 19337 35649 19349 35652
rect 19383 35649 19395 35683
rect 19337 35643 19395 35649
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 19521 35643 19579 35649
rect 21266 35640 21272 35692
rect 21324 35640 21330 35692
rect 21744 35680 21772 35720
rect 22005 35683 22063 35689
rect 22005 35680 22017 35683
rect 21744 35652 22017 35680
rect 22005 35649 22017 35652
rect 22051 35649 22063 35683
rect 22296 35680 22324 35788
rect 23014 35776 23020 35828
rect 23072 35816 23078 35828
rect 23109 35819 23167 35825
rect 23109 35816 23121 35819
rect 23072 35788 23121 35816
rect 23072 35776 23078 35788
rect 23109 35785 23121 35788
rect 23155 35785 23167 35819
rect 23109 35779 23167 35785
rect 23477 35819 23535 35825
rect 23477 35785 23489 35819
rect 23523 35816 23535 35819
rect 23566 35816 23572 35828
rect 23523 35788 23572 35816
rect 23523 35785 23535 35788
rect 23477 35779 23535 35785
rect 23566 35776 23572 35788
rect 23624 35776 23630 35828
rect 25314 35748 25320 35760
rect 23676 35720 25320 35748
rect 23676 35689 23704 35720
rect 25314 35708 25320 35720
rect 25372 35708 25378 35760
rect 22557 35683 22615 35689
rect 22557 35680 22569 35683
rect 22296 35652 22569 35680
rect 22005 35643 22063 35649
rect 22557 35649 22569 35652
rect 22603 35649 22615 35683
rect 22833 35683 22891 35689
rect 22833 35680 22845 35683
rect 22557 35643 22615 35649
rect 22664 35652 22845 35680
rect 19245 35615 19303 35621
rect 19245 35581 19257 35615
rect 19291 35612 19303 35615
rect 19429 35615 19487 35621
rect 19429 35612 19441 35615
rect 19291 35584 19441 35612
rect 19291 35581 19303 35584
rect 19245 35575 19303 35581
rect 19429 35581 19441 35584
rect 19475 35581 19487 35615
rect 22370 35612 22376 35624
rect 19429 35575 19487 35581
rect 22066 35584 22376 35612
rect 18601 35547 18659 35553
rect 18601 35513 18613 35547
rect 18647 35513 18659 35547
rect 22066 35544 22094 35584
rect 22370 35572 22376 35584
rect 22428 35612 22434 35624
rect 22664 35612 22692 35652
rect 22833 35649 22845 35652
rect 22879 35649 22891 35683
rect 22833 35643 22891 35649
rect 23293 35683 23351 35689
rect 23293 35649 23305 35683
rect 23339 35649 23351 35683
rect 23293 35643 23351 35649
rect 23661 35683 23719 35689
rect 23661 35649 23673 35683
rect 23707 35649 23719 35683
rect 23661 35643 23719 35649
rect 22428 35584 22692 35612
rect 22428 35572 22434 35584
rect 18601 35507 18659 35513
rect 18708 35516 22094 35544
rect 22649 35547 22707 35553
rect 18708 35476 18736 35516
rect 22649 35513 22661 35547
rect 22695 35544 22707 35547
rect 23308 35544 23336 35643
rect 23934 35640 23940 35692
rect 23992 35640 23998 35692
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35649 24179 35683
rect 24121 35643 24179 35649
rect 24136 35612 24164 35643
rect 22695 35516 23336 35544
rect 23676 35584 24164 35612
rect 22695 35513 22707 35516
rect 22649 35507 22707 35513
rect 15948 35448 18736 35476
rect 19058 35436 19064 35488
rect 19116 35436 19122 35488
rect 19153 35479 19211 35485
rect 19153 35445 19165 35479
rect 19199 35476 19211 35479
rect 21174 35476 21180 35488
rect 19199 35448 21180 35476
rect 19199 35445 19211 35448
rect 19153 35439 19211 35445
rect 21174 35436 21180 35448
rect 21232 35436 21238 35488
rect 22373 35479 22431 35485
rect 22373 35445 22385 35479
rect 22419 35476 22431 35479
rect 23676 35476 23704 35584
rect 22419 35448 23704 35476
rect 22419 35445 22431 35448
rect 22373 35439 22431 35445
rect 23750 35436 23756 35488
rect 23808 35436 23814 35488
rect 24394 35436 24400 35488
rect 24452 35436 24458 35488
rect 1104 35386 24840 35408
rect 1104 35334 3917 35386
rect 3969 35334 3981 35386
rect 4033 35334 4045 35386
rect 4097 35334 4109 35386
rect 4161 35334 4173 35386
rect 4225 35334 9851 35386
rect 9903 35334 9915 35386
rect 9967 35334 9979 35386
rect 10031 35334 10043 35386
rect 10095 35334 10107 35386
rect 10159 35334 15785 35386
rect 15837 35334 15849 35386
rect 15901 35334 15913 35386
rect 15965 35334 15977 35386
rect 16029 35334 16041 35386
rect 16093 35334 21719 35386
rect 21771 35334 21783 35386
rect 21835 35334 21847 35386
rect 21899 35334 21911 35386
rect 21963 35334 21975 35386
rect 22027 35334 24840 35386
rect 1104 35312 24840 35334
rect 3234 35272 3240 35284
rect 1688 35244 3240 35272
rect 1688 35145 1716 35244
rect 3234 35232 3240 35244
rect 3292 35232 3298 35284
rect 5261 35275 5319 35281
rect 5261 35241 5273 35275
rect 5307 35241 5319 35275
rect 5261 35235 5319 35241
rect 3329 35207 3387 35213
rect 3329 35173 3341 35207
rect 3375 35173 3387 35207
rect 3329 35167 3387 35173
rect 1673 35139 1731 35145
rect 1673 35105 1685 35139
rect 1719 35105 1731 35139
rect 3344 35136 3372 35167
rect 5276 35148 5304 35235
rect 5534 35232 5540 35284
rect 5592 35272 5598 35284
rect 6178 35272 6184 35284
rect 5592 35244 6184 35272
rect 5592 35232 5598 35244
rect 6178 35232 6184 35244
rect 6236 35232 6242 35284
rect 6270 35232 6276 35284
rect 6328 35272 6334 35284
rect 6457 35275 6515 35281
rect 6457 35272 6469 35275
rect 6328 35244 6469 35272
rect 6328 35232 6334 35244
rect 6457 35241 6469 35244
rect 6503 35241 6515 35275
rect 9582 35272 9588 35284
rect 6457 35235 6515 35241
rect 7208 35244 9588 35272
rect 5552 35204 5580 35232
rect 5460 35176 5580 35204
rect 3344 35108 3818 35136
rect 1673 35099 1731 35105
rect 5258 35096 5264 35148
rect 5316 35096 5322 35148
rect 5460 35145 5488 35176
rect 5445 35139 5503 35145
rect 5445 35105 5457 35139
rect 5491 35105 5503 35139
rect 5445 35099 5503 35105
rect 750 35028 756 35080
rect 808 35068 814 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 808 35040 1409 35068
rect 808 35028 814 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 2314 35028 2320 35080
rect 2372 35028 2378 35080
rect 2498 35028 2504 35080
rect 2556 35068 2562 35080
rect 2591 35071 2649 35077
rect 2591 35068 2603 35071
rect 2556 35040 2603 35068
rect 2556 35028 2562 35040
rect 2591 35037 2603 35040
rect 2637 35037 2649 35071
rect 3234 35068 3240 35080
rect 2591 35031 2649 35037
rect 2700 35040 3240 35068
rect 2332 35000 2360 35028
rect 2700 35000 2728 35040
rect 3234 35028 3240 35040
rect 3292 35028 3298 35080
rect 4246 35028 4252 35080
rect 4304 35028 4310 35080
rect 5718 35068 5724 35080
rect 5679 35040 5724 35068
rect 5718 35028 5724 35040
rect 5776 35068 5782 35080
rect 7208 35068 7236 35244
rect 9582 35232 9588 35244
rect 9640 35232 9646 35284
rect 10410 35232 10416 35284
rect 10468 35232 10474 35284
rect 11054 35272 11060 35284
rect 10520 35244 11060 35272
rect 7926 35164 7932 35216
rect 7984 35204 7990 35216
rect 10428 35204 10456 35232
rect 7984 35176 10456 35204
rect 7984 35164 7990 35176
rect 7282 35096 7288 35148
rect 7340 35136 7346 35148
rect 10045 35139 10103 35145
rect 10045 35136 10057 35139
rect 7340 35108 10057 35136
rect 7340 35096 7346 35108
rect 10045 35105 10057 35108
rect 10091 35136 10103 35139
rect 10410 35136 10416 35148
rect 10091 35108 10416 35136
rect 10091 35105 10103 35108
rect 10045 35099 10103 35105
rect 10410 35096 10416 35108
rect 10468 35096 10474 35148
rect 10520 35145 10548 35244
rect 11054 35232 11060 35244
rect 11112 35232 11118 35284
rect 11701 35275 11759 35281
rect 11701 35241 11713 35275
rect 11747 35272 11759 35275
rect 11747 35244 12756 35272
rect 11747 35241 11759 35244
rect 11701 35235 11759 35241
rect 12728 35204 12756 35244
rect 12802 35232 12808 35284
rect 12860 35232 12866 35284
rect 13538 35232 13544 35284
rect 13596 35272 13602 35284
rect 18233 35275 18291 35281
rect 13596 35244 16344 35272
rect 13596 35232 13602 35244
rect 13814 35204 13820 35216
rect 12728 35176 13820 35204
rect 13814 35164 13820 35176
rect 13872 35164 13878 35216
rect 10505 35139 10563 35145
rect 10505 35105 10517 35139
rect 10551 35105 10563 35139
rect 10505 35099 10563 35105
rect 10919 35139 10977 35145
rect 10919 35105 10931 35139
rect 10965 35136 10977 35139
rect 11606 35136 11612 35148
rect 10965 35108 11612 35136
rect 10965 35105 10977 35108
rect 10919 35099 10977 35105
rect 11606 35096 11612 35108
rect 11664 35096 11670 35148
rect 15470 35096 15476 35148
rect 15528 35136 15534 35148
rect 15657 35139 15715 35145
rect 15657 35136 15669 35139
rect 15528 35108 15669 35136
rect 15528 35096 15534 35108
rect 15657 35105 15669 35108
rect 15703 35105 15715 35139
rect 16316 35136 16344 35244
rect 18233 35241 18245 35275
rect 18279 35272 18291 35275
rect 19058 35272 19064 35284
rect 18279 35244 19064 35272
rect 18279 35241 18291 35244
rect 18233 35235 18291 35241
rect 19058 35232 19064 35244
rect 19116 35232 19122 35284
rect 19978 35272 19984 35284
rect 19352 35244 19984 35272
rect 16666 35164 16672 35216
rect 16724 35204 16730 35216
rect 17126 35204 17132 35216
rect 16724 35176 17132 35204
rect 16724 35164 16730 35176
rect 17126 35164 17132 35176
rect 17184 35164 17190 35216
rect 17586 35164 17592 35216
rect 17644 35204 17650 35216
rect 19352 35204 19380 35244
rect 19978 35232 19984 35244
rect 20036 35232 20042 35284
rect 22278 35232 22284 35284
rect 22336 35272 22342 35284
rect 23201 35275 23259 35281
rect 23201 35272 23213 35275
rect 22336 35244 23213 35272
rect 22336 35232 22342 35244
rect 23201 35241 23213 35244
rect 23247 35241 23259 35275
rect 23201 35235 23259 35241
rect 23658 35232 23664 35284
rect 23716 35272 23722 35284
rect 24578 35272 24584 35284
rect 23716 35244 24584 35272
rect 23716 35232 23722 35244
rect 24578 35232 24584 35244
rect 24636 35232 24642 35284
rect 20622 35204 20628 35216
rect 17644 35176 19380 35204
rect 19812 35176 20628 35204
rect 17644 35164 17650 35176
rect 19812 35136 19840 35176
rect 20622 35164 20628 35176
rect 20680 35164 20686 35216
rect 20809 35207 20867 35213
rect 20809 35173 20821 35207
rect 20855 35204 20867 35207
rect 20855 35176 23980 35204
rect 20855 35173 20867 35176
rect 20809 35167 20867 35173
rect 16316 35108 19840 35136
rect 15657 35099 15715 35105
rect 21174 35096 21180 35148
rect 21232 35136 21238 35148
rect 21232 35108 22094 35136
rect 21232 35096 21238 35108
rect 5776 35040 7236 35068
rect 5776 35028 5782 35040
rect 8938 35028 8944 35080
rect 8996 35068 9002 35080
rect 9766 35068 9772 35080
rect 8996 35040 9772 35068
rect 8996 35028 9002 35040
rect 9766 35028 9772 35040
rect 9824 35068 9830 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9824 35040 9873 35068
rect 9824 35028 9830 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 10778 35028 10784 35080
rect 10836 35028 10842 35080
rect 11054 35028 11060 35080
rect 11112 35028 11118 35080
rect 11793 35071 11851 35077
rect 11793 35037 11805 35071
rect 11839 35037 11851 35071
rect 12066 35068 12072 35080
rect 12027 35040 12072 35068
rect 11793 35031 11851 35037
rect 2332 34972 2728 35000
rect 4338 34960 4344 35012
rect 4396 34960 4402 35012
rect 4614 34960 4620 35012
rect 4672 35000 4678 35012
rect 4709 35003 4767 35009
rect 4709 35000 4721 35003
rect 4672 34972 4721 35000
rect 4672 34960 4678 34972
rect 4709 34969 4721 34972
rect 4755 34969 4767 35003
rect 5258 35000 5264 35012
rect 4709 34963 4767 34969
rect 5000 34972 5264 35000
rect 3326 34892 3332 34944
rect 3384 34932 3390 34944
rect 3786 34932 3792 34944
rect 3384 34904 3792 34932
rect 3384 34892 3390 34904
rect 3786 34892 3792 34904
rect 3844 34932 3850 34944
rect 3973 34935 4031 34941
rect 3973 34932 3985 34935
rect 3844 34904 3985 34932
rect 3844 34892 3850 34904
rect 3973 34901 3985 34904
rect 4019 34901 4031 34935
rect 3973 34895 4031 34901
rect 4430 34892 4436 34944
rect 4488 34932 4494 34944
rect 5000 34932 5028 34972
rect 5258 34960 5264 34972
rect 5316 34960 5322 35012
rect 7558 35000 7564 35012
rect 5368 34972 7564 35000
rect 4488 34904 5028 34932
rect 5077 34935 5135 34941
rect 4488 34892 4494 34904
rect 5077 34901 5089 34935
rect 5123 34932 5135 34935
rect 5166 34932 5172 34944
rect 5123 34904 5172 34932
rect 5123 34901 5135 34904
rect 5077 34895 5135 34901
rect 5166 34892 5172 34904
rect 5224 34932 5230 34944
rect 5368 34932 5396 34972
rect 7558 34960 7564 34972
rect 7616 34960 7622 35012
rect 11808 35000 11836 35031
rect 12066 35028 12072 35040
rect 12124 35028 12130 35080
rect 14093 35071 14151 35077
rect 14093 35037 14105 35071
rect 14139 35037 14151 35071
rect 14093 35031 14151 35037
rect 14367 35071 14425 35077
rect 14367 35037 14379 35071
rect 14413 35068 14425 35071
rect 14413 35040 15608 35068
rect 14413 35037 14425 35040
rect 14367 35031 14425 35037
rect 14108 35000 14136 35031
rect 14182 35000 14188 35012
rect 11808 34972 14188 35000
rect 14182 34960 14188 34972
rect 14240 34960 14246 35012
rect 5224 34904 5396 34932
rect 5224 34892 5230 34904
rect 5810 34892 5816 34944
rect 5868 34932 5874 34944
rect 14382 34932 14410 35031
rect 5868 34904 14410 34932
rect 5868 34892 5874 34904
rect 14458 34892 14464 34944
rect 14516 34932 14522 34944
rect 15105 34935 15163 34941
rect 15105 34932 15117 34935
rect 14516 34904 15117 34932
rect 14516 34892 14522 34904
rect 15105 34901 15117 34904
rect 15151 34901 15163 34935
rect 15580 34932 15608 35040
rect 15915 35041 15973 35047
rect 15915 35007 15927 35041
rect 15961 35038 15973 35041
rect 15961 35007 15974 35038
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 18141 35071 18199 35077
rect 18141 35068 18153 35071
rect 18012 35040 18153 35068
rect 18012 35028 18018 35040
rect 18141 35037 18153 35040
rect 18187 35037 18199 35071
rect 18141 35031 18199 35037
rect 18230 35028 18236 35080
rect 18288 35068 18294 35080
rect 19334 35068 19340 35080
rect 18288 35040 19340 35068
rect 18288 35028 18294 35040
rect 19334 35028 19340 35040
rect 19392 35068 19398 35080
rect 19705 35071 19763 35077
rect 19705 35068 19717 35071
rect 19392 35040 19717 35068
rect 19392 35028 19398 35040
rect 19705 35037 19717 35040
rect 19751 35037 19763 35071
rect 20073 35071 20131 35077
rect 20073 35068 20085 35071
rect 19705 35031 19763 35037
rect 19996 35040 20085 35068
rect 15915 35001 15974 35007
rect 15946 35000 15974 35001
rect 16390 35000 16396 35012
rect 15946 34972 16396 35000
rect 16390 34960 16396 34972
rect 16448 34960 16454 35012
rect 19242 34960 19248 35012
rect 19300 34960 19306 35012
rect 19426 34960 19432 35012
rect 19484 35000 19490 35012
rect 19996 35000 20024 35040
rect 20073 35037 20085 35040
rect 20119 35037 20131 35071
rect 20993 35071 21051 35077
rect 20993 35068 21005 35071
rect 20073 35031 20131 35037
rect 20456 35040 21005 35068
rect 19484 34972 20024 35000
rect 19484 34960 19490 34972
rect 19260 34932 19288 34960
rect 15580 34904 19288 34932
rect 19521 34935 19579 34941
rect 15105 34895 15163 34901
rect 19521 34901 19533 34935
rect 19567 34932 19579 34935
rect 19610 34932 19616 34944
rect 19567 34904 19616 34932
rect 19567 34901 19579 34904
rect 19521 34895 19579 34901
rect 19610 34892 19616 34904
rect 19668 34892 19674 34944
rect 19889 34935 19947 34941
rect 19889 34901 19901 34935
rect 19935 34932 19947 34935
rect 20456 34932 20484 35040
rect 20993 35037 21005 35040
rect 21039 35037 21051 35071
rect 22066 35068 22094 35108
rect 22278 35096 22284 35148
rect 22336 35136 22342 35148
rect 22646 35136 22652 35148
rect 22336 35108 22652 35136
rect 22336 35096 22342 35108
rect 22646 35096 22652 35108
rect 22704 35096 22710 35148
rect 22756 35108 23796 35136
rect 22756 35068 22784 35108
rect 22066 35040 22784 35068
rect 20993 35031 21051 35037
rect 23382 35028 23388 35080
rect 23440 35028 23446 35080
rect 23661 35071 23719 35077
rect 23661 35037 23673 35071
rect 23707 35037 23719 35071
rect 23661 35031 23719 35037
rect 20622 34960 20628 35012
rect 20680 35000 20686 35012
rect 23676 35000 23704 35031
rect 20680 34972 23704 35000
rect 23768 35000 23796 35108
rect 23952 35077 23980 35176
rect 23937 35071 23995 35077
rect 23937 35037 23949 35071
rect 23983 35037 23995 35071
rect 23937 35031 23995 35037
rect 24210 35000 24216 35012
rect 23768 34972 24216 35000
rect 20680 34960 20686 34972
rect 24210 34960 24216 34972
rect 24268 34960 24274 35012
rect 19935 34904 20484 34932
rect 19935 34901 19947 34904
rect 19889 34895 19947 34901
rect 23474 34892 23480 34944
rect 23532 34892 23538 34944
rect 24121 34935 24179 34941
rect 24121 34901 24133 34935
rect 24167 34932 24179 34935
rect 25222 34932 25228 34944
rect 24167 34904 25228 34932
rect 24167 34901 24179 34904
rect 24121 34895 24179 34901
rect 25222 34892 25228 34904
rect 25280 34892 25286 34944
rect 1104 34842 25000 34864
rect 1104 34790 6884 34842
rect 6936 34790 6948 34842
rect 7000 34790 7012 34842
rect 7064 34790 7076 34842
rect 7128 34790 7140 34842
rect 7192 34790 12818 34842
rect 12870 34790 12882 34842
rect 12934 34790 12946 34842
rect 12998 34790 13010 34842
rect 13062 34790 13074 34842
rect 13126 34790 18752 34842
rect 18804 34790 18816 34842
rect 18868 34790 18880 34842
rect 18932 34790 18944 34842
rect 18996 34790 19008 34842
rect 19060 34790 24686 34842
rect 24738 34790 24750 34842
rect 24802 34790 24814 34842
rect 24866 34790 24878 34842
rect 24930 34790 24942 34842
rect 24994 34790 25000 34842
rect 1104 34768 25000 34790
rect 2130 34688 2136 34740
rect 2188 34728 2194 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 2188 34700 2421 34728
rect 2188 34688 2194 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 2409 34691 2467 34697
rect 2590 34688 2596 34740
rect 2648 34728 2654 34740
rect 2774 34728 2780 34740
rect 2648 34700 2780 34728
rect 2648 34688 2654 34700
rect 2774 34688 2780 34700
rect 2832 34688 2838 34740
rect 3068 34700 4292 34728
rect 3068 34669 3096 34700
rect 3053 34663 3111 34669
rect 3053 34629 3065 34663
rect 3099 34629 3111 34663
rect 3053 34623 3111 34629
rect 3602 34620 3608 34672
rect 3660 34660 3666 34672
rect 3970 34660 3976 34672
rect 3660 34632 3976 34660
rect 3660 34620 3666 34632
rect 3970 34620 3976 34632
rect 4028 34620 4034 34672
rect 4264 34660 4292 34700
rect 4338 34688 4344 34740
rect 4396 34728 4402 34740
rect 4525 34731 4583 34737
rect 4525 34728 4537 34731
rect 4396 34700 4537 34728
rect 4396 34688 4402 34700
rect 4525 34697 4537 34700
rect 4571 34697 4583 34731
rect 4525 34691 4583 34697
rect 4614 34688 4620 34740
rect 4672 34728 4678 34740
rect 4672 34700 8340 34728
rect 4672 34688 4678 34700
rect 8312 34660 8340 34700
rect 9030 34688 9036 34740
rect 9088 34688 9094 34740
rect 14182 34728 14188 34740
rect 9140 34700 14188 34728
rect 9140 34660 9168 34700
rect 14182 34688 14188 34700
rect 14240 34688 14246 34740
rect 15197 34731 15255 34737
rect 15197 34697 15209 34731
rect 15243 34728 15255 34731
rect 15286 34728 15292 34740
rect 15243 34700 15292 34728
rect 15243 34697 15255 34700
rect 15197 34691 15255 34697
rect 15286 34688 15292 34700
rect 15344 34688 15350 34740
rect 15378 34688 15384 34740
rect 15436 34728 15442 34740
rect 16945 34731 17003 34737
rect 16945 34728 16957 34731
rect 15436 34700 16957 34728
rect 15436 34688 15442 34700
rect 16945 34697 16957 34700
rect 16991 34697 17003 34731
rect 16945 34691 17003 34697
rect 18785 34731 18843 34737
rect 18785 34697 18797 34731
rect 18831 34728 18843 34731
rect 19426 34728 19432 34740
rect 18831 34700 19432 34728
rect 18831 34697 18843 34700
rect 18785 34691 18843 34697
rect 19426 34688 19432 34700
rect 19484 34688 19490 34740
rect 21453 34731 21511 34737
rect 19536 34700 21128 34728
rect 4264 34632 8248 34660
rect 8312 34632 9168 34660
rect 1671 34595 1729 34601
rect 1671 34561 1683 34595
rect 1717 34592 1729 34595
rect 2406 34592 2412 34604
rect 1717 34564 2412 34592
rect 1717 34561 1729 34564
rect 1671 34555 1729 34561
rect 2406 34552 2412 34564
rect 2464 34552 2470 34604
rect 2774 34552 2780 34604
rect 2832 34552 2838 34604
rect 3326 34552 3332 34604
rect 3384 34592 3390 34604
rect 3513 34595 3571 34601
rect 3513 34592 3525 34595
rect 3384 34564 3525 34592
rect 3384 34552 3390 34564
rect 3513 34561 3525 34564
rect 3559 34561 3571 34595
rect 3513 34555 3571 34561
rect 3787 34595 3845 34601
rect 3787 34561 3799 34595
rect 3833 34592 3845 34595
rect 3988 34592 4016 34620
rect 3833 34564 4016 34592
rect 3833 34561 3845 34564
rect 3787 34555 3845 34561
rect 4154 34552 4160 34604
rect 4212 34592 4218 34604
rect 4893 34595 4951 34601
rect 4893 34592 4905 34595
rect 4212 34564 4905 34592
rect 4212 34552 4218 34564
rect 4893 34561 4905 34564
rect 4939 34561 4951 34595
rect 4893 34555 4951 34561
rect 5534 34552 5540 34604
rect 5592 34592 5598 34604
rect 6638 34601 6644 34604
rect 6607 34595 6644 34601
rect 6607 34592 6619 34595
rect 5592 34564 6619 34592
rect 5592 34552 5598 34564
rect 6607 34561 6619 34564
rect 6607 34555 6644 34561
rect 6638 34552 6644 34555
rect 6696 34552 6702 34604
rect 8220 34592 8248 34632
rect 9674 34620 9680 34672
rect 9732 34660 9738 34672
rect 9732 34632 11928 34660
rect 9732 34620 9738 34632
rect 8478 34592 8484 34604
rect 8220 34564 8484 34592
rect 8478 34552 8484 34564
rect 8536 34552 8542 34604
rect 8757 34595 8815 34601
rect 8757 34561 8769 34595
rect 8803 34592 8815 34595
rect 9309 34595 9367 34601
rect 9309 34592 9321 34595
rect 8803 34564 9321 34592
rect 8803 34561 8815 34564
rect 8757 34555 8815 34561
rect 9309 34561 9321 34564
rect 9355 34561 9367 34595
rect 9309 34555 9367 34561
rect 1394 34484 1400 34536
rect 1452 34484 1458 34536
rect 5077 34527 5135 34533
rect 5077 34493 5089 34527
rect 5123 34524 5135 34527
rect 5902 34524 5908 34536
rect 5123 34496 5908 34524
rect 5123 34493 5135 34496
rect 5077 34487 5135 34493
rect 5902 34484 5908 34496
rect 5960 34484 5966 34536
rect 6178 34484 6184 34536
rect 6236 34524 6242 34536
rect 6365 34527 6423 34533
rect 6365 34524 6377 34527
rect 6236 34496 6377 34524
rect 6236 34484 6242 34496
rect 6365 34493 6377 34496
rect 6411 34493 6423 34527
rect 9033 34527 9091 34533
rect 9033 34524 9045 34527
rect 6365 34487 6423 34493
rect 8772 34496 9045 34524
rect 1762 34348 1768 34400
rect 1820 34388 1826 34400
rect 5166 34388 5172 34400
rect 1820 34360 5172 34388
rect 1820 34348 1826 34360
rect 5166 34348 5172 34360
rect 5224 34348 5230 34400
rect 7374 34348 7380 34400
rect 7432 34348 7438 34400
rect 8772 34388 8800 34496
rect 9033 34493 9045 34496
rect 9079 34493 9091 34527
rect 9324 34524 9352 34555
rect 9490 34552 9496 34604
rect 9548 34552 9554 34604
rect 9582 34552 9588 34604
rect 9640 34552 9646 34604
rect 10060 34601 10088 34632
rect 10045 34595 10103 34601
rect 10045 34561 10057 34595
rect 10091 34561 10103 34595
rect 10045 34555 10103 34561
rect 10287 34595 10345 34601
rect 10287 34561 10299 34595
rect 10333 34592 10345 34595
rect 10686 34592 10692 34604
rect 10333 34564 10692 34592
rect 10333 34561 10345 34564
rect 10287 34555 10345 34561
rect 10686 34552 10692 34564
rect 10744 34552 10750 34604
rect 11900 34536 11928 34632
rect 14568 34632 15056 34660
rect 14459 34605 14517 34611
rect 14459 34571 14471 34605
rect 14505 34592 14517 34605
rect 14568 34592 14596 34632
rect 15028 34604 15056 34632
rect 16666 34620 16672 34672
rect 16724 34620 16730 34672
rect 16758 34620 16764 34672
rect 16816 34660 16822 34672
rect 16816 34632 16988 34660
rect 16816 34620 16822 34632
rect 16670 34617 16728 34620
rect 14505 34571 14596 34592
rect 14459 34565 14596 34571
rect 14474 34564 14596 34565
rect 14826 34552 14832 34604
rect 14884 34552 14890 34604
rect 15010 34552 15016 34604
rect 15068 34552 15074 34604
rect 16670 34583 16682 34617
rect 16716 34583 16728 34617
rect 16670 34577 16728 34583
rect 16960 34590 16988 34632
rect 17126 34620 17132 34672
rect 17184 34620 17190 34672
rect 19334 34669 19340 34672
rect 19328 34660 19340 34669
rect 17880 34632 19104 34660
rect 19295 34632 19340 34660
rect 17037 34595 17095 34601
rect 17037 34590 17049 34595
rect 16960 34562 17049 34590
rect 17037 34561 17049 34562
rect 17083 34561 17095 34595
rect 17144 34592 17172 34620
rect 17880 34604 17908 34632
rect 17313 34595 17371 34601
rect 17313 34592 17325 34595
rect 17144 34564 17325 34592
rect 17037 34555 17095 34561
rect 17313 34561 17325 34564
rect 17359 34561 17371 34595
rect 17313 34555 17371 34561
rect 17494 34552 17500 34604
rect 17552 34552 17558 34604
rect 17862 34552 17868 34604
rect 17920 34552 17926 34604
rect 18966 34552 18972 34604
rect 19024 34552 19030 34604
rect 19076 34592 19104 34632
rect 19328 34623 19340 34632
rect 19334 34620 19340 34623
rect 19392 34620 19398 34672
rect 19536 34592 19564 34700
rect 19610 34620 19616 34672
rect 19668 34620 19674 34672
rect 20438 34620 20444 34672
rect 20496 34660 20502 34672
rect 21100 34660 21128 34700
rect 21453 34697 21465 34731
rect 21499 34728 21511 34731
rect 21499 34700 22784 34728
rect 21499 34697 21511 34700
rect 21453 34691 21511 34697
rect 20496 34632 21036 34660
rect 21100 34632 21680 34660
rect 20496 34620 20502 34632
rect 19076 34564 19564 34592
rect 19628 34592 19656 34620
rect 21008 34601 21036 34632
rect 21652 34601 21680 34632
rect 22079 34625 22137 34631
rect 20533 34595 20591 34601
rect 20533 34592 20545 34595
rect 19628 34564 20545 34592
rect 20533 34561 20545 34564
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34561 21051 34595
rect 20993 34555 21051 34561
rect 21637 34595 21695 34601
rect 21637 34561 21649 34595
rect 21683 34561 21695 34595
rect 22079 34591 22091 34625
rect 22125 34622 22137 34625
rect 22125 34592 22140 34622
rect 22186 34592 22192 34604
rect 22125 34591 22192 34592
rect 22079 34585 22192 34591
rect 22112 34564 22192 34585
rect 21637 34555 21695 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 22756 34592 22784 34700
rect 23290 34688 23296 34740
rect 23348 34728 23354 34740
rect 23348 34700 23520 34728
rect 23348 34688 23354 34700
rect 23492 34660 23520 34700
rect 23658 34688 23664 34740
rect 23716 34688 23722 34740
rect 23750 34688 23756 34740
rect 23808 34728 23814 34740
rect 23808 34700 24164 34728
rect 23808 34688 23814 34700
rect 23492 34632 23888 34660
rect 23860 34601 23888 34632
rect 23934 34620 23940 34672
rect 23992 34620 23998 34672
rect 24136 34669 24164 34700
rect 24121 34663 24179 34669
rect 24121 34629 24133 34663
rect 24167 34629 24179 34663
rect 24121 34623 24179 34629
rect 23385 34595 23443 34601
rect 23385 34592 23397 34595
rect 22756 34564 23397 34592
rect 23385 34561 23397 34564
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 23845 34595 23903 34601
rect 23845 34561 23857 34595
rect 23891 34561 23903 34595
rect 23845 34555 23903 34561
rect 9324 34516 9444 34524
rect 9600 34516 9812 34524
rect 9324 34496 9812 34516
rect 9033 34487 9091 34493
rect 9416 34488 9628 34496
rect 8849 34459 8907 34465
rect 8849 34425 8861 34459
rect 8895 34456 8907 34459
rect 9677 34459 9735 34465
rect 9677 34456 9689 34459
rect 8895 34428 9689 34456
rect 8895 34425 8907 34428
rect 8849 34419 8907 34425
rect 9677 34425 9689 34428
rect 9723 34425 9735 34459
rect 9677 34419 9735 34425
rect 9784 34400 9812 34496
rect 11882 34484 11888 34536
rect 11940 34484 11946 34536
rect 13906 34484 13912 34536
rect 13964 34524 13970 34536
rect 14185 34527 14243 34533
rect 14185 34524 14197 34527
rect 13964 34496 14197 34524
rect 13964 34484 13970 34496
rect 14185 34493 14197 34496
rect 14231 34493 14243 34527
rect 14185 34487 14243 34493
rect 11698 34416 11704 34468
rect 11756 34456 11762 34468
rect 11756 34428 13676 34456
rect 11756 34416 11762 34428
rect 9401 34391 9459 34397
rect 9401 34388 9413 34391
rect 8772 34360 9413 34388
rect 9401 34357 9413 34360
rect 9447 34357 9459 34391
rect 9401 34351 9459 34357
rect 9766 34348 9772 34400
rect 9824 34348 9830 34400
rect 11054 34348 11060 34400
rect 11112 34348 11118 34400
rect 13648 34388 13676 34428
rect 14844 34388 14872 34552
rect 16945 34527 17003 34533
rect 16945 34493 16957 34527
rect 16991 34524 17003 34527
rect 17405 34527 17463 34533
rect 17405 34524 17417 34527
rect 16991 34496 17417 34524
rect 16991 34493 17003 34496
rect 16945 34487 17003 34493
rect 17405 34493 17417 34496
rect 17451 34493 17463 34527
rect 19058 34524 19064 34536
rect 17405 34487 17463 34493
rect 18156 34496 19064 34524
rect 16761 34459 16819 34465
rect 16761 34425 16773 34459
rect 16807 34456 16819 34459
rect 17129 34459 17187 34465
rect 17129 34456 17141 34459
rect 16807 34428 17141 34456
rect 16807 34425 16819 34428
rect 16761 34419 16819 34425
rect 17129 34425 17141 34428
rect 17175 34425 17187 34459
rect 17129 34419 17187 34425
rect 17218 34416 17224 34468
rect 17276 34456 17282 34468
rect 18156 34456 18184 34496
rect 19058 34484 19064 34496
rect 19116 34484 19122 34536
rect 20625 34527 20683 34533
rect 20625 34493 20637 34527
rect 20671 34524 20683 34527
rect 21082 34524 21088 34536
rect 20671 34496 21088 34524
rect 20671 34493 20683 34496
rect 20625 34487 20683 34493
rect 21082 34484 21088 34496
rect 21140 34484 21146 34536
rect 21821 34527 21879 34533
rect 21821 34524 21833 34527
rect 21192 34496 21833 34524
rect 21192 34456 21220 34496
rect 21821 34493 21833 34496
rect 21867 34493 21879 34527
rect 23952 34524 23980 34620
rect 21821 34487 21879 34493
rect 23216 34496 23980 34524
rect 23216 34465 23244 34496
rect 24394 34484 24400 34536
rect 24452 34484 24458 34536
rect 17276 34428 18184 34456
rect 19996 34428 21220 34456
rect 23201 34459 23259 34465
rect 17276 34416 17282 34428
rect 19996 34400 20024 34428
rect 23201 34425 23213 34459
rect 23247 34425 23259 34459
rect 23201 34419 23259 34425
rect 13648 34360 14872 34388
rect 15010 34348 15016 34400
rect 15068 34388 15074 34400
rect 19794 34388 19800 34400
rect 15068 34360 19800 34388
rect 15068 34348 15074 34360
rect 19794 34348 19800 34360
rect 19852 34348 19858 34400
rect 19978 34348 19984 34400
rect 20036 34348 20042 34400
rect 20438 34348 20444 34400
rect 20496 34348 20502 34400
rect 20806 34348 20812 34400
rect 20864 34348 20870 34400
rect 22833 34391 22891 34397
rect 22833 34357 22845 34391
rect 22879 34388 22891 34391
rect 23106 34388 23112 34400
rect 22879 34360 23112 34388
rect 22879 34357 22891 34360
rect 22833 34351 22891 34357
rect 23106 34348 23112 34360
rect 23164 34348 23170 34400
rect 1104 34298 24840 34320
rect 1104 34246 3917 34298
rect 3969 34246 3981 34298
rect 4033 34246 4045 34298
rect 4097 34246 4109 34298
rect 4161 34246 4173 34298
rect 4225 34246 9851 34298
rect 9903 34246 9915 34298
rect 9967 34246 9979 34298
rect 10031 34246 10043 34298
rect 10095 34246 10107 34298
rect 10159 34246 15785 34298
rect 15837 34246 15849 34298
rect 15901 34246 15913 34298
rect 15965 34246 15977 34298
rect 16029 34246 16041 34298
rect 16093 34246 21719 34298
rect 21771 34246 21783 34298
rect 21835 34246 21847 34298
rect 21899 34246 21911 34298
rect 21963 34246 21975 34298
rect 22027 34246 24840 34298
rect 1104 34224 24840 34246
rect 198 34144 204 34196
rect 256 34184 262 34196
rect 1762 34184 1768 34196
rect 256 34156 1768 34184
rect 256 34144 262 34156
rect 1762 34144 1768 34156
rect 1820 34144 1826 34196
rect 2958 34144 2964 34196
rect 3016 34144 3022 34196
rect 5534 34184 5540 34196
rect 3068 34156 5540 34184
rect 2976 34048 3004 34144
rect 3068 34057 3096 34156
rect 5534 34144 5540 34156
rect 5592 34144 5598 34196
rect 9398 34184 9404 34196
rect 7024 34156 9404 34184
rect 2700 34020 3004 34048
rect 3053 34051 3111 34057
rect 750 33940 756 33992
rect 808 33980 814 33992
rect 1394 33980 1400 33992
rect 808 33952 1400 33980
rect 808 33940 814 33952
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 1671 33983 1729 33989
rect 1671 33949 1683 33983
rect 1717 33980 1729 33983
rect 2700 33980 2728 34020
rect 3053 34017 3065 34051
rect 3099 34017 3111 34051
rect 3053 34011 3111 34017
rect 6454 34008 6460 34060
rect 6512 34048 6518 34060
rect 6822 34048 6828 34060
rect 6512 34020 6828 34048
rect 6512 34008 6518 34020
rect 6822 34008 6828 34020
rect 6880 34008 6886 34060
rect 7024 34057 7052 34156
rect 9398 34144 9404 34156
rect 9456 34184 9462 34196
rect 9456 34156 9674 34184
rect 9456 34144 9462 34156
rect 7374 34076 7380 34128
rect 7432 34116 7438 34128
rect 7469 34119 7527 34125
rect 7469 34116 7481 34119
rect 7432 34088 7481 34116
rect 7432 34076 7438 34088
rect 7469 34085 7481 34088
rect 7515 34085 7527 34119
rect 7469 34079 7527 34085
rect 8478 34076 8484 34128
rect 8536 34116 8542 34128
rect 9646 34116 9674 34156
rect 9766 34144 9772 34196
rect 9824 34184 9830 34196
rect 9953 34187 10011 34193
rect 9953 34184 9965 34187
rect 9824 34156 9965 34184
rect 9824 34144 9830 34156
rect 9953 34153 9965 34156
rect 9999 34153 10011 34187
rect 16206 34184 16212 34196
rect 9953 34147 10011 34153
rect 10796 34156 16212 34184
rect 10796 34128 10824 34156
rect 16206 34144 16212 34156
rect 16264 34144 16270 34196
rect 17313 34187 17371 34193
rect 17313 34153 17325 34187
rect 17359 34184 17371 34187
rect 17494 34184 17500 34196
rect 17359 34156 17500 34184
rect 17359 34153 17371 34156
rect 17313 34147 17371 34153
rect 17494 34144 17500 34156
rect 17552 34144 17558 34196
rect 20530 34184 20536 34196
rect 17604 34156 20536 34184
rect 10686 34116 10692 34128
rect 8536 34088 8800 34116
rect 9646 34088 10692 34116
rect 8536 34076 8542 34088
rect 7009 34051 7067 34057
rect 7009 34017 7021 34051
rect 7055 34017 7067 34051
rect 7745 34051 7803 34057
rect 7745 34048 7757 34051
rect 7009 34011 7067 34017
rect 7114 34020 7757 34048
rect 1717 33952 2728 33980
rect 1717 33949 1729 33952
rect 1671 33943 1729 33949
rect 2774 33940 2780 33992
rect 2832 33940 2838 33992
rect 3789 33983 3847 33989
rect 3789 33980 3801 33983
rect 2976 33952 3801 33980
rect 1302 33872 1308 33924
rect 1360 33912 1366 33924
rect 2976 33912 3004 33952
rect 3789 33949 3801 33952
rect 3835 33949 3847 33983
rect 3789 33943 3847 33949
rect 4525 33983 4583 33989
rect 4525 33949 4537 33983
rect 4571 33949 4583 33983
rect 4525 33943 4583 33949
rect 4767 33983 4825 33989
rect 4767 33949 4779 33983
rect 4813 33980 4825 33983
rect 5258 33980 5264 33992
rect 4813 33952 5264 33980
rect 4813 33949 4825 33952
rect 4767 33943 4825 33949
rect 1360 33884 3004 33912
rect 1360 33872 1366 33884
rect 4062 33872 4068 33924
rect 4120 33872 4126 33924
rect 4540 33912 4568 33943
rect 5258 33940 5264 33952
rect 5316 33980 5322 33992
rect 6362 33980 6368 33992
rect 5316 33952 6368 33980
rect 5316 33940 5322 33952
rect 6362 33940 6368 33952
rect 6420 33940 6426 33992
rect 7114 33980 7142 34020
rect 7745 34017 7757 34020
rect 7791 34017 7803 34051
rect 7745 34011 7803 34017
rect 7898 34020 8616 34048
rect 7898 33989 7926 34020
rect 6472 33952 7142 33980
rect 7883 33983 7941 33989
rect 4890 33912 4896 33924
rect 4540 33884 4896 33912
rect 4890 33872 4896 33884
rect 4948 33912 4954 33924
rect 6178 33912 6184 33924
rect 4948 33884 6184 33912
rect 4948 33872 4954 33884
rect 6178 33872 6184 33884
rect 6236 33872 6242 33924
rect 6472 33856 6500 33952
rect 7883 33949 7895 33983
rect 7929 33949 7941 33983
rect 7883 33943 7941 33949
rect 8018 33940 8024 33992
rect 8076 33940 8082 33992
rect 8588 33912 8616 34020
rect 8772 33980 8800 34088
rect 10686 34076 10692 34088
rect 10744 34076 10750 34128
rect 10778 34076 10784 34128
rect 10836 34076 10842 34128
rect 13541 34119 13599 34125
rect 13541 34085 13553 34119
rect 13587 34116 13599 34119
rect 13722 34116 13728 34128
rect 13587 34088 13728 34116
rect 13587 34085 13599 34088
rect 13541 34079 13599 34085
rect 13722 34076 13728 34088
rect 13780 34076 13786 34128
rect 16758 34076 16764 34128
rect 16816 34116 16822 34128
rect 17604 34116 17632 34156
rect 20530 34144 20536 34156
rect 20588 34144 20594 34196
rect 20806 34144 20812 34196
rect 20864 34144 20870 34196
rect 21082 34144 21088 34196
rect 21140 34144 21146 34196
rect 22373 34187 22431 34193
rect 22373 34153 22385 34187
rect 22419 34184 22431 34187
rect 23382 34184 23388 34196
rect 22419 34156 23388 34184
rect 22419 34153 22431 34156
rect 22373 34147 22431 34153
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 16816 34088 17632 34116
rect 17681 34119 17739 34125
rect 16816 34076 16822 34088
rect 17681 34085 17693 34119
rect 17727 34085 17739 34119
rect 17681 34079 17739 34085
rect 20625 34119 20683 34125
rect 20625 34085 20637 34119
rect 20671 34085 20683 34119
rect 20824 34116 20852 34144
rect 23109 34119 23167 34125
rect 20824 34088 21588 34116
rect 20625 34079 20683 34085
rect 8846 34008 8852 34060
rect 8904 34048 8910 34060
rect 8941 34051 8999 34057
rect 8941 34048 8953 34051
rect 8904 34020 8953 34048
rect 8904 34008 8910 34020
rect 8941 34017 8953 34020
rect 8987 34017 8999 34051
rect 11606 34048 11612 34060
rect 8941 34011 8999 34017
rect 10428 34020 11612 34048
rect 9183 33983 9241 33989
rect 9183 33980 9195 33983
rect 8772 33952 9195 33980
rect 9183 33949 9195 33952
rect 9229 33949 9241 33983
rect 10428 33980 10456 34020
rect 11606 34008 11612 34020
rect 11664 34008 11670 34060
rect 11882 34008 11888 34060
rect 11940 34048 11946 34060
rect 12526 34048 12532 34060
rect 11940 34020 12532 34048
rect 11940 34008 11946 34020
rect 12526 34008 12532 34020
rect 12584 34008 12590 34060
rect 15194 34008 15200 34060
rect 15252 34048 15258 34060
rect 15470 34048 15476 34060
rect 15252 34020 15476 34048
rect 15252 34008 15258 34020
rect 15470 34008 15476 34020
rect 15528 34048 15534 34060
rect 15933 34051 15991 34057
rect 15933 34048 15945 34051
rect 15528 34020 15945 34048
rect 15528 34008 15534 34020
rect 15933 34017 15945 34020
rect 15979 34017 15991 34051
rect 15933 34011 15991 34017
rect 17310 34008 17316 34060
rect 17368 34048 17374 34060
rect 17696 34048 17724 34079
rect 17368 34020 17632 34048
rect 17696 34020 18184 34048
rect 17368 34008 17374 34020
rect 9183 33943 9241 33949
rect 9324 33952 10456 33980
rect 12803 33983 12861 33989
rect 9324 33912 9352 33952
rect 12803 33949 12815 33983
rect 12849 33980 12861 33983
rect 13538 33980 13544 33992
rect 12849 33952 13544 33980
rect 12849 33949 12861 33952
rect 12803 33943 12861 33949
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 13906 33940 13912 33992
rect 13964 33980 13970 33992
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 13964 33952 14105 33980
rect 13964 33940 13970 33952
rect 14093 33949 14105 33952
rect 14139 33949 14151 33983
rect 14351 33983 14409 33989
rect 14351 33980 14363 33983
rect 14093 33943 14151 33949
rect 14292 33952 14363 33980
rect 8588 33884 8800 33912
rect 290 33804 296 33856
rect 348 33844 354 33856
rect 566 33844 572 33856
rect 348 33816 572 33844
rect 348 33804 354 33816
rect 566 33804 572 33816
rect 624 33804 630 33856
rect 1762 33804 1768 33856
rect 1820 33844 1826 33856
rect 2409 33847 2467 33853
rect 2409 33844 2421 33847
rect 1820 33816 2421 33844
rect 1820 33804 1826 33816
rect 2409 33813 2421 33816
rect 2455 33813 2467 33847
rect 2409 33807 2467 33813
rect 5534 33804 5540 33856
rect 5592 33804 5598 33856
rect 6454 33804 6460 33856
rect 6512 33804 6518 33856
rect 8662 33804 8668 33856
rect 8720 33804 8726 33856
rect 8772 33844 8800 33884
rect 9048 33884 9352 33912
rect 9048 33844 9076 33884
rect 9490 33872 9496 33924
rect 9548 33912 9554 33924
rect 12342 33912 12348 33924
rect 9548 33884 12348 33912
rect 9548 33872 9554 33884
rect 12342 33872 12348 33884
rect 12400 33872 12406 33924
rect 12618 33872 12624 33924
rect 12676 33912 12682 33924
rect 13998 33912 14004 33924
rect 12676 33884 14004 33912
rect 12676 33872 12682 33884
rect 13998 33872 14004 33884
rect 14056 33872 14062 33924
rect 14292 33912 14320 33952
rect 14351 33949 14363 33952
rect 14397 33980 14409 33983
rect 15378 33980 15384 33992
rect 14397 33952 15384 33980
rect 14397 33949 14409 33952
rect 14351 33943 14409 33949
rect 15378 33940 15384 33952
rect 15436 33940 15442 33992
rect 16206 33940 16212 33992
rect 16264 33980 16270 33992
rect 16850 33980 16856 33992
rect 16264 33952 16856 33980
rect 16264 33940 16270 33952
rect 16850 33940 16856 33952
rect 16908 33940 16914 33992
rect 17494 33940 17500 33992
rect 17552 33940 17558 33992
rect 17604 33980 17632 34020
rect 18156 33989 18184 34020
rect 17865 33983 17923 33989
rect 17865 33980 17877 33983
rect 17604 33952 17877 33980
rect 17865 33949 17877 33952
rect 17911 33949 17923 33983
rect 17865 33943 17923 33949
rect 18141 33983 18199 33989
rect 18141 33949 18153 33983
rect 18187 33949 18199 33983
rect 18141 33943 18199 33949
rect 19613 33983 19671 33989
rect 19613 33949 19625 33983
rect 19659 33949 19671 33983
rect 19613 33943 19671 33949
rect 14108 33884 14320 33912
rect 8772 33816 9076 33844
rect 9398 33804 9404 33856
rect 9456 33844 9462 33856
rect 14108 33844 14136 33884
rect 17034 33872 17040 33924
rect 17092 33912 17098 33924
rect 19518 33912 19524 33924
rect 17092 33884 19524 33912
rect 17092 33872 17098 33884
rect 19518 33872 19524 33884
rect 19576 33872 19582 33924
rect 19628 33912 19656 33943
rect 19794 33940 19800 33992
rect 19852 33980 19858 33992
rect 19887 33983 19945 33989
rect 19887 33980 19899 33983
rect 19852 33952 19899 33980
rect 19852 33940 19858 33952
rect 19887 33949 19899 33952
rect 19933 33949 19945 33983
rect 20640 33980 20668 34079
rect 21269 34051 21327 34057
rect 21269 34017 21281 34051
rect 21315 34048 21327 34051
rect 21453 34051 21511 34057
rect 21453 34048 21465 34051
rect 21315 34020 21465 34048
rect 21315 34017 21327 34020
rect 21269 34011 21327 34017
rect 21453 34017 21465 34020
rect 21499 34017 21511 34051
rect 21453 34011 21511 34017
rect 21560 33989 21588 34088
rect 23109 34085 23121 34119
rect 23155 34085 23167 34119
rect 23109 34079 23167 34085
rect 23124 34048 23152 34079
rect 23124 34020 23980 34048
rect 20993 33983 21051 33989
rect 20993 33980 21005 33983
rect 20640 33952 21005 33980
rect 19887 33943 19945 33949
rect 20993 33949 21005 33952
rect 21039 33980 21051 33983
rect 21361 33983 21419 33989
rect 21361 33980 21373 33983
rect 21039 33952 21373 33980
rect 21039 33949 21051 33952
rect 20993 33943 21051 33949
rect 21361 33949 21373 33952
rect 21407 33949 21419 33983
rect 21361 33943 21419 33949
rect 21545 33983 21603 33989
rect 21545 33949 21557 33983
rect 21591 33949 21603 33983
rect 21545 33943 21603 33949
rect 22554 33940 22560 33992
rect 22612 33940 22618 33992
rect 22830 33940 22836 33992
rect 22888 33940 22894 33992
rect 23293 33983 23351 33989
rect 23293 33980 23305 33983
rect 23124 33952 23305 33980
rect 19628 33884 19932 33912
rect 19904 33856 19932 33884
rect 9456 33816 14136 33844
rect 9456 33804 9462 33816
rect 14274 33804 14280 33856
rect 14332 33844 14338 33856
rect 15010 33844 15016 33856
rect 14332 33816 15016 33844
rect 14332 33804 14338 33816
rect 15010 33804 15016 33816
rect 15068 33804 15074 33856
rect 15102 33804 15108 33856
rect 15160 33804 15166 33856
rect 16942 33804 16948 33856
rect 17000 33804 17006 33856
rect 18230 33804 18236 33856
rect 18288 33804 18294 33856
rect 19886 33804 19892 33856
rect 19944 33804 19950 33856
rect 21269 33847 21327 33853
rect 21269 33813 21281 33847
rect 21315 33844 21327 33847
rect 21634 33844 21640 33856
rect 21315 33816 21640 33844
rect 21315 33813 21327 33816
rect 21269 33807 21327 33813
rect 21634 33804 21640 33816
rect 21692 33804 21698 33856
rect 22646 33804 22652 33856
rect 22704 33804 22710 33856
rect 23124 33844 23152 33952
rect 23293 33949 23305 33952
rect 23339 33949 23351 33983
rect 23293 33943 23351 33949
rect 23474 33940 23480 33992
rect 23532 33980 23538 33992
rect 23952 33989 23980 34020
rect 23569 33983 23627 33989
rect 23569 33980 23581 33983
rect 23532 33952 23581 33980
rect 23532 33940 23538 33952
rect 23569 33949 23581 33952
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 23845 33983 23903 33989
rect 23845 33949 23857 33983
rect 23891 33949 23903 33983
rect 23845 33943 23903 33949
rect 23937 33983 23995 33989
rect 23937 33949 23949 33983
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 23198 33872 23204 33924
rect 23256 33912 23262 33924
rect 23860 33912 23888 33943
rect 23256 33884 23888 33912
rect 23256 33872 23262 33884
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 23124 33816 23397 33844
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 23658 33804 23664 33856
rect 23716 33804 23722 33856
rect 24121 33847 24179 33853
rect 24121 33813 24133 33847
rect 24167 33844 24179 33847
rect 25222 33844 25228 33856
rect 24167 33816 25228 33844
rect 24167 33813 24179 33816
rect 24121 33807 24179 33813
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 1104 33754 25000 33776
rect 1104 33702 6884 33754
rect 6936 33702 6948 33754
rect 7000 33702 7012 33754
rect 7064 33702 7076 33754
rect 7128 33702 7140 33754
rect 7192 33702 12818 33754
rect 12870 33702 12882 33754
rect 12934 33702 12946 33754
rect 12998 33702 13010 33754
rect 13062 33702 13074 33754
rect 13126 33702 18752 33754
rect 18804 33702 18816 33754
rect 18868 33702 18880 33754
rect 18932 33702 18944 33754
rect 18996 33702 19008 33754
rect 19060 33702 24686 33754
rect 24738 33702 24750 33754
rect 24802 33702 24814 33754
rect 24866 33702 24878 33754
rect 24930 33702 24942 33754
rect 24994 33702 25000 33754
rect 1104 33680 25000 33702
rect 1210 33600 1216 33652
rect 1268 33640 1274 33652
rect 1268 33612 1716 33640
rect 1268 33600 1274 33612
rect 1688 33504 1716 33612
rect 2682 33600 2688 33652
rect 2740 33640 2746 33652
rect 2958 33640 2964 33652
rect 2740 33612 2964 33640
rect 2740 33600 2746 33612
rect 2958 33600 2964 33612
rect 3016 33640 3022 33652
rect 3786 33640 3792 33652
rect 3016 33612 3792 33640
rect 3016 33600 3022 33612
rect 3786 33600 3792 33612
rect 3844 33600 3850 33652
rect 5166 33600 5172 33652
rect 5224 33640 5230 33652
rect 7098 33640 7104 33652
rect 5224 33612 7104 33640
rect 5224 33600 5230 33612
rect 7098 33600 7104 33612
rect 7156 33600 7162 33652
rect 8662 33600 8668 33652
rect 8720 33600 8726 33652
rect 8849 33643 8907 33649
rect 8849 33609 8861 33643
rect 8895 33640 8907 33643
rect 9030 33640 9036 33652
rect 8895 33612 9036 33640
rect 8895 33609 8907 33612
rect 8849 33603 8907 33609
rect 9030 33600 9036 33612
rect 9088 33600 9094 33652
rect 9125 33643 9183 33649
rect 9125 33609 9137 33643
rect 9171 33640 9183 33643
rect 9582 33640 9588 33652
rect 9171 33612 9588 33640
rect 9171 33609 9183 33612
rect 9125 33603 9183 33609
rect 9582 33600 9588 33612
rect 9640 33600 9646 33652
rect 11606 33600 11612 33652
rect 11664 33640 11670 33652
rect 11790 33640 11796 33652
rect 11664 33612 11796 33640
rect 11664 33600 11670 33612
rect 11790 33600 11796 33612
rect 11848 33640 11854 33652
rect 12710 33640 12716 33652
rect 11848 33612 12716 33640
rect 11848 33600 11854 33612
rect 12710 33600 12716 33612
rect 12768 33600 12774 33652
rect 13722 33600 13728 33652
rect 13780 33600 13786 33652
rect 13998 33600 14004 33652
rect 14056 33640 14062 33652
rect 16758 33640 16764 33652
rect 14056 33612 16764 33640
rect 14056 33600 14062 33612
rect 3050 33532 3056 33584
rect 3108 33532 3114 33584
rect 3329 33575 3387 33581
rect 3329 33541 3341 33575
rect 3375 33572 3387 33575
rect 4157 33575 4215 33581
rect 3375 33544 4108 33572
rect 3375 33541 3387 33544
rect 3329 33535 3387 33541
rect 1747 33507 1805 33513
rect 1747 33504 1759 33507
rect 1688 33476 1759 33504
rect 1747 33473 1759 33476
rect 1793 33504 1805 33507
rect 3234 33504 3240 33516
rect 1793 33476 2268 33504
rect 1793 33473 1805 33476
rect 1747 33467 1805 33473
rect 1394 33396 1400 33448
rect 1452 33436 1458 33448
rect 1489 33439 1547 33445
rect 1489 33436 1501 33439
rect 1452 33408 1501 33436
rect 1452 33396 1458 33408
rect 1489 33405 1501 33408
rect 1535 33405 1547 33439
rect 2240 33436 2268 33476
rect 2424 33476 3240 33504
rect 2424 33436 2452 33476
rect 3234 33464 3240 33476
rect 3292 33464 3298 33516
rect 3418 33464 3424 33516
rect 3476 33464 3482 33516
rect 3786 33464 3792 33516
rect 3844 33464 3850 33516
rect 4080 33504 4108 33544
rect 4157 33541 4169 33575
rect 4203 33572 4215 33575
rect 4522 33572 4528 33584
rect 4203 33544 4528 33572
rect 4203 33541 4215 33544
rect 4157 33535 4215 33541
rect 4522 33532 4528 33544
rect 4580 33572 4586 33584
rect 5350 33572 5356 33584
rect 4580 33544 4752 33572
rect 4580 33532 4586 33544
rect 4614 33504 4620 33516
rect 4080 33476 4620 33504
rect 4614 33464 4620 33476
rect 4672 33464 4678 33516
rect 2240 33408 2452 33436
rect 2746 33408 2898 33436
rect 1489 33399 1547 33405
rect 2501 33371 2559 33377
rect 2501 33337 2513 33371
rect 2547 33368 2559 33371
rect 2746 33368 2774 33408
rect 2547 33340 2774 33368
rect 2547 33337 2559 33340
rect 2501 33331 2559 33337
rect 4338 33328 4344 33380
rect 4396 33328 4402 33380
rect 2406 33260 2412 33312
rect 2464 33300 2470 33312
rect 2682 33300 2688 33312
rect 2464 33272 2688 33300
rect 2464 33260 2470 33272
rect 2682 33260 2688 33272
rect 2740 33260 2746 33312
rect 4724 33300 4752 33544
rect 5184 33544 5356 33572
rect 5184 33543 5212 33544
rect 5151 33537 5212 33543
rect 4890 33464 4896 33516
rect 4948 33464 4954 33516
rect 5151 33503 5163 33537
rect 5197 33506 5212 33537
rect 5350 33532 5356 33544
rect 5408 33532 5414 33584
rect 5197 33503 5209 33506
rect 7282 33504 7288 33516
rect 5151 33497 5209 33503
rect 6932 33476 7288 33504
rect 6932 33448 6960 33476
rect 7282 33464 7288 33476
rect 7340 33464 7346 33516
rect 8110 33464 8116 33516
rect 8168 33464 8174 33516
rect 8680 33504 8708 33600
rect 10962 33572 10968 33584
rect 9692 33544 10968 33572
rect 9033 33507 9091 33513
rect 9033 33504 9045 33507
rect 8680 33476 9045 33504
rect 9033 33473 9045 33476
rect 9079 33473 9091 33507
rect 9033 33467 9091 33473
rect 9309 33507 9367 33513
rect 9309 33473 9321 33507
rect 9355 33473 9367 33507
rect 9692 33504 9720 33544
rect 10962 33532 10968 33544
rect 11020 33572 11026 33584
rect 11020 33544 12020 33572
rect 11020 33532 11026 33544
rect 9766 33513 9772 33516
rect 9309 33467 9367 33473
rect 9416 33476 9720 33504
rect 9751 33507 9772 33513
rect 6914 33396 6920 33448
rect 6972 33396 6978 33448
rect 7101 33439 7159 33445
rect 7101 33405 7113 33439
rect 7147 33405 7159 33439
rect 7101 33399 7159 33405
rect 5166 33300 5172 33312
rect 4724 33272 5172 33300
rect 5166 33260 5172 33272
rect 5224 33260 5230 33312
rect 5350 33260 5356 33312
rect 5408 33300 5414 33312
rect 5905 33303 5963 33309
rect 5905 33300 5917 33303
rect 5408 33272 5917 33300
rect 5408 33260 5414 33272
rect 5905 33269 5917 33272
rect 5951 33269 5963 33303
rect 7116 33300 7144 33399
rect 7190 33396 7196 33448
rect 7248 33436 7254 33448
rect 7837 33439 7895 33445
rect 7837 33436 7849 33439
rect 7248 33408 7849 33436
rect 7248 33396 7254 33408
rect 7837 33405 7849 33408
rect 7883 33405 7895 33439
rect 7837 33399 7895 33405
rect 7926 33396 7932 33448
rect 7984 33445 7990 33448
rect 7984 33439 8012 33445
rect 8000 33405 8012 33439
rect 7984 33399 8012 33405
rect 8757 33439 8815 33445
rect 8757 33405 8769 33439
rect 8803 33436 8815 33439
rect 9324 33436 9352 33467
rect 8803 33408 9352 33436
rect 8803 33405 8815 33408
rect 8757 33399 8815 33405
rect 7984 33396 7990 33399
rect 7374 33328 7380 33380
rect 7432 33368 7438 33380
rect 7561 33371 7619 33377
rect 7561 33368 7573 33371
rect 7432 33340 7573 33368
rect 7432 33328 7438 33340
rect 7561 33337 7573 33340
rect 7607 33337 7619 33371
rect 9416 33368 9444 33476
rect 9751 33473 9763 33507
rect 9751 33467 9772 33473
rect 9766 33464 9772 33467
rect 9824 33464 9830 33516
rect 9858 33464 9864 33516
rect 9916 33504 9922 33516
rect 11992 33513 12020 33544
rect 11977 33507 12035 33513
rect 9916 33476 11928 33504
rect 9916 33464 9922 33476
rect 9493 33439 9551 33445
rect 9493 33405 9505 33439
rect 9539 33405 9551 33439
rect 9493 33399 9551 33405
rect 7561 33331 7619 33337
rect 8588 33340 9444 33368
rect 8588 33300 8616 33340
rect 7116 33272 8616 33300
rect 9508 33300 9536 33399
rect 11054 33396 11060 33448
rect 11112 33436 11118 33448
rect 11793 33439 11851 33445
rect 11793 33436 11805 33439
rect 11112 33408 11805 33436
rect 11112 33396 11118 33408
rect 11793 33405 11805 33408
rect 11839 33405 11851 33439
rect 11900 33436 11928 33476
rect 11977 33473 11989 33507
rect 12023 33504 12035 33507
rect 12158 33504 12164 33516
rect 12023 33476 12164 33504
rect 12023 33473 12035 33476
rect 11977 33467 12035 33473
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 12710 33464 12716 33516
rect 12768 33464 12774 33516
rect 12830 33439 12888 33445
rect 12830 33436 12842 33439
rect 11900 33408 12842 33436
rect 11793 33399 11851 33405
rect 12830 33405 12842 33408
rect 12876 33405 12888 33439
rect 12830 33399 12888 33405
rect 12989 33439 13047 33445
rect 12989 33405 13001 33439
rect 13035 33436 13047 33439
rect 13740 33436 13768 33600
rect 13906 33464 13912 33516
rect 13964 33504 13970 33516
rect 14366 33504 14372 33516
rect 13964 33476 14372 33504
rect 13964 33464 13970 33476
rect 14366 33464 14372 33476
rect 14424 33504 14430 33516
rect 15194 33504 15200 33516
rect 14424 33476 15200 33504
rect 14424 33464 14430 33476
rect 15194 33464 15200 33476
rect 15252 33464 15258 33516
rect 15396 33504 15424 33612
rect 16758 33600 16764 33612
rect 16816 33600 16822 33652
rect 16945 33643 17003 33649
rect 16945 33609 16957 33643
rect 16991 33609 17003 33643
rect 16945 33603 17003 33609
rect 16574 33532 16580 33584
rect 16632 33572 16638 33584
rect 16960 33572 16988 33603
rect 18230 33600 18236 33652
rect 18288 33600 18294 33652
rect 18601 33643 18659 33649
rect 18601 33609 18613 33643
rect 18647 33640 18659 33643
rect 18647 33612 19564 33640
rect 18647 33609 18659 33612
rect 18601 33603 18659 33609
rect 16632 33544 16988 33572
rect 18248 33572 18276 33600
rect 18248 33544 18828 33572
rect 16632 33532 16638 33544
rect 15455 33507 15513 33513
rect 15455 33504 15467 33507
rect 15396 33476 15467 33504
rect 15455 33473 15467 33476
rect 15501 33473 15513 33507
rect 15455 33467 15513 33473
rect 17126 33464 17132 33516
rect 17184 33464 17190 33516
rect 17218 33464 17224 33516
rect 17276 33464 17282 33516
rect 17310 33464 17316 33516
rect 17368 33504 17374 33516
rect 18800 33513 18828 33544
rect 18966 33532 18972 33584
rect 19024 33532 19030 33584
rect 17477 33507 17535 33513
rect 17477 33504 17489 33507
rect 17368 33476 17489 33504
rect 17368 33464 17374 33476
rect 17477 33473 17489 33476
rect 17523 33473 17535 33507
rect 18693 33507 18751 33513
rect 18693 33504 18705 33507
rect 17477 33467 17535 33473
rect 18616 33476 18705 33504
rect 18616 33448 18644 33476
rect 18693 33473 18705 33476
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 18785 33507 18843 33513
rect 18785 33473 18797 33507
rect 18831 33473 18843 33507
rect 19061 33507 19119 33513
rect 19061 33504 19073 33507
rect 18785 33467 18843 33473
rect 18892 33476 19073 33504
rect 13035 33408 13768 33436
rect 13035 33405 13047 33408
rect 12989 33399 13047 33405
rect 18598 33396 18604 33448
rect 18656 33436 18662 33448
rect 18892 33436 18920 33476
rect 19061 33473 19073 33476
rect 19107 33473 19119 33507
rect 19061 33467 19119 33473
rect 19150 33464 19156 33516
rect 19208 33464 19214 33516
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33504 19303 33507
rect 19426 33504 19432 33516
rect 19291 33476 19432 33504
rect 19291 33473 19303 33476
rect 19245 33467 19303 33473
rect 19426 33464 19432 33476
rect 19484 33464 19490 33516
rect 19536 33513 19564 33612
rect 22646 33600 22652 33652
rect 22704 33600 22710 33652
rect 22830 33600 22836 33652
rect 22888 33640 22894 33652
rect 23201 33643 23259 33649
rect 23201 33640 23213 33643
rect 22888 33612 23213 33640
rect 22888 33600 22894 33612
rect 23201 33609 23213 33612
rect 23247 33609 23259 33643
rect 23201 33603 23259 33609
rect 23658 33600 23664 33652
rect 23716 33600 23722 33652
rect 19521 33507 19579 33513
rect 19521 33473 19533 33507
rect 19567 33473 19579 33507
rect 19521 33467 19579 33473
rect 20990 33464 20996 33516
rect 21048 33504 21054 33516
rect 21637 33507 21695 33513
rect 21637 33504 21649 33507
rect 21048 33476 21649 33504
rect 21048 33464 21054 33476
rect 21637 33473 21649 33476
rect 21683 33504 21695 33507
rect 22077 33507 22135 33513
rect 22077 33504 22089 33507
rect 21683 33476 22089 33504
rect 21683 33473 21695 33476
rect 21637 33467 21695 33473
rect 22077 33473 22089 33476
rect 22123 33473 22135 33507
rect 22664 33504 22692 33600
rect 23676 33572 23704 33600
rect 24121 33575 24179 33581
rect 24121 33572 24133 33575
rect 23676 33544 24133 33572
rect 24121 33541 24133 33544
rect 24167 33541 24179 33575
rect 24121 33535 24179 33541
rect 22664 33476 23060 33504
rect 22077 33467 22135 33473
rect 18656 33408 18920 33436
rect 18969 33439 19027 33445
rect 18656 33396 18662 33408
rect 18969 33405 18981 33439
rect 19015 33405 19027 33439
rect 19168 33436 19196 33464
rect 21542 33436 21548 33448
rect 19168 33408 21548 33436
rect 18969 33399 19027 33405
rect 11514 33328 11520 33380
rect 11572 33368 11578 33380
rect 12158 33368 12164 33380
rect 11572 33340 12164 33368
rect 11572 33328 11578 33340
rect 12158 33328 12164 33340
rect 12216 33328 12222 33380
rect 12437 33371 12495 33377
rect 12437 33337 12449 33371
rect 12483 33337 12495 33371
rect 18984 33368 19012 33399
rect 21542 33396 21548 33408
rect 21600 33436 21606 33448
rect 21821 33439 21879 33445
rect 21821 33436 21833 33439
rect 21600 33408 21833 33436
rect 21600 33396 21606 33408
rect 21821 33405 21833 33408
rect 21867 33405 21879 33439
rect 21821 33399 21879 33405
rect 19153 33371 19211 33377
rect 19153 33368 19165 33371
rect 12437 33331 12495 33337
rect 16132 33340 17264 33368
rect 18984 33340 19165 33368
rect 10318 33300 10324 33312
rect 9508 33272 10324 33300
rect 5905 33263 5963 33269
rect 10318 33260 10324 33272
rect 10376 33260 10382 33312
rect 10502 33260 10508 33312
rect 10560 33260 10566 33312
rect 12452 33300 12480 33331
rect 12894 33300 12900 33312
rect 12452 33272 12900 33300
rect 12894 33260 12900 33272
rect 12952 33260 12958 33312
rect 13633 33303 13691 33309
rect 13633 33269 13645 33303
rect 13679 33300 13691 33303
rect 16132 33300 16160 33340
rect 13679 33272 16160 33300
rect 13679 33269 13691 33272
rect 13633 33263 13691 33269
rect 16206 33260 16212 33312
rect 16264 33260 16270 33312
rect 17236 33300 17264 33340
rect 19153 33337 19165 33340
rect 19199 33337 19211 33371
rect 19153 33331 19211 33337
rect 19337 33371 19395 33377
rect 19337 33337 19349 33371
rect 19383 33368 19395 33371
rect 19426 33368 19432 33380
rect 19383 33340 19432 33368
rect 19383 33337 19395 33340
rect 19337 33331 19395 33337
rect 19426 33328 19432 33340
rect 19484 33328 19490 33380
rect 23032 33368 23060 33476
rect 23106 33464 23112 33516
rect 23164 33504 23170 33516
rect 23293 33507 23351 33513
rect 23293 33504 23305 33507
rect 23164 33476 23305 33504
rect 23164 33464 23170 33476
rect 23293 33473 23305 33476
rect 23339 33504 23351 33507
rect 23661 33507 23719 33513
rect 23661 33504 23673 33507
rect 23339 33476 23673 33504
rect 23339 33473 23351 33476
rect 23293 33467 23351 33473
rect 23661 33473 23673 33476
rect 23707 33473 23719 33507
rect 23661 33467 23719 33473
rect 23845 33507 23903 33513
rect 23845 33473 23857 33507
rect 23891 33473 23903 33507
rect 23845 33467 23903 33473
rect 23569 33439 23627 33445
rect 23569 33405 23581 33439
rect 23615 33436 23627 33439
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 23615 33408 23765 33436
rect 23615 33405 23627 33408
rect 23569 33399 23627 33405
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 23860 33368 23888 33467
rect 25406 33368 25412 33380
rect 23032 33340 23888 33368
rect 24320 33340 25412 33368
rect 20990 33300 20996 33312
rect 17236 33272 20996 33300
rect 20990 33260 20996 33272
rect 21048 33260 21054 33312
rect 21453 33303 21511 33309
rect 21453 33269 21465 33303
rect 21499 33300 21511 33303
rect 22186 33300 22192 33312
rect 21499 33272 22192 33300
rect 21499 33269 21511 33272
rect 21453 33263 21511 33269
rect 22186 33260 22192 33272
rect 22244 33260 22250 33312
rect 23382 33260 23388 33312
rect 23440 33260 23446 33312
rect 23477 33303 23535 33309
rect 23477 33269 23489 33303
rect 23523 33300 23535 33303
rect 24320 33300 24348 33340
rect 25406 33328 25412 33340
rect 25464 33328 25470 33380
rect 23523 33272 24348 33300
rect 23523 33269 23535 33272
rect 23477 33263 23535 33269
rect 24394 33260 24400 33312
rect 24452 33260 24458 33312
rect 1104 33210 24840 33232
rect 1104 33158 3917 33210
rect 3969 33158 3981 33210
rect 4033 33158 4045 33210
rect 4097 33158 4109 33210
rect 4161 33158 4173 33210
rect 4225 33158 9851 33210
rect 9903 33158 9915 33210
rect 9967 33158 9979 33210
rect 10031 33158 10043 33210
rect 10095 33158 10107 33210
rect 10159 33158 15785 33210
rect 15837 33158 15849 33210
rect 15901 33158 15913 33210
rect 15965 33158 15977 33210
rect 16029 33158 16041 33210
rect 16093 33158 21719 33210
rect 21771 33158 21783 33210
rect 21835 33158 21847 33210
rect 21899 33158 21911 33210
rect 21963 33158 21975 33210
rect 22027 33158 24840 33210
rect 1104 33136 24840 33158
rect 3329 33099 3387 33105
rect 2424 33068 3004 33096
rect 1394 32988 1400 33040
rect 1452 33028 1458 33040
rect 2424 33028 2452 33068
rect 1452 33000 2452 33028
rect 1452 32988 1458 33000
rect 2332 32969 2360 33000
rect 2317 32963 2375 32969
rect 2317 32929 2329 32963
rect 2363 32929 2375 32963
rect 2976 32960 3004 33068
rect 3329 33065 3341 33099
rect 3375 33096 3387 33099
rect 3418 33096 3424 33108
rect 3375 33068 3424 33096
rect 3375 33065 3387 33068
rect 3329 33059 3387 33065
rect 3418 33056 3424 33068
rect 3476 33056 3482 33108
rect 6362 33056 6368 33108
rect 6420 33096 6426 33108
rect 6420 33068 8064 33096
rect 6420 33056 6426 33068
rect 8036 33028 8064 33068
rect 8110 33056 8116 33108
rect 8168 33096 8174 33108
rect 8205 33099 8263 33105
rect 8205 33096 8217 33099
rect 8168 33068 8217 33096
rect 8168 33056 8174 33068
rect 8205 33065 8217 33068
rect 8251 33065 8263 33099
rect 11054 33096 11060 33108
rect 8205 33059 8263 33065
rect 10152 33068 11060 33096
rect 9398 33028 9404 33040
rect 8036 33000 9404 33028
rect 9398 32988 9404 33000
rect 9456 32988 9462 33040
rect 3326 32960 3332 32972
rect 2976 32932 3332 32960
rect 2317 32923 2375 32929
rect 3326 32920 3332 32932
rect 3384 32920 3390 32972
rect 4154 32960 4160 32972
rect 3620 32932 4160 32960
rect 1394 32852 1400 32904
rect 1452 32852 1458 32904
rect 2591 32895 2649 32901
rect 2591 32861 2603 32895
rect 2637 32892 2649 32895
rect 3620 32892 3648 32932
rect 4154 32920 4160 32932
rect 4212 32920 4218 32972
rect 5534 32920 5540 32972
rect 5592 32920 5598 32972
rect 6178 32920 6184 32972
rect 6236 32960 6242 32972
rect 10152 32969 10180 33068
rect 11054 33056 11060 33068
rect 11112 33056 11118 33108
rect 11793 33099 11851 33105
rect 11793 33065 11805 33099
rect 11839 33096 11851 33099
rect 11839 33068 12848 33096
rect 11839 33065 11851 33068
rect 11793 33059 11851 33065
rect 7193 32963 7251 32969
rect 7193 32960 7205 32963
rect 6236 32932 7205 32960
rect 6236 32920 6242 32932
rect 7193 32929 7205 32932
rect 7239 32929 7251 32963
rect 10137 32963 10195 32969
rect 10137 32960 10149 32963
rect 7193 32923 7251 32929
rect 9232 32932 10149 32960
rect 2637 32864 3648 32892
rect 3712 32864 5212 32892
rect 2637 32861 2649 32864
rect 2591 32855 2649 32861
rect 1673 32827 1731 32833
rect 1673 32793 1685 32827
rect 1719 32824 1731 32827
rect 3712 32824 3740 32864
rect 1719 32796 3740 32824
rect 3789 32827 3847 32833
rect 1719 32793 1731 32796
rect 1673 32787 1731 32793
rect 3789 32793 3801 32827
rect 3835 32793 3847 32827
rect 3789 32787 3847 32793
rect 1302 32716 1308 32768
rect 1360 32756 1366 32768
rect 3804 32756 3832 32787
rect 4522 32784 4528 32836
rect 4580 32784 4586 32836
rect 1360 32728 3832 32756
rect 1360 32716 1366 32728
rect 4890 32716 4896 32768
rect 4948 32756 4954 32768
rect 4985 32759 5043 32765
rect 4985 32756 4997 32759
rect 4948 32728 4997 32756
rect 4948 32716 4954 32728
rect 4985 32725 4997 32728
rect 5031 32725 5043 32759
rect 5184 32756 5212 32864
rect 5258 32852 5264 32904
rect 5316 32852 5322 32904
rect 5350 32852 5356 32904
rect 5408 32852 5414 32904
rect 5442 32852 5448 32904
rect 5500 32892 5506 32904
rect 5721 32895 5779 32901
rect 5721 32892 5733 32895
rect 5500 32864 5733 32892
rect 5500 32852 5506 32864
rect 5721 32861 5733 32864
rect 5767 32861 5779 32895
rect 5721 32855 5779 32861
rect 5810 32852 5816 32904
rect 5868 32892 5874 32904
rect 6196 32892 6224 32920
rect 9232 32904 9260 32932
rect 10137 32929 10149 32932
rect 10183 32929 10195 32963
rect 10137 32923 10195 32929
rect 10502 32920 10508 32972
rect 10560 32960 10566 32972
rect 10597 32963 10655 32969
rect 10597 32960 10609 32963
rect 10560 32932 10609 32960
rect 10560 32920 10566 32932
rect 10597 32929 10609 32932
rect 10643 32929 10655 32963
rect 10597 32923 10655 32929
rect 10686 32920 10692 32972
rect 10744 32960 10750 32972
rect 10873 32963 10931 32969
rect 10873 32960 10885 32963
rect 10744 32932 10885 32960
rect 10744 32920 10750 32932
rect 10873 32929 10885 32932
rect 10919 32929 10931 32963
rect 10873 32923 10931 32929
rect 11011 32963 11069 32969
rect 11011 32929 11023 32963
rect 11057 32960 11069 32963
rect 11330 32960 11336 32972
rect 11057 32932 11336 32960
rect 11057 32929 11069 32932
rect 11011 32923 11069 32929
rect 11330 32920 11336 32932
rect 11388 32960 11394 32972
rect 11514 32960 11520 32972
rect 11388 32932 11520 32960
rect 11388 32920 11394 32932
rect 11514 32920 11520 32932
rect 11572 32920 11578 32972
rect 11882 32920 11888 32972
rect 11940 32920 11946 32972
rect 12820 32960 12848 33068
rect 12894 33056 12900 33108
rect 12952 33056 12958 33108
rect 15102 33096 15108 33108
rect 14752 33068 15108 33096
rect 14752 33037 14780 33068
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 15378 33056 15384 33108
rect 15436 33096 15442 33108
rect 15933 33099 15991 33105
rect 15436 33068 15884 33096
rect 15436 33056 15442 33068
rect 14737 33031 14795 33037
rect 14737 32997 14749 33031
rect 14783 32997 14795 33031
rect 15856 33028 15884 33068
rect 15933 33065 15945 33099
rect 15979 33096 15991 33099
rect 16114 33096 16120 33108
rect 15979 33068 16120 33096
rect 15979 33065 15991 33068
rect 15933 33059 15991 33065
rect 16114 33056 16120 33068
rect 16172 33056 16178 33108
rect 18598 33056 18604 33108
rect 18656 33056 18662 33108
rect 22281 33099 22339 33105
rect 22281 33065 22293 33099
rect 22327 33096 22339 33099
rect 23382 33096 23388 33108
rect 22327 33068 23388 33096
rect 22327 33065 22339 33068
rect 22281 33059 22339 33065
rect 23382 33056 23388 33068
rect 23440 33056 23446 33108
rect 21913 33031 21971 33037
rect 15856 33000 17448 33028
rect 14737 32991 14795 32997
rect 17310 32960 17316 32972
rect 12820 32932 17316 32960
rect 17310 32920 17316 32932
rect 17368 32920 17374 32972
rect 17420 32904 17448 33000
rect 21913 32997 21925 33031
rect 21959 33028 21971 33031
rect 23661 33031 23719 33037
rect 21959 33000 23060 33028
rect 21959 32997 21971 33000
rect 21913 32991 21971 32997
rect 17586 32920 17592 32972
rect 17644 32920 17650 32972
rect 7466 32892 7472 32904
rect 5868 32864 6224 32892
rect 7427 32864 7472 32892
rect 5868 32852 5874 32864
rect 7466 32852 7472 32864
rect 7524 32892 7530 32904
rect 8110 32892 8116 32904
rect 7524 32864 8116 32892
rect 7524 32852 7530 32864
rect 8110 32852 8116 32864
rect 8168 32852 8174 32904
rect 9214 32852 9220 32904
rect 9272 32852 9278 32904
rect 9766 32852 9772 32904
rect 9824 32892 9830 32904
rect 9953 32895 10011 32901
rect 9953 32892 9965 32895
rect 9824 32864 9965 32892
rect 9824 32852 9830 32864
rect 9953 32861 9965 32864
rect 9999 32861 10011 32895
rect 9953 32855 10011 32861
rect 11146 32852 11152 32904
rect 11204 32852 11210 32904
rect 12159 32895 12217 32901
rect 12159 32861 12171 32895
rect 12205 32892 12217 32895
rect 12205 32864 12572 32892
rect 12205 32861 12217 32864
rect 12159 32855 12217 32861
rect 10134 32824 10140 32836
rect 5644 32796 10140 32824
rect 5644 32756 5672 32796
rect 10134 32784 10140 32796
rect 10192 32784 10198 32836
rect 12544 32824 12572 32864
rect 12618 32852 12624 32904
rect 12676 32892 12682 32904
rect 14093 32895 14151 32901
rect 14093 32892 14105 32895
rect 12676 32864 14105 32892
rect 12676 32852 12682 32864
rect 14093 32861 14105 32864
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 12710 32824 12716 32836
rect 11624 32796 12434 32824
rect 12544 32796 12716 32824
rect 5184 32728 5672 32756
rect 6089 32759 6147 32765
rect 4985 32719 5043 32725
rect 6089 32725 6101 32759
rect 6135 32756 6147 32759
rect 6178 32756 6184 32768
rect 6135 32728 6184 32756
rect 6135 32725 6147 32728
rect 6089 32719 6147 32725
rect 6178 32716 6184 32728
rect 6236 32716 6242 32768
rect 6273 32759 6331 32765
rect 6273 32725 6285 32759
rect 6319 32756 6331 32759
rect 11624 32756 11652 32796
rect 6319 32728 11652 32756
rect 12406 32756 12434 32796
rect 12710 32784 12716 32796
rect 12768 32824 12774 32836
rect 13538 32824 13544 32836
rect 12768 32796 13544 32824
rect 12768 32784 12774 32796
rect 13538 32784 13544 32796
rect 13596 32784 13602 32836
rect 13998 32756 14004 32768
rect 12406 32728 14004 32756
rect 6319 32725 6331 32728
rect 6273 32719 6331 32725
rect 13998 32716 14004 32728
rect 14056 32716 14062 32768
rect 14292 32756 14320 32855
rect 15010 32852 15016 32904
rect 15068 32852 15074 32904
rect 15102 32852 15108 32904
rect 15160 32901 15166 32904
rect 15160 32895 15188 32901
rect 15176 32861 15188 32895
rect 15160 32855 15188 32861
rect 15160 32852 15166 32855
rect 15286 32852 15292 32904
rect 15344 32852 15350 32904
rect 17402 32852 17408 32904
rect 17460 32892 17466 32904
rect 17862 32901 17868 32904
rect 17831 32895 17868 32901
rect 17831 32892 17843 32895
rect 17460 32864 17843 32892
rect 17460 32852 17466 32864
rect 17831 32861 17843 32864
rect 17831 32855 17868 32861
rect 17862 32852 17868 32855
rect 17920 32852 17926 32904
rect 22097 32895 22155 32901
rect 22097 32861 22109 32895
rect 22143 32861 22155 32895
rect 22097 32855 22155 32861
rect 16850 32784 16856 32836
rect 16908 32824 16914 32836
rect 19702 32824 19708 32836
rect 16908 32796 19708 32824
rect 16908 32784 16914 32796
rect 19702 32784 19708 32796
rect 19760 32784 19766 32836
rect 15286 32756 15292 32768
rect 14292 32728 15292 32756
rect 15286 32716 15292 32728
rect 15344 32716 15350 32768
rect 15378 32716 15384 32768
rect 15436 32756 15442 32768
rect 22112 32756 22140 32855
rect 22186 32852 22192 32904
rect 22244 32852 22250 32904
rect 23032 32901 23060 33000
rect 23661 32997 23673 33031
rect 23707 32997 23719 33031
rect 23661 32991 23719 32997
rect 23017 32895 23075 32901
rect 23017 32861 23029 32895
rect 23063 32861 23075 32895
rect 23017 32855 23075 32861
rect 23569 32895 23627 32901
rect 23569 32861 23581 32895
rect 23615 32892 23627 32895
rect 23676 32892 23704 32991
rect 23615 32864 23704 32892
rect 23845 32895 23903 32901
rect 23615 32861 23627 32864
rect 23569 32855 23627 32861
rect 23845 32861 23857 32895
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 23198 32784 23204 32836
rect 23256 32784 23262 32836
rect 23290 32784 23296 32836
rect 23348 32784 23354 32836
rect 23860 32824 23888 32855
rect 23934 32852 23940 32904
rect 23992 32852 23998 32904
rect 25130 32824 25136 32836
rect 23860 32796 25136 32824
rect 25130 32784 25136 32796
rect 25188 32784 25194 32836
rect 22646 32756 22652 32768
rect 15436 32728 22652 32756
rect 15436 32716 15442 32728
rect 22646 32716 22652 32728
rect 22704 32716 22710 32768
rect 22833 32759 22891 32765
rect 22833 32725 22845 32759
rect 22879 32756 22891 32759
rect 23216 32756 23244 32784
rect 22879 32728 23244 32756
rect 23308 32756 23336 32784
rect 23385 32759 23443 32765
rect 23385 32756 23397 32759
rect 23308 32728 23397 32756
rect 22879 32725 22891 32728
rect 22833 32719 22891 32725
rect 23385 32725 23397 32728
rect 23431 32725 23443 32759
rect 23385 32719 23443 32725
rect 24121 32759 24179 32765
rect 24121 32725 24133 32759
rect 24167 32756 24179 32759
rect 25222 32756 25228 32768
rect 24167 32728 25228 32756
rect 24167 32725 24179 32728
rect 24121 32719 24179 32725
rect 25222 32716 25228 32728
rect 25280 32716 25286 32768
rect 1104 32666 25000 32688
rect 1104 32614 6884 32666
rect 6936 32614 6948 32666
rect 7000 32614 7012 32666
rect 7064 32614 7076 32666
rect 7128 32614 7140 32666
rect 7192 32614 12818 32666
rect 12870 32614 12882 32666
rect 12934 32614 12946 32666
rect 12998 32614 13010 32666
rect 13062 32614 13074 32666
rect 13126 32614 18752 32666
rect 18804 32614 18816 32666
rect 18868 32614 18880 32666
rect 18932 32614 18944 32666
rect 18996 32614 19008 32666
rect 19060 32614 24686 32666
rect 24738 32614 24750 32666
rect 24802 32614 24814 32666
rect 24866 32614 24878 32666
rect 24930 32614 24942 32666
rect 24994 32614 25000 32666
rect 1104 32592 25000 32614
rect 1210 32512 1216 32564
rect 1268 32552 1274 32564
rect 1268 32524 3924 32552
rect 1268 32512 1274 32524
rect 3237 32487 3295 32493
rect 3237 32453 3249 32487
rect 3283 32484 3295 32487
rect 3694 32484 3700 32496
rect 3283 32456 3700 32484
rect 3283 32453 3295 32456
rect 3237 32447 3295 32453
rect 3694 32444 3700 32456
rect 3752 32444 3758 32496
rect 2314 32376 2320 32428
rect 2372 32376 2378 32428
rect 2434 32419 2492 32425
rect 2434 32416 2446 32419
rect 2424 32385 2446 32416
rect 2480 32385 2492 32419
rect 2424 32379 2492 32385
rect 1397 32351 1455 32357
rect 1397 32317 1409 32351
rect 1443 32348 1455 32351
rect 1486 32348 1492 32360
rect 1443 32320 1492 32348
rect 1443 32317 1455 32320
rect 1397 32311 1455 32317
rect 1486 32308 1492 32320
rect 1544 32308 1550 32360
rect 1578 32308 1584 32360
rect 1636 32308 1642 32360
rect 1762 32308 1768 32360
rect 1820 32348 1826 32360
rect 2041 32351 2099 32357
rect 2041 32348 2053 32351
rect 1820 32320 2053 32348
rect 1820 32308 1826 32320
rect 2041 32317 2053 32320
rect 2087 32317 2099 32351
rect 2424 32348 2452 32379
rect 2588 32376 2594 32428
rect 2646 32376 2652 32428
rect 3326 32376 3332 32428
rect 3384 32376 3390 32428
rect 3896 32425 3924 32524
rect 4522 32512 4528 32564
rect 4580 32512 4586 32564
rect 5166 32512 5172 32564
rect 5224 32552 5230 32564
rect 5350 32552 5356 32564
rect 5224 32524 5356 32552
rect 5224 32512 5230 32524
rect 5350 32512 5356 32524
rect 5408 32552 5414 32564
rect 6178 32552 6184 32564
rect 5408 32524 6184 32552
rect 5408 32512 5414 32524
rect 6178 32512 6184 32524
rect 6236 32512 6242 32564
rect 10134 32512 10140 32564
rect 10192 32552 10198 32564
rect 10594 32552 10600 32564
rect 10192 32524 10600 32552
rect 10192 32512 10198 32524
rect 10594 32512 10600 32524
rect 10652 32512 10658 32564
rect 11057 32555 11115 32561
rect 11057 32521 11069 32555
rect 11103 32552 11115 32555
rect 11146 32552 11152 32564
rect 11103 32524 11152 32552
rect 11103 32521 11115 32524
rect 11057 32515 11115 32521
rect 11146 32512 11152 32524
rect 11204 32512 11210 32564
rect 15010 32552 15016 32564
rect 14384 32524 15016 32552
rect 4540 32484 4568 32512
rect 6730 32484 6736 32496
rect 4540 32456 6736 32484
rect 6730 32444 6736 32456
rect 6788 32444 6794 32496
rect 8570 32484 8576 32496
rect 8036 32456 8576 32484
rect 3881 32419 3939 32425
rect 3881 32385 3893 32419
rect 3927 32385 3939 32419
rect 4154 32416 4160 32428
rect 3881 32379 3939 32385
rect 3988 32388 4160 32416
rect 2041 32311 2099 32317
rect 2148 32320 2452 32348
rect 3605 32351 3663 32357
rect 1854 32240 1860 32292
rect 1912 32280 1918 32292
rect 2148 32280 2176 32320
rect 3605 32317 3617 32351
rect 3651 32348 3663 32351
rect 3988 32348 4016 32388
rect 4154 32376 4160 32388
rect 4212 32376 4218 32428
rect 4614 32376 4620 32428
rect 4672 32376 4678 32428
rect 4890 32376 4896 32428
rect 4948 32416 4954 32428
rect 6086 32416 6092 32428
rect 4948 32388 6092 32416
rect 4948 32376 4954 32388
rect 6086 32376 6092 32388
rect 6144 32376 6150 32428
rect 6178 32376 6184 32428
rect 6236 32416 6242 32428
rect 6454 32416 6460 32428
rect 6236 32388 6460 32416
rect 6236 32376 6242 32388
rect 6454 32376 6460 32388
rect 6512 32376 6518 32428
rect 8036 32425 8064 32456
rect 8570 32444 8576 32456
rect 8628 32484 8634 32496
rect 14384 32493 14412 32524
rect 15010 32512 15016 32524
rect 15068 32512 15074 32564
rect 15197 32555 15255 32561
rect 15197 32521 15209 32555
rect 15243 32552 15255 32555
rect 15286 32552 15292 32564
rect 15243 32524 15292 32552
rect 15243 32521 15255 32524
rect 15197 32515 15255 32521
rect 15286 32512 15292 32524
rect 15344 32512 15350 32564
rect 15381 32555 15439 32561
rect 15381 32521 15393 32555
rect 15427 32552 15439 32555
rect 21266 32552 21272 32564
rect 15427 32524 21272 32552
rect 15427 32521 15439 32524
rect 15381 32515 15439 32521
rect 21266 32512 21272 32524
rect 21324 32512 21330 32564
rect 22649 32555 22707 32561
rect 22649 32521 22661 32555
rect 22695 32552 22707 32555
rect 23661 32555 23719 32561
rect 22695 32524 23612 32552
rect 22695 32521 22707 32524
rect 22649 32515 22707 32521
rect 14093 32487 14151 32493
rect 8628 32456 9168 32484
rect 8628 32444 8634 32456
rect 9140 32428 9168 32456
rect 10060 32456 10456 32484
rect 8021 32419 8079 32425
rect 8021 32385 8033 32419
rect 8067 32385 8079 32419
rect 8021 32379 8079 32385
rect 8202 32376 8208 32428
rect 8260 32416 8266 32428
rect 8295 32419 8353 32425
rect 8295 32416 8307 32419
rect 8260 32388 8307 32416
rect 8260 32376 8266 32388
rect 8295 32385 8307 32388
rect 8341 32416 8353 32419
rect 8386 32416 8392 32428
rect 8341 32388 8392 32416
rect 8341 32385 8353 32388
rect 8295 32379 8353 32385
rect 8386 32376 8392 32388
rect 8444 32376 8450 32428
rect 9122 32376 9128 32428
rect 9180 32376 9186 32428
rect 10060 32425 10088 32456
rect 10428 32428 10456 32456
rect 14093 32453 14105 32487
rect 14139 32453 14151 32487
rect 14093 32447 14151 32453
rect 14369 32487 14427 32493
rect 14369 32453 14381 32487
rect 14415 32453 14427 32487
rect 14369 32447 14427 32453
rect 10045 32419 10103 32425
rect 10045 32385 10057 32419
rect 10091 32385 10103 32419
rect 10318 32416 10324 32428
rect 10279 32388 10324 32416
rect 10045 32379 10103 32385
rect 10318 32376 10324 32388
rect 10376 32376 10382 32428
rect 10410 32376 10416 32428
rect 10468 32416 10474 32428
rect 11974 32416 11980 32428
rect 10468 32388 11980 32416
rect 10468 32376 10474 32388
rect 11974 32376 11980 32388
rect 12032 32376 12038 32428
rect 14108 32416 14136 32447
rect 14458 32444 14464 32496
rect 14516 32444 14522 32496
rect 15102 32484 15108 32496
rect 14660 32456 15108 32484
rect 14660 32416 14688 32456
rect 15102 32444 15108 32456
rect 15160 32484 15166 32496
rect 15160 32456 16712 32484
rect 15160 32444 15166 32456
rect 14108 32388 14688 32416
rect 14826 32376 14832 32428
rect 14884 32376 14890 32428
rect 3651 32320 4016 32348
rect 3651 32317 3663 32320
rect 3605 32311 3663 32317
rect 4062 32308 4068 32360
rect 4120 32308 4126 32360
rect 4172 32348 4200 32376
rect 15108 32360 15160 32366
rect 16684 32360 16712 32456
rect 19334 32444 19340 32496
rect 19392 32484 19398 32496
rect 19392 32456 19472 32484
rect 19392 32444 19398 32456
rect 17678 32376 17684 32428
rect 17736 32416 17742 32428
rect 19150 32416 19156 32428
rect 17736 32388 19156 32416
rect 17736 32376 17742 32388
rect 19150 32376 19156 32388
rect 19208 32376 19214 32428
rect 19444 32425 19472 32456
rect 19420 32419 19478 32425
rect 19420 32385 19432 32419
rect 19466 32385 19478 32419
rect 19420 32379 19478 32385
rect 19702 32376 19708 32428
rect 19760 32416 19766 32428
rect 23584 32425 23612 32524
rect 23661 32521 23673 32555
rect 23707 32552 23719 32555
rect 23934 32552 23940 32564
rect 23707 32524 23940 32552
rect 23707 32521 23719 32524
rect 23661 32515 23719 32521
rect 23934 32512 23940 32524
rect 23992 32512 23998 32564
rect 22005 32419 22063 32425
rect 22005 32416 22017 32419
rect 19760 32388 22017 32416
rect 19760 32376 19766 32388
rect 22005 32385 22017 32388
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22557 32419 22615 32425
rect 22557 32385 22569 32419
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32385 22891 32419
rect 23293 32419 23351 32425
rect 23293 32416 23305 32419
rect 22833 32379 22891 32385
rect 22940 32388 23305 32416
rect 4982 32348 4988 32360
rect 4172 32320 4988 32348
rect 4982 32308 4988 32320
rect 5040 32348 5046 32360
rect 5166 32348 5172 32360
rect 5040 32320 5172 32348
rect 5040 32308 5046 32320
rect 5166 32308 5172 32320
rect 5224 32308 5230 32360
rect 15194 32308 15200 32360
rect 15252 32348 15258 32360
rect 15252 32320 16436 32348
rect 15252 32308 15258 32320
rect 15108 32302 15160 32308
rect 16408 32292 16436 32320
rect 16666 32308 16672 32360
rect 16724 32308 16730 32360
rect 22572 32348 22600 32379
rect 22066 32320 22600 32348
rect 1912 32252 2176 32280
rect 1912 32240 1918 32252
rect 2148 32212 2176 32252
rect 16390 32240 16396 32292
rect 16448 32280 16454 32292
rect 21821 32283 21879 32289
rect 16448 32252 18644 32280
rect 16448 32240 16454 32252
rect 18616 32224 18644 32252
rect 20088 32252 20668 32280
rect 3050 32212 3056 32224
rect 2148 32184 3056 32212
rect 3050 32172 3056 32184
rect 3108 32172 3114 32224
rect 4062 32172 4068 32224
rect 4120 32212 4126 32224
rect 5718 32212 5724 32224
rect 4120 32184 5724 32212
rect 4120 32172 4126 32184
rect 5718 32172 5724 32184
rect 5776 32172 5782 32224
rect 9030 32172 9036 32224
rect 9088 32172 9094 32224
rect 16574 32172 16580 32224
rect 16632 32212 16638 32224
rect 17034 32212 17040 32224
rect 16632 32184 17040 32212
rect 16632 32172 16638 32184
rect 17034 32172 17040 32184
rect 17092 32172 17098 32224
rect 18598 32172 18604 32224
rect 18656 32212 18662 32224
rect 20088 32212 20116 32252
rect 18656 32184 20116 32212
rect 18656 32172 18662 32184
rect 20530 32172 20536 32224
rect 20588 32172 20594 32224
rect 20640 32212 20668 32252
rect 21821 32249 21833 32283
rect 21867 32280 21879 32283
rect 22066 32280 22094 32320
rect 22848 32280 22876 32379
rect 21867 32252 22094 32280
rect 22296 32252 22876 32280
rect 21867 32249 21879 32252
rect 21821 32243 21879 32249
rect 22296 32212 22324 32252
rect 20640 32184 22324 32212
rect 22373 32215 22431 32221
rect 22373 32181 22385 32215
rect 22419 32212 22431 32215
rect 22940 32212 22968 32388
rect 23293 32385 23305 32388
rect 23339 32385 23351 32419
rect 23293 32379 23351 32385
rect 23569 32419 23627 32425
rect 23569 32385 23581 32419
rect 23615 32385 23627 32419
rect 23569 32379 23627 32385
rect 23845 32419 23903 32425
rect 23845 32385 23857 32419
rect 23891 32385 23903 32419
rect 23845 32379 23903 32385
rect 23860 32348 23888 32379
rect 24118 32376 24124 32428
rect 24176 32376 24182 32428
rect 24213 32419 24271 32425
rect 24213 32385 24225 32419
rect 24259 32385 24271 32419
rect 24213 32379 24271 32385
rect 23400 32320 23888 32348
rect 23400 32289 23428 32320
rect 23385 32283 23443 32289
rect 23385 32249 23397 32283
rect 23431 32249 23443 32283
rect 24228 32280 24256 32379
rect 23385 32243 23443 32249
rect 23860 32252 24256 32280
rect 22419 32184 22968 32212
rect 23109 32215 23167 32221
rect 22419 32181 22431 32184
rect 22373 32175 22431 32181
rect 23109 32181 23121 32215
rect 23155 32212 23167 32215
rect 23860 32212 23888 32252
rect 23155 32184 23888 32212
rect 23937 32215 23995 32221
rect 23155 32181 23167 32184
rect 23109 32175 23167 32181
rect 23937 32181 23949 32215
rect 23983 32212 23995 32215
rect 24026 32212 24032 32224
rect 23983 32184 24032 32212
rect 23983 32181 23995 32184
rect 23937 32175 23995 32181
rect 24026 32172 24032 32184
rect 24084 32172 24090 32224
rect 24394 32172 24400 32224
rect 24452 32172 24458 32224
rect 1104 32122 24840 32144
rect 1104 32070 3917 32122
rect 3969 32070 3981 32122
rect 4033 32070 4045 32122
rect 4097 32070 4109 32122
rect 4161 32070 4173 32122
rect 4225 32070 9851 32122
rect 9903 32070 9915 32122
rect 9967 32070 9979 32122
rect 10031 32070 10043 32122
rect 10095 32070 10107 32122
rect 10159 32070 15785 32122
rect 15837 32070 15849 32122
rect 15901 32070 15913 32122
rect 15965 32070 15977 32122
rect 16029 32070 16041 32122
rect 16093 32070 21719 32122
rect 21771 32070 21783 32122
rect 21835 32070 21847 32122
rect 21899 32070 21911 32122
rect 21963 32070 21975 32122
rect 22027 32070 24840 32122
rect 1104 32048 24840 32070
rect 1486 31968 1492 32020
rect 1544 32008 1550 32020
rect 2409 32011 2467 32017
rect 1544 31980 2084 32008
rect 1544 31968 1550 31980
rect 2056 31872 2084 31980
rect 2409 31977 2421 32011
rect 2455 32008 2467 32011
rect 2590 32008 2596 32020
rect 2455 31980 2596 32008
rect 2455 31977 2467 31980
rect 2409 31971 2467 31977
rect 2590 31968 2596 31980
rect 2648 31968 2654 32020
rect 3234 31968 3240 32020
rect 3292 32008 3298 32020
rect 3510 32008 3516 32020
rect 3292 31980 3516 32008
rect 3292 31968 3298 31980
rect 3510 31968 3516 31980
rect 3568 31968 3574 32020
rect 4709 32011 4767 32017
rect 4709 31977 4721 32011
rect 4755 32008 4767 32011
rect 5074 32008 5080 32020
rect 4755 31980 5080 32008
rect 4755 31977 4767 31980
rect 4709 31971 4767 31977
rect 5074 31968 5080 31980
rect 5132 31968 5138 32020
rect 10502 32008 10508 32020
rect 5920 31980 10508 32008
rect 5920 31940 5948 31980
rect 10502 31968 10508 31980
rect 10560 31968 10566 32020
rect 11072 31980 13308 32008
rect 3068 31912 5948 31940
rect 3068 31881 3096 31912
rect 6822 31900 6828 31952
rect 6880 31900 6886 31952
rect 9674 31900 9680 31952
rect 9732 31940 9738 31952
rect 10318 31940 10324 31952
rect 9732 31912 10324 31940
rect 9732 31900 9738 31912
rect 10318 31900 10324 31912
rect 10376 31900 10382 31952
rect 3053 31875 3111 31881
rect 2056 31844 3004 31872
rect 750 31764 756 31816
rect 808 31804 814 31816
rect 1302 31804 1308 31816
rect 808 31776 1308 31804
rect 808 31764 814 31776
rect 1302 31764 1308 31776
rect 1360 31804 1366 31816
rect 1397 31807 1455 31813
rect 1397 31804 1409 31807
rect 1360 31776 1409 31804
rect 1360 31764 1366 31776
rect 1397 31773 1409 31776
rect 1443 31773 1455 31807
rect 2130 31804 2136 31816
rect 1688 31783 2136 31804
rect 1397 31767 1455 31773
rect 1655 31777 2136 31783
rect 1655 31743 1667 31777
rect 1701 31776 2136 31777
rect 1701 31746 1716 31776
rect 2130 31764 2136 31776
rect 2188 31764 2194 31816
rect 2774 31764 2780 31816
rect 2832 31764 2838 31816
rect 2976 31804 3004 31844
rect 3053 31841 3065 31875
rect 3099 31841 3111 31875
rect 3053 31835 3111 31841
rect 3510 31832 3516 31884
rect 3568 31872 3574 31884
rect 3973 31875 4031 31881
rect 3973 31872 3985 31875
rect 3568 31844 3985 31872
rect 3568 31832 3574 31844
rect 3973 31841 3985 31844
rect 4019 31841 4031 31875
rect 3973 31835 4031 31841
rect 5810 31832 5816 31884
rect 5868 31832 5874 31884
rect 8294 31832 8300 31884
rect 8352 31872 8358 31884
rect 8478 31872 8484 31884
rect 8352 31844 8484 31872
rect 8352 31832 8358 31844
rect 8478 31832 8484 31844
rect 8536 31832 8542 31884
rect 11072 31881 11100 31980
rect 13280 31952 13308 31980
rect 13906 31968 13912 32020
rect 13964 31968 13970 32020
rect 13998 31968 14004 32020
rect 14056 32008 14062 32020
rect 14056 31980 14780 32008
rect 14056 31968 14062 31980
rect 13262 31900 13268 31952
rect 13320 31900 13326 31952
rect 13924 31940 13952 31968
rect 14752 31940 14780 31980
rect 15102 31968 15108 32020
rect 15160 31968 15166 32020
rect 15286 31968 15292 32020
rect 15344 32008 15350 32020
rect 15746 32008 15752 32020
rect 15344 31980 15752 32008
rect 15344 31968 15350 31980
rect 15746 31968 15752 31980
rect 15804 31968 15810 32020
rect 19794 32008 19800 32020
rect 15856 31980 17172 32008
rect 15856 31940 15884 31980
rect 13924 31912 14136 31940
rect 14752 31912 15884 31940
rect 14108 31881 14136 31912
rect 16206 31900 16212 31952
rect 16264 31900 16270 31952
rect 17144 31940 17172 31980
rect 17512 31980 19800 32008
rect 17512 31940 17540 31980
rect 19794 31968 19800 31980
rect 19852 31968 19858 32020
rect 20530 31968 20536 32020
rect 20588 31968 20594 32020
rect 21637 32011 21695 32017
rect 21637 31977 21649 32011
rect 21683 32008 21695 32011
rect 23477 32011 23535 32017
rect 21683 31980 22094 32008
rect 21683 31977 21695 31980
rect 21637 31971 21695 31977
rect 17144 31912 17540 31940
rect 19334 31900 19340 31952
rect 19392 31940 19398 31952
rect 19521 31943 19579 31949
rect 19392 31912 19472 31940
rect 19392 31900 19398 31912
rect 11057 31875 11115 31881
rect 11057 31841 11069 31875
rect 11103 31841 11115 31875
rect 14093 31875 14151 31881
rect 11057 31835 11115 31841
rect 12452 31844 13952 31872
rect 3234 31804 3240 31816
rect 2976 31776 3240 31804
rect 3234 31764 3240 31776
rect 3292 31804 3298 31816
rect 3292 31776 3464 31804
rect 3292 31764 3298 31776
rect 1701 31743 1713 31746
rect 1655 31737 1713 31743
rect 3436 31736 3464 31776
rect 3786 31764 3792 31816
rect 3844 31764 3850 31816
rect 4890 31764 4896 31816
rect 4948 31764 4954 31816
rect 5534 31764 5540 31816
rect 5592 31804 5598 31816
rect 5592 31777 6130 31804
rect 5592 31776 6083 31777
rect 5592 31764 5598 31776
rect 5718 31736 5724 31748
rect 3436 31708 5724 31736
rect 5718 31696 5724 31708
rect 5776 31696 5782 31748
rect 6071 31743 6083 31776
rect 6117 31746 6130 31777
rect 6454 31764 6460 31816
rect 6512 31804 6518 31816
rect 11331 31807 11389 31813
rect 11331 31804 11343 31807
rect 6512 31776 11343 31804
rect 6512 31764 6518 31776
rect 11331 31773 11343 31776
rect 11377 31804 11389 31807
rect 12452 31804 12480 31844
rect 11377 31776 12480 31804
rect 11377 31773 11389 31776
rect 11331 31767 11389 31773
rect 12526 31764 12532 31816
rect 12584 31804 12590 31816
rect 13081 31807 13139 31813
rect 13081 31804 13093 31807
rect 12584 31776 13093 31804
rect 12584 31764 12590 31776
rect 13081 31773 13093 31776
rect 13127 31773 13139 31807
rect 13081 31767 13139 31773
rect 13173 31807 13231 31813
rect 13173 31773 13185 31807
rect 13219 31804 13231 31807
rect 13814 31804 13820 31816
rect 13219 31776 13820 31804
rect 13219 31773 13231 31776
rect 13173 31767 13231 31773
rect 13814 31764 13820 31776
rect 13872 31764 13878 31816
rect 13924 31804 13952 31844
rect 14093 31841 14105 31875
rect 14139 31841 14151 31875
rect 16602 31875 16660 31881
rect 16602 31872 16614 31875
rect 14093 31835 14151 31841
rect 15304 31844 16614 31872
rect 13924 31776 14228 31804
rect 6117 31743 6129 31746
rect 6071 31737 6129 31743
rect 6638 31696 6644 31748
rect 6696 31736 6702 31748
rect 14200 31736 14228 31776
rect 14274 31764 14280 31816
rect 14332 31804 14338 31816
rect 14367 31807 14425 31813
rect 14367 31804 14379 31807
rect 14332 31776 14379 31804
rect 14332 31764 14338 31776
rect 14367 31773 14379 31776
rect 14413 31773 14425 31807
rect 15194 31804 15200 31816
rect 14367 31767 14425 31773
rect 14458 31776 15200 31804
rect 14458 31736 14486 31776
rect 15194 31764 15200 31776
rect 15252 31764 15258 31816
rect 6696 31708 14136 31736
rect 14200 31708 14486 31736
rect 6696 31696 6702 31708
rect 1762 31628 1768 31680
rect 1820 31668 1826 31680
rect 7650 31668 7656 31680
rect 1820 31640 7656 31668
rect 1820 31628 1826 31640
rect 7650 31628 7656 31640
rect 7708 31628 7714 31680
rect 8478 31628 8484 31680
rect 8536 31668 8542 31680
rect 9214 31668 9220 31680
rect 8536 31640 9220 31668
rect 8536 31628 8542 31640
rect 9214 31628 9220 31640
rect 9272 31628 9278 31680
rect 12066 31628 12072 31680
rect 12124 31628 12130 31680
rect 14108 31668 14136 31708
rect 14826 31696 14832 31748
rect 14884 31736 14890 31748
rect 15304 31736 15332 31844
rect 16602 31841 16614 31844
rect 16648 31841 16660 31875
rect 16602 31835 16660 31841
rect 16761 31875 16819 31881
rect 16761 31841 16773 31875
rect 16807 31872 16819 31875
rect 16942 31872 16948 31884
rect 16807 31844 16948 31872
rect 16807 31841 16819 31844
rect 16761 31835 16819 31841
rect 16942 31832 16948 31844
rect 17000 31832 17006 31884
rect 17126 31832 17132 31884
rect 17184 31872 17190 31884
rect 17405 31875 17463 31881
rect 17405 31872 17417 31875
rect 17184 31844 17417 31872
rect 17184 31832 17190 31844
rect 17405 31841 17417 31844
rect 17451 31841 17463 31875
rect 17405 31835 17463 31841
rect 15470 31764 15476 31816
rect 15528 31804 15534 31816
rect 15565 31807 15623 31813
rect 15565 31804 15577 31807
rect 15528 31776 15577 31804
rect 15528 31764 15534 31776
rect 15565 31773 15577 31776
rect 15611 31773 15623 31807
rect 15565 31767 15623 31773
rect 15746 31764 15752 31816
rect 15804 31764 15810 31816
rect 16482 31764 16488 31816
rect 16540 31764 16546 31816
rect 19444 31804 19472 31912
rect 19521 31909 19533 31943
rect 19567 31909 19579 31943
rect 19521 31903 19579 31909
rect 19536 31872 19564 31903
rect 19536 31844 20116 31872
rect 20088 31813 20116 31844
rect 19705 31807 19763 31813
rect 19705 31804 19717 31807
rect 19444 31776 19717 31804
rect 19705 31773 19717 31776
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 20073 31807 20131 31813
rect 20073 31773 20085 31807
rect 20119 31773 20131 31807
rect 20073 31767 20131 31773
rect 20165 31807 20223 31813
rect 20165 31773 20177 31807
rect 20211 31804 20223 31807
rect 20548 31804 20576 31968
rect 20625 31943 20683 31949
rect 20625 31909 20637 31943
rect 20671 31940 20683 31943
rect 20714 31940 20720 31952
rect 20671 31912 20720 31940
rect 20671 31909 20683 31912
rect 20625 31903 20683 31909
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 20901 31943 20959 31949
rect 20901 31909 20913 31943
rect 20947 31909 20959 31943
rect 20901 31903 20959 31909
rect 21177 31943 21235 31949
rect 21177 31909 21189 31943
rect 21223 31940 21235 31943
rect 21223 31912 21864 31940
rect 21223 31909 21235 31912
rect 21177 31903 21235 31909
rect 20916 31872 20944 31903
rect 20916 31844 21404 31872
rect 20809 31807 20867 31813
rect 20809 31804 20821 31807
rect 20211 31776 20484 31804
rect 20548 31776 20821 31804
rect 20211 31773 20223 31776
rect 20165 31767 20223 31773
rect 14884 31708 15332 31736
rect 20456 31736 20484 31776
rect 20809 31773 20821 31776
rect 20855 31773 20867 31807
rect 20809 31767 20867 31773
rect 20898 31764 20904 31816
rect 20956 31804 20962 31816
rect 21376 31813 21404 31844
rect 21836 31813 21864 31912
rect 22066 31872 22094 31980
rect 23477 31977 23489 32011
rect 23523 32008 23535 32011
rect 24118 32008 24124 32020
rect 23523 31980 24124 32008
rect 23523 31977 23535 31980
rect 23477 31971 23535 31977
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 22066 31844 23888 31872
rect 21085 31807 21143 31813
rect 21085 31804 21097 31807
rect 20956 31776 21097 31804
rect 20956 31764 20962 31776
rect 21085 31773 21097 31776
rect 21131 31773 21143 31807
rect 21085 31767 21143 31773
rect 21361 31807 21419 31813
rect 21361 31773 21373 31807
rect 21407 31773 21419 31807
rect 21361 31767 21419 31773
rect 21821 31807 21879 31813
rect 21821 31773 21833 31807
rect 21867 31773 21879 31807
rect 21821 31767 21879 31773
rect 23198 31764 23204 31816
rect 23256 31804 23262 31816
rect 23860 31813 23888 31844
rect 23661 31807 23719 31813
rect 23661 31804 23673 31807
rect 23256 31776 23673 31804
rect 23256 31764 23262 31776
rect 23661 31773 23673 31776
rect 23707 31773 23719 31807
rect 23661 31767 23719 31773
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 24213 31807 24271 31813
rect 24213 31773 24225 31807
rect 24259 31804 24271 31807
rect 25130 31804 25136 31816
rect 24259 31776 25136 31804
rect 24259 31773 24271 31776
rect 24213 31767 24271 31773
rect 25130 31764 25136 31776
rect 25188 31764 25194 31816
rect 21542 31736 21548 31748
rect 20456 31708 21548 31736
rect 14884 31696 14890 31708
rect 21542 31696 21548 31708
rect 21600 31696 21606 31748
rect 22186 31696 22192 31748
rect 22244 31736 22250 31748
rect 22370 31736 22376 31748
rect 22244 31708 22376 31736
rect 22244 31696 22250 31708
rect 22370 31696 22376 31708
rect 22428 31696 22434 31748
rect 15746 31668 15752 31680
rect 14108 31640 15752 31668
rect 15746 31628 15752 31640
rect 15804 31628 15810 31680
rect 16022 31628 16028 31680
rect 16080 31668 16086 31680
rect 22094 31668 22100 31680
rect 16080 31640 22100 31668
rect 16080 31628 16086 31640
rect 22094 31628 22100 31640
rect 22152 31628 22158 31680
rect 1104 31578 25000 31600
rect 1104 31526 6884 31578
rect 6936 31526 6948 31578
rect 7000 31526 7012 31578
rect 7064 31526 7076 31578
rect 7128 31526 7140 31578
rect 7192 31526 12818 31578
rect 12870 31526 12882 31578
rect 12934 31526 12946 31578
rect 12998 31526 13010 31578
rect 13062 31526 13074 31578
rect 13126 31526 18752 31578
rect 18804 31526 18816 31578
rect 18868 31526 18880 31578
rect 18932 31526 18944 31578
rect 18996 31526 19008 31578
rect 19060 31526 24686 31578
rect 24738 31526 24750 31578
rect 24802 31526 24814 31578
rect 24866 31526 24878 31578
rect 24930 31526 24942 31578
rect 24994 31526 25000 31578
rect 1104 31504 25000 31526
rect 2498 31464 2504 31476
rect 1686 31436 2504 31464
rect 1686 31347 1714 31436
rect 2498 31424 2504 31436
rect 2556 31424 2562 31476
rect 3142 31424 3148 31476
rect 3200 31464 3206 31476
rect 3881 31467 3939 31473
rect 3881 31464 3893 31467
rect 3200 31436 3893 31464
rect 3200 31424 3206 31436
rect 3881 31433 3893 31436
rect 3927 31433 3939 31467
rect 5626 31464 5632 31476
rect 3881 31427 3939 31433
rect 4448 31436 5632 31464
rect 4154 31356 4160 31408
rect 4212 31356 4218 31408
rect 4448 31405 4476 31436
rect 5626 31424 5632 31436
rect 5684 31424 5690 31476
rect 5718 31424 5724 31476
rect 5776 31464 5782 31476
rect 5776 31436 7328 31464
rect 5776 31424 5782 31436
rect 4433 31399 4491 31405
rect 4433 31365 4445 31399
rect 4479 31365 4491 31399
rect 4433 31359 4491 31365
rect 4525 31399 4583 31405
rect 4525 31365 4537 31399
rect 4571 31396 4583 31399
rect 4614 31396 4620 31408
rect 4571 31368 4620 31396
rect 4571 31365 4583 31368
rect 4525 31359 4583 31365
rect 4614 31356 4620 31368
rect 4672 31356 4678 31408
rect 5261 31399 5319 31405
rect 5261 31396 5273 31399
rect 4816 31368 5273 31396
rect 1671 31341 1729 31347
rect 1671 31307 1683 31341
rect 1717 31307 1729 31341
rect 1671 31301 1729 31307
rect 3697 31331 3755 31337
rect 3697 31297 3709 31331
rect 3743 31328 3755 31331
rect 4816 31328 4844 31368
rect 5261 31365 5273 31368
rect 5307 31396 5319 31399
rect 5307 31368 5672 31396
rect 5307 31365 5319 31368
rect 5261 31359 5319 31365
rect 5644 31340 5672 31368
rect 5994 31356 6000 31408
rect 6052 31396 6058 31408
rect 7300 31405 7328 31436
rect 7650 31424 7656 31476
rect 7708 31424 7714 31476
rect 8665 31467 8723 31473
rect 8665 31433 8677 31467
rect 8711 31464 8723 31467
rect 15562 31464 15568 31476
rect 8711 31436 15568 31464
rect 8711 31433 8723 31436
rect 8665 31427 8723 31433
rect 6549 31399 6607 31405
rect 6549 31396 6561 31399
rect 6052 31368 6561 31396
rect 6052 31356 6058 31368
rect 6549 31365 6561 31368
rect 6595 31396 6607 31399
rect 7285 31399 7343 31405
rect 6595 31368 7236 31396
rect 6595 31365 6607 31368
rect 6549 31359 6607 31365
rect 3743 31300 4844 31328
rect 3743 31297 3755 31300
rect 3697 31291 3755 31297
rect 4890 31288 4896 31340
rect 4948 31288 4954 31340
rect 5626 31288 5632 31340
rect 5684 31288 5690 31340
rect 6178 31288 6184 31340
rect 6236 31328 6242 31340
rect 6638 31328 6644 31340
rect 6236 31300 6644 31328
rect 6236 31288 6242 31300
rect 6638 31288 6644 31300
rect 6696 31328 6702 31340
rect 6825 31331 6883 31337
rect 6825 31328 6837 31331
rect 6696 31300 6837 31328
rect 6696 31288 6702 31300
rect 6825 31297 6837 31300
rect 6871 31297 6883 31331
rect 6825 31291 6883 31297
rect 6917 31331 6975 31337
rect 6917 31297 6929 31331
rect 6963 31328 6975 31331
rect 7098 31328 7104 31340
rect 6963 31300 7104 31328
rect 6963 31297 6975 31300
rect 6917 31291 6975 31297
rect 7098 31288 7104 31300
rect 7156 31288 7162 31340
rect 7208 31328 7236 31368
rect 7285 31365 7297 31399
rect 7331 31365 7343 31399
rect 7285 31359 7343 31365
rect 8941 31399 8999 31405
rect 8941 31365 8953 31399
rect 8987 31396 8999 31399
rect 9306 31396 9312 31408
rect 8987 31368 9312 31396
rect 8987 31365 8999 31368
rect 8941 31359 8999 31365
rect 9306 31356 9312 31368
rect 9364 31356 9370 31408
rect 11146 31356 11152 31408
rect 11204 31396 11210 31408
rect 11606 31396 11612 31408
rect 11204 31368 11612 31396
rect 11204 31356 11210 31368
rect 11606 31356 11612 31368
rect 11664 31356 11670 31408
rect 12268 31405 12296 31436
rect 15562 31424 15568 31436
rect 15620 31424 15626 31476
rect 17218 31424 17224 31476
rect 17276 31464 17282 31476
rect 17954 31464 17960 31476
rect 17276 31436 17960 31464
rect 17276 31424 17282 31436
rect 17954 31424 17960 31436
rect 18012 31424 18018 31476
rect 12253 31399 12311 31405
rect 12253 31365 12265 31399
rect 12299 31365 12311 31399
rect 12253 31359 12311 31365
rect 12544 31368 13308 31396
rect 7926 31328 7932 31340
rect 7208 31300 7932 31328
rect 7926 31288 7932 31300
rect 7984 31288 7990 31340
rect 9030 31288 9036 31340
rect 9088 31288 9094 31340
rect 9398 31288 9404 31340
rect 9456 31288 9462 31340
rect 9766 31288 9772 31340
rect 9824 31337 9830 31340
rect 9824 31331 9841 31337
rect 9829 31297 9841 31331
rect 9824 31291 9841 31297
rect 9824 31288 9830 31291
rect 12434 31288 12440 31340
rect 12492 31328 12498 31340
rect 12544 31337 12572 31368
rect 13280 31340 13308 31368
rect 13464 31368 16620 31396
rect 12529 31331 12587 31337
rect 12529 31328 12541 31331
rect 12492 31300 12541 31328
rect 12492 31288 12498 31300
rect 12529 31297 12541 31300
rect 12575 31297 12587 31331
rect 12529 31291 12587 31297
rect 12802 31288 12808 31340
rect 12860 31328 12866 31340
rect 12860 31300 12903 31328
rect 12860 31288 12866 31300
rect 13262 31288 13268 31340
rect 13320 31288 13326 31340
rect 1394 31220 1400 31272
rect 1452 31220 1458 31272
rect 2777 31263 2835 31269
rect 2777 31229 2789 31263
rect 2823 31229 2835 31263
rect 2777 31223 2835 31229
rect 3053 31263 3111 31269
rect 3053 31229 3065 31263
rect 3099 31229 3111 31263
rect 3053 31223 3111 31229
rect 2792 31192 2820 31223
rect 2056 31164 2820 31192
rect 3068 31192 3096 31223
rect 3326 31220 3332 31272
rect 3384 31260 3390 31272
rect 3384 31232 4002 31260
rect 3384 31220 3390 31232
rect 6730 31220 6736 31272
rect 6788 31220 6794 31272
rect 9122 31220 9128 31272
rect 9180 31220 9186 31272
rect 3694 31192 3700 31204
rect 3068 31164 3700 31192
rect 1302 31084 1308 31136
rect 1360 31124 1366 31136
rect 2056 31124 2084 31164
rect 3694 31152 3700 31164
rect 3752 31152 3758 31204
rect 10410 31152 10416 31204
rect 10468 31192 10474 31204
rect 10686 31192 10692 31204
rect 10468 31164 10692 31192
rect 10468 31152 10474 31164
rect 10686 31152 10692 31164
rect 10744 31152 10750 31204
rect 12437 31195 12495 31201
rect 12437 31161 12449 31195
rect 12483 31161 12495 31195
rect 12437 31155 12495 31161
rect 1360 31096 2084 31124
rect 1360 31084 1366 31096
rect 2130 31084 2136 31136
rect 2188 31124 2194 31136
rect 2409 31127 2467 31133
rect 2409 31124 2421 31127
rect 2188 31096 2421 31124
rect 2188 31084 2194 31096
rect 2409 31093 2421 31096
rect 2455 31093 2467 31127
rect 2409 31087 2467 31093
rect 5445 31127 5503 31133
rect 5445 31093 5457 31127
rect 5491 31124 5503 31127
rect 6086 31124 6092 31136
rect 5491 31096 6092 31124
rect 5491 31093 5503 31096
rect 5445 31087 5503 31093
rect 6086 31084 6092 31096
rect 6144 31084 6150 31136
rect 7834 31084 7840 31136
rect 7892 31084 7898 31136
rect 8202 31084 8208 31136
rect 8260 31124 8266 31136
rect 8662 31124 8668 31136
rect 8260 31096 8668 31124
rect 8260 31084 8266 31096
rect 8662 31084 8668 31096
rect 8720 31084 8726 31136
rect 9953 31127 10011 31133
rect 9953 31093 9965 31127
rect 9999 31124 10011 31127
rect 10318 31124 10324 31136
rect 9999 31096 10324 31124
rect 9999 31093 10011 31096
rect 9953 31087 10011 31093
rect 10318 31084 10324 31096
rect 10376 31084 10382 31136
rect 11698 31084 11704 31136
rect 11756 31084 11762 31136
rect 12452 31124 12480 31155
rect 13262 31152 13268 31204
rect 13320 31192 13326 31204
rect 13464 31192 13492 31368
rect 13906 31328 13912 31340
rect 13556 31300 13912 31328
rect 13556 31201 13584 31300
rect 13906 31288 13912 31300
rect 13964 31288 13970 31340
rect 14093 31331 14151 31337
rect 14093 31297 14105 31331
rect 14139 31297 14151 31331
rect 14093 31291 14151 31297
rect 15379 31331 15437 31337
rect 15379 31297 15391 31331
rect 15425 31328 15437 31331
rect 15746 31328 15752 31340
rect 15425 31300 15752 31328
rect 15425 31297 15437 31300
rect 15379 31291 15437 31297
rect 13722 31220 13728 31272
rect 13780 31260 13786 31272
rect 14108 31260 14136 31291
rect 15746 31288 15752 31300
rect 15804 31328 15810 31340
rect 16482 31328 16488 31340
rect 15804 31300 16488 31328
rect 15804 31288 15810 31300
rect 16482 31288 16488 31300
rect 16540 31288 16546 31340
rect 16592 31328 16620 31368
rect 16942 31368 23336 31396
rect 16942 31337 16970 31368
rect 16911 31331 16970 31337
rect 16911 31328 16923 31331
rect 16592 31300 16923 31328
rect 16911 31297 16923 31300
rect 16957 31300 16970 31331
rect 16957 31297 16969 31300
rect 16911 31291 16969 31297
rect 17770 31288 17776 31340
rect 17828 31288 17834 31340
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18233 31331 18291 31337
rect 18233 31328 18245 31331
rect 18012 31300 18245 31328
rect 18012 31288 18018 31300
rect 18233 31297 18245 31300
rect 18279 31297 18291 31331
rect 18233 31291 18291 31297
rect 18509 31331 18567 31337
rect 18509 31297 18521 31331
rect 18555 31297 18567 31331
rect 18509 31291 18567 31297
rect 13780 31232 14136 31260
rect 15105 31263 15163 31269
rect 13780 31220 13786 31232
rect 15105 31229 15117 31263
rect 15151 31229 15163 31263
rect 15105 31223 15163 31229
rect 16669 31263 16727 31269
rect 16669 31229 16681 31263
rect 16715 31229 16727 31263
rect 16669 31223 16727 31229
rect 13320 31164 13492 31192
rect 13541 31195 13599 31201
rect 13320 31152 13326 31164
rect 13541 31161 13553 31195
rect 13587 31161 13599 31195
rect 13541 31155 13599 31161
rect 13722 31124 13728 31136
rect 12452 31096 13728 31124
rect 13722 31084 13728 31096
rect 13780 31084 13786 31136
rect 13998 31084 14004 31136
rect 14056 31084 14062 31136
rect 15120 31124 15148 31223
rect 16684 31192 16712 31223
rect 17788 31192 17816 31288
rect 18524 31260 18552 31291
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19763 31331 19821 31337
rect 19763 31328 19775 31331
rect 19484 31300 19775 31328
rect 19484 31288 19490 31300
rect 19763 31297 19775 31300
rect 19809 31297 19821 31331
rect 19763 31291 19821 31297
rect 21085 31331 21143 31337
rect 21085 31297 21097 31331
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 18064 31232 18552 31260
rect 18064 31201 18092 31232
rect 19334 31220 19340 31272
rect 19392 31260 19398 31272
rect 19521 31263 19579 31269
rect 19521 31260 19533 31263
rect 19392 31232 19533 31260
rect 19392 31220 19398 31232
rect 19521 31229 19533 31232
rect 19567 31229 19579 31263
rect 19521 31223 19579 31229
rect 20901 31263 20959 31269
rect 20901 31229 20913 31263
rect 20947 31229 20959 31263
rect 21100 31260 21128 31291
rect 21450 31288 21456 31340
rect 21508 31288 21514 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 22112 31300 22477 31328
rect 22112 31272 22140 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 23109 31331 23167 31337
rect 23109 31297 23121 31331
rect 23155 31297 23167 31331
rect 23109 31291 23167 31297
rect 21542 31260 21548 31272
rect 21100 31232 21548 31260
rect 20901 31223 20959 31229
rect 15764 31164 16804 31192
rect 15764 31124 15792 31164
rect 15120 31096 15792 31124
rect 16114 31084 16120 31136
rect 16172 31084 16178 31136
rect 16776 31124 16804 31164
rect 17328 31164 17816 31192
rect 18049 31195 18107 31201
rect 17126 31124 17132 31136
rect 16776 31096 17132 31124
rect 17126 31084 17132 31096
rect 17184 31124 17190 31136
rect 17328 31124 17356 31164
rect 18049 31161 18061 31195
rect 18095 31161 18107 31195
rect 18049 31155 18107 31161
rect 20533 31195 20591 31201
rect 20533 31161 20545 31195
rect 20579 31192 20591 31195
rect 20622 31192 20628 31204
rect 20579 31164 20628 31192
rect 20579 31161 20591 31164
rect 20533 31155 20591 31161
rect 20622 31152 20628 31164
rect 20680 31192 20686 31204
rect 20916 31192 20944 31223
rect 21542 31220 21548 31232
rect 21600 31220 21606 31272
rect 22094 31220 22100 31272
rect 22152 31220 22158 31272
rect 23124 31260 23152 31291
rect 23308 31272 23336 31368
rect 23753 31331 23811 31337
rect 23753 31328 23765 31331
rect 23400 31300 23765 31328
rect 22296 31232 23152 31260
rect 20680 31164 20944 31192
rect 20680 31152 20686 31164
rect 21082 31152 21088 31204
rect 21140 31152 21146 31204
rect 22296 31201 22324 31232
rect 23290 31220 23296 31272
rect 23348 31220 23354 31272
rect 22281 31195 22339 31201
rect 22281 31161 22293 31195
rect 22327 31161 22339 31195
rect 22281 31155 22339 31161
rect 22925 31195 22983 31201
rect 22925 31161 22937 31195
rect 22971 31192 22983 31195
rect 23400 31192 23428 31300
rect 23753 31297 23765 31300
rect 23799 31297 23811 31331
rect 23753 31291 23811 31297
rect 23842 31288 23848 31340
rect 23900 31328 23906 31340
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 23900 31300 24133 31328
rect 23900 31288 23906 31300
rect 24121 31297 24133 31300
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24213 31331 24271 31337
rect 24213 31297 24225 31331
rect 24259 31297 24271 31331
rect 24213 31291 24271 31297
rect 24228 31260 24256 31291
rect 23584 31232 24256 31260
rect 23584 31201 23612 31232
rect 22971 31164 23428 31192
rect 23569 31195 23627 31201
rect 22971 31161 22983 31164
rect 22925 31155 22983 31161
rect 23569 31161 23581 31195
rect 23615 31161 23627 31195
rect 23569 31155 23627 31161
rect 17184 31096 17356 31124
rect 17184 31084 17190 31096
rect 17402 31084 17408 31136
rect 17460 31124 17466 31136
rect 17681 31127 17739 31133
rect 17681 31124 17693 31127
rect 17460 31096 17693 31124
rect 17460 31084 17466 31096
rect 17681 31093 17693 31096
rect 17727 31093 17739 31127
rect 17681 31087 17739 31093
rect 18598 31084 18604 31136
rect 18656 31084 18662 31136
rect 23934 31084 23940 31136
rect 23992 31084 23998 31136
rect 24394 31084 24400 31136
rect 24452 31084 24458 31136
rect 1104 31034 24840 31056
rect 1104 30982 3917 31034
rect 3969 30982 3981 31034
rect 4033 30982 4045 31034
rect 4097 30982 4109 31034
rect 4161 30982 4173 31034
rect 4225 30982 9851 31034
rect 9903 30982 9915 31034
rect 9967 30982 9979 31034
rect 10031 30982 10043 31034
rect 10095 30982 10107 31034
rect 10159 30982 15785 31034
rect 15837 30982 15849 31034
rect 15901 30982 15913 31034
rect 15965 30982 15977 31034
rect 16029 30982 16041 31034
rect 16093 30982 21719 31034
rect 21771 30982 21783 31034
rect 21835 30982 21847 31034
rect 21899 30982 21911 31034
rect 21963 30982 21975 31034
rect 22027 30982 24840 31034
rect 1104 30960 24840 30982
rect 2424 30892 3004 30920
rect 1946 30812 1952 30864
rect 2004 30852 2010 30864
rect 2424 30852 2452 30892
rect 2004 30824 2452 30852
rect 2004 30812 2010 30824
rect 2332 30793 2360 30824
rect 2317 30787 2375 30793
rect 2317 30753 2329 30787
rect 2363 30753 2375 30787
rect 2976 30784 3004 30892
rect 3326 30880 3332 30932
rect 3384 30880 3390 30932
rect 4614 30880 4620 30932
rect 4672 30920 4678 30932
rect 5261 30923 5319 30929
rect 5261 30920 5273 30923
rect 4672 30892 5273 30920
rect 4672 30880 4678 30892
rect 5261 30889 5273 30892
rect 5307 30889 5319 30923
rect 5261 30883 5319 30889
rect 6086 30880 6092 30932
rect 6144 30920 6150 30932
rect 6638 30920 6644 30932
rect 6144 30892 6644 30920
rect 6144 30880 6150 30892
rect 6638 30880 6644 30892
rect 6696 30880 6702 30932
rect 7098 30880 7104 30932
rect 7156 30920 7162 30932
rect 7377 30923 7435 30929
rect 7377 30920 7389 30923
rect 7156 30892 7389 30920
rect 7156 30880 7162 30892
rect 7377 30889 7389 30892
rect 7423 30889 7435 30923
rect 7377 30883 7435 30889
rect 9030 30880 9036 30932
rect 9088 30920 9094 30932
rect 9953 30923 10011 30929
rect 9953 30920 9965 30923
rect 9088 30892 9965 30920
rect 9088 30880 9094 30892
rect 9953 30889 9965 30892
rect 9999 30889 10011 30923
rect 9953 30883 10011 30889
rect 10612 30892 12480 30920
rect 10612 30852 10640 30892
rect 10962 30852 10968 30864
rect 9646 30824 10640 30852
rect 10704 30824 10968 30852
rect 4249 30787 4307 30793
rect 4249 30784 4261 30787
rect 2976 30756 4261 30784
rect 2317 30747 2375 30753
rect 4249 30753 4261 30756
rect 4295 30753 4307 30787
rect 4249 30747 4307 30753
rect 2590 30716 2596 30728
rect 2551 30688 2596 30716
rect 2590 30676 2596 30688
rect 2648 30676 2654 30728
rect 3786 30676 3792 30728
rect 3844 30676 3850 30728
rect 4154 30676 4160 30728
rect 4212 30716 4218 30728
rect 4264 30716 4292 30747
rect 5810 30744 5816 30796
rect 5868 30784 5874 30796
rect 6362 30784 6368 30796
rect 5868 30756 6368 30784
rect 5868 30744 5874 30756
rect 6362 30744 6368 30756
rect 6420 30744 6426 30796
rect 8570 30744 8576 30796
rect 8628 30784 8634 30796
rect 8941 30787 8999 30793
rect 8941 30784 8953 30787
rect 8628 30756 8953 30784
rect 8628 30744 8634 30756
rect 8941 30753 8953 30756
rect 8987 30753 8999 30787
rect 8941 30747 8999 30753
rect 4522 30716 4528 30728
rect 4212 30688 4292 30716
rect 4483 30688 4528 30716
rect 4212 30676 4218 30688
rect 4522 30676 4528 30688
rect 4580 30676 4586 30728
rect 4614 30676 4620 30728
rect 4672 30716 4678 30728
rect 5074 30716 5080 30728
rect 4672 30688 5080 30716
rect 4672 30676 4678 30688
rect 5074 30676 5080 30688
rect 5132 30676 5138 30728
rect 6546 30676 6552 30728
rect 6604 30716 6610 30728
rect 6639 30719 6697 30725
rect 6639 30716 6651 30719
rect 6604 30688 6651 30716
rect 6604 30676 6610 30688
rect 6639 30685 6651 30688
rect 6685 30685 6697 30719
rect 9214 30716 9220 30728
rect 9175 30688 9220 30716
rect 6639 30679 6697 30685
rect 9214 30676 9220 30688
rect 9272 30676 9278 30728
rect 1486 30608 1492 30660
rect 1544 30608 1550 30660
rect 1673 30651 1731 30657
rect 1673 30617 1685 30651
rect 1719 30648 1731 30651
rect 4246 30648 4252 30660
rect 1719 30620 4252 30648
rect 1719 30617 1731 30620
rect 1673 30611 1731 30617
rect 4246 30608 4252 30620
rect 4304 30608 4310 30660
rect 7282 30608 7288 30660
rect 7340 30648 7346 30660
rect 8110 30648 8116 30660
rect 7340 30620 8116 30648
rect 7340 30608 7346 30620
rect 8110 30608 8116 30620
rect 8168 30648 8174 30660
rect 9646 30648 9674 30824
rect 10704 30728 10732 30824
rect 10962 30812 10968 30824
rect 11020 30812 11026 30864
rect 12452 30852 12480 30892
rect 12526 30880 12532 30932
rect 12584 30880 12590 30932
rect 12805 30923 12863 30929
rect 12805 30889 12817 30923
rect 12851 30920 12863 30923
rect 13630 30920 13636 30932
rect 12851 30892 13636 30920
rect 12851 30889 12863 30892
rect 12805 30883 12863 30889
rect 13630 30880 13636 30892
rect 13688 30880 13694 30932
rect 13998 30880 14004 30932
rect 14056 30880 14062 30932
rect 16114 30880 16120 30932
rect 16172 30880 16178 30932
rect 17402 30880 17408 30932
rect 17460 30880 17466 30932
rect 17589 30923 17647 30929
rect 17589 30889 17601 30923
rect 17635 30920 17647 30923
rect 17954 30920 17960 30932
rect 17635 30892 17960 30920
rect 17635 30889 17647 30892
rect 17589 30883 17647 30889
rect 13170 30852 13176 30864
rect 12452 30824 13176 30852
rect 13170 30812 13176 30824
rect 13228 30812 13234 30864
rect 11146 30744 11152 30796
rect 11204 30744 11210 30796
rect 11238 30744 11244 30796
rect 11296 30784 11302 30796
rect 11425 30787 11483 30793
rect 11425 30784 11437 30787
rect 11296 30756 11437 30784
rect 11296 30744 11302 30756
rect 11425 30753 11437 30756
rect 11471 30753 11483 30787
rect 11425 30747 11483 30753
rect 11514 30744 11520 30796
rect 11572 30793 11578 30796
rect 11572 30787 11600 30793
rect 11588 30753 11600 30787
rect 11572 30747 11600 30753
rect 11701 30787 11759 30793
rect 11701 30753 11713 30787
rect 11747 30784 11759 30787
rect 12066 30784 12072 30796
rect 11747 30756 12072 30784
rect 11747 30753 11759 30756
rect 11701 30747 11759 30753
rect 11572 30744 11578 30747
rect 12066 30744 12072 30756
rect 12124 30744 12130 30796
rect 13906 30744 13912 30796
rect 13964 30744 13970 30796
rect 14016 30784 14044 30880
rect 14826 30812 14832 30864
rect 14884 30852 14890 30864
rect 16132 30852 16160 30880
rect 16393 30855 16451 30861
rect 16393 30852 16405 30855
rect 14884 30824 16068 30852
rect 16132 30824 16405 30852
rect 14884 30812 14890 30824
rect 14016 30756 14964 30784
rect 9766 30676 9772 30728
rect 9824 30716 9830 30728
rect 10505 30719 10563 30725
rect 10505 30716 10517 30719
rect 9824 30688 10517 30716
rect 9824 30676 9830 30688
rect 10505 30685 10517 30688
rect 10551 30685 10563 30719
rect 10505 30679 10563 30685
rect 10686 30676 10692 30728
rect 10744 30676 10750 30728
rect 12345 30719 12403 30725
rect 12345 30685 12357 30719
rect 12391 30716 12403 30719
rect 12713 30719 12771 30725
rect 12713 30716 12725 30719
rect 12391 30688 12725 30716
rect 12391 30685 12403 30688
rect 12345 30679 12403 30685
rect 12713 30685 12725 30688
rect 12759 30685 12771 30719
rect 12713 30679 12771 30685
rect 12989 30719 13047 30725
rect 12989 30685 13001 30719
rect 13035 30685 13047 30719
rect 13924 30716 13952 30744
rect 14936 30725 14964 30756
rect 15470 30744 15476 30796
rect 15528 30784 15534 30796
rect 16040 30784 16068 30824
rect 16393 30821 16405 30824
rect 16439 30821 16451 30855
rect 16393 30815 16451 30821
rect 16786 30787 16844 30793
rect 16786 30784 16798 30787
rect 15528 30756 15976 30784
rect 16040 30756 16798 30784
rect 15528 30744 15534 30756
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 13924 30688 14105 30716
rect 12989 30679 13047 30685
rect 14093 30685 14105 30688
rect 14139 30685 14151 30719
rect 14093 30679 14151 30685
rect 14461 30719 14519 30725
rect 14461 30685 14473 30719
rect 14507 30685 14519 30719
rect 14461 30679 14519 30685
rect 14921 30719 14979 30725
rect 14921 30685 14933 30719
rect 14967 30685 14979 30719
rect 14921 30679 14979 30685
rect 8168 30620 9674 30648
rect 8168 30608 8174 30620
rect 566 30540 572 30592
rect 624 30580 630 30592
rect 1578 30580 1584 30592
rect 624 30552 1584 30580
rect 624 30540 630 30552
rect 1578 30540 1584 30552
rect 1636 30540 1642 30592
rect 3973 30583 4031 30589
rect 3973 30549 3985 30583
rect 4019 30580 4031 30583
rect 4522 30580 4528 30592
rect 4019 30552 4528 30580
rect 4019 30549 4031 30552
rect 3973 30543 4031 30549
rect 4522 30540 4528 30552
rect 4580 30580 4586 30592
rect 5258 30580 5264 30592
rect 4580 30552 5264 30580
rect 4580 30540 4586 30552
rect 5258 30540 5264 30552
rect 5316 30540 5322 30592
rect 7466 30540 7472 30592
rect 7524 30580 7530 30592
rect 11514 30580 11520 30592
rect 7524 30552 11520 30580
rect 7524 30540 7530 30552
rect 11514 30540 11520 30552
rect 11572 30540 11578 30592
rect 12342 30540 12348 30592
rect 12400 30580 12406 30592
rect 13004 30580 13032 30679
rect 13814 30608 13820 30660
rect 13872 30648 13878 30660
rect 14476 30648 14504 30679
rect 15562 30676 15568 30728
rect 15620 30716 15626 30728
rect 15948 30725 15976 30756
rect 16786 30753 16798 30756
rect 16832 30753 16844 30787
rect 16786 30747 16844 30753
rect 16945 30787 17003 30793
rect 16945 30753 16957 30787
rect 16991 30784 17003 30787
rect 17420 30784 17448 30880
rect 16991 30756 17448 30784
rect 16991 30753 17003 30756
rect 16945 30747 17003 30753
rect 15749 30719 15807 30725
rect 15749 30716 15761 30719
rect 15620 30688 15761 30716
rect 15620 30676 15626 30688
rect 15749 30685 15761 30688
rect 15795 30685 15807 30719
rect 15749 30679 15807 30685
rect 15933 30719 15991 30725
rect 15933 30685 15945 30719
rect 15979 30716 15991 30719
rect 16114 30716 16120 30728
rect 15979 30688 16120 30716
rect 15979 30685 15991 30688
rect 15933 30679 15991 30685
rect 16114 30676 16120 30688
rect 16172 30676 16178 30728
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 17604 30716 17632 30883
rect 17954 30880 17960 30892
rect 18012 30880 18018 30932
rect 18598 30880 18604 30932
rect 18656 30920 18662 30932
rect 19337 30923 19395 30929
rect 19337 30920 19349 30923
rect 18656 30892 19349 30920
rect 18656 30880 18662 30892
rect 19337 30889 19349 30892
rect 19383 30889 19395 30923
rect 19337 30883 19395 30889
rect 19812 30892 20116 30920
rect 19061 30855 19119 30861
rect 19061 30821 19073 30855
rect 19107 30852 19119 30855
rect 19812 30852 19840 30892
rect 19107 30824 19840 30852
rect 19889 30855 19947 30861
rect 19107 30821 19119 30824
rect 19061 30815 19119 30821
rect 19889 30821 19901 30855
rect 19935 30821 19947 30855
rect 19889 30815 19947 30821
rect 17678 30744 17684 30796
rect 17736 30744 17742 30796
rect 19521 30787 19579 30793
rect 19521 30753 19533 30787
rect 19567 30784 19579 30787
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19567 30756 19717 30784
rect 19567 30753 19579 30756
rect 19521 30747 19579 30753
rect 19705 30753 19717 30756
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 17937 30719 17995 30725
rect 17937 30716 17949 30719
rect 17604 30688 17949 30716
rect 17937 30685 17949 30688
rect 17983 30685 17995 30719
rect 17937 30679 17995 30685
rect 19245 30719 19303 30725
rect 19245 30685 19257 30719
rect 19291 30716 19303 30719
rect 19613 30719 19671 30725
rect 19613 30716 19625 30719
rect 19291 30688 19625 30716
rect 19291 30685 19303 30688
rect 19245 30679 19303 30685
rect 19613 30685 19625 30688
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 19904 30716 19932 30815
rect 20088 30725 20116 30892
rect 20622 30880 20628 30932
rect 20680 30880 20686 30932
rect 20717 30923 20775 30929
rect 20717 30889 20729 30923
rect 20763 30920 20775 30923
rect 21450 30920 21456 30932
rect 20763 30892 21456 30920
rect 20763 30889 20775 30892
rect 20717 30883 20775 30889
rect 21450 30880 21456 30892
rect 21508 30880 21514 30932
rect 23109 30923 23167 30929
rect 23109 30889 23121 30923
rect 23155 30920 23167 30923
rect 23155 30892 23704 30920
rect 23155 30889 23167 30892
rect 23109 30883 23167 30889
rect 20640 30725 20668 30880
rect 22833 30855 22891 30861
rect 22833 30821 22845 30855
rect 22879 30821 22891 30855
rect 22833 30815 22891 30821
rect 23477 30855 23535 30861
rect 23477 30821 23489 30855
rect 23523 30821 23535 30855
rect 23477 30815 23535 30821
rect 19843 30688 19932 30716
rect 20073 30719 20131 30725
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 20073 30685 20085 30719
rect 20119 30685 20131 30719
rect 20073 30679 20131 30685
rect 20625 30719 20683 30725
rect 20625 30685 20637 30719
rect 20671 30685 20683 30719
rect 20625 30679 20683 30685
rect 13872 30620 14504 30648
rect 15197 30651 15255 30657
rect 13872 30608 13878 30620
rect 15197 30617 15209 30651
rect 15243 30617 15255 30651
rect 15197 30611 15255 30617
rect 12400 30552 13032 30580
rect 15212 30580 15240 30611
rect 19260 30592 19288 30679
rect 20806 30676 20812 30728
rect 20864 30676 20870 30728
rect 22278 30676 22284 30728
rect 22336 30676 22342 30728
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30648 19579 30651
rect 22848 30648 22876 30815
rect 23492 30784 23520 30815
rect 23032 30756 23520 30784
rect 23032 30725 23060 30756
rect 23017 30719 23075 30725
rect 23017 30685 23029 30719
rect 23063 30685 23075 30719
rect 23017 30679 23075 30685
rect 23290 30676 23296 30728
rect 23348 30676 23354 30728
rect 23676 30725 23704 30892
rect 23661 30719 23719 30725
rect 23661 30685 23673 30719
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 23845 30651 23903 30657
rect 23845 30648 23857 30651
rect 19567 30620 22784 30648
rect 22848 30620 23857 30648
rect 19567 30617 19579 30620
rect 19521 30611 19579 30617
rect 16390 30580 16396 30592
rect 15212 30552 16396 30580
rect 12400 30540 12406 30552
rect 16390 30540 16396 30552
rect 16448 30540 16454 30592
rect 19242 30540 19248 30592
rect 19300 30540 19306 30592
rect 22097 30583 22155 30589
rect 22097 30549 22109 30583
rect 22143 30580 22155 30583
rect 22554 30580 22560 30592
rect 22143 30552 22560 30580
rect 22143 30549 22155 30552
rect 22097 30543 22155 30549
rect 22554 30540 22560 30552
rect 22612 30540 22618 30592
rect 22756 30580 22784 30620
rect 23845 30617 23857 30620
rect 23891 30617 23903 30651
rect 23845 30611 23903 30617
rect 24213 30651 24271 30657
rect 24213 30617 24225 30651
rect 24259 30648 24271 30651
rect 25130 30648 25136 30660
rect 24259 30620 25136 30648
rect 24259 30617 24271 30620
rect 24213 30611 24271 30617
rect 25130 30608 25136 30620
rect 25188 30608 25194 30660
rect 25682 30608 25688 30660
rect 25740 30608 25746 30660
rect 25700 30580 25728 30608
rect 22756 30552 25728 30580
rect 1104 30490 25000 30512
rect 1104 30438 6884 30490
rect 6936 30438 6948 30490
rect 7000 30438 7012 30490
rect 7064 30438 7076 30490
rect 7128 30438 7140 30490
rect 7192 30438 12818 30490
rect 12870 30438 12882 30490
rect 12934 30438 12946 30490
rect 12998 30438 13010 30490
rect 13062 30438 13074 30490
rect 13126 30438 18752 30490
rect 18804 30438 18816 30490
rect 18868 30438 18880 30490
rect 18932 30438 18944 30490
rect 18996 30438 19008 30490
rect 19060 30438 24686 30490
rect 24738 30438 24750 30490
rect 24802 30438 24814 30490
rect 24866 30438 24878 30490
rect 24930 30438 24942 30490
rect 24994 30438 25000 30490
rect 1104 30416 25000 30438
rect 658 30336 664 30388
rect 716 30376 722 30388
rect 716 30348 3372 30376
rect 716 30336 722 30348
rect 3344 30317 3372 30348
rect 3694 30336 3700 30388
rect 3752 30376 3758 30388
rect 10965 30379 11023 30385
rect 3752 30348 10916 30376
rect 3752 30336 3758 30348
rect 3329 30311 3387 30317
rect 3329 30277 3341 30311
rect 3375 30277 3387 30311
rect 4706 30308 4712 30320
rect 4446 30280 4712 30308
rect 4446 30279 4474 30280
rect 3329 30271 3387 30277
rect 4415 30273 4474 30279
rect 2682 30200 2688 30252
rect 2740 30200 2746 30252
rect 3418 30200 3424 30252
rect 3476 30200 3482 30252
rect 4415 30239 4427 30273
rect 4461 30242 4474 30273
rect 4706 30268 4712 30280
rect 4764 30308 4770 30320
rect 5902 30308 5908 30320
rect 4764 30280 5908 30308
rect 4764 30268 4770 30280
rect 5902 30268 5908 30280
rect 5960 30268 5966 30320
rect 6822 30268 6828 30320
rect 6880 30308 6886 30320
rect 10888 30308 10916 30348
rect 10965 30345 10977 30379
rect 11011 30376 11023 30379
rect 11146 30376 11152 30388
rect 11011 30348 11152 30376
rect 11011 30345 11023 30348
rect 10965 30339 11023 30345
rect 11146 30336 11152 30348
rect 11204 30336 11210 30388
rect 13906 30336 13912 30388
rect 13964 30376 13970 30388
rect 14366 30376 14372 30388
rect 13964 30348 14372 30376
rect 13964 30336 13970 30348
rect 14366 30336 14372 30348
rect 14424 30336 14430 30388
rect 18969 30379 19027 30385
rect 18156 30348 18368 30376
rect 13998 30308 14004 30320
rect 6880 30280 10824 30308
rect 10888 30280 14004 30308
rect 6880 30268 6886 30280
rect 7099 30243 7157 30249
rect 4461 30239 4473 30242
rect 4415 30233 4473 30239
rect 7099 30209 7111 30243
rect 7145 30240 7157 30243
rect 7558 30240 7564 30252
rect 7145 30212 7564 30240
rect 7145 30209 7157 30212
rect 7099 30203 7157 30209
rect 7558 30200 7564 30212
rect 7616 30240 7622 30252
rect 8018 30240 8024 30252
rect 7616 30212 8024 30240
rect 7616 30200 7622 30212
rect 8018 30200 8024 30212
rect 8076 30200 8082 30252
rect 10134 30200 10140 30252
rect 10192 30240 10198 30252
rect 10227 30243 10285 30249
rect 10227 30240 10239 30243
rect 10192 30212 10239 30240
rect 10192 30200 10198 30212
rect 10227 30209 10239 30212
rect 10273 30209 10285 30243
rect 10227 30203 10285 30209
rect 1489 30175 1547 30181
rect 1489 30141 1501 30175
rect 1535 30141 1547 30175
rect 1489 30135 1547 30141
rect 1504 30104 1532 30135
rect 1670 30132 1676 30184
rect 1728 30132 1734 30184
rect 2130 30132 2136 30184
rect 2188 30132 2194 30184
rect 2222 30132 2228 30184
rect 2280 30172 2286 30184
rect 2590 30181 2596 30184
rect 2409 30175 2467 30181
rect 2409 30172 2421 30175
rect 2280 30144 2421 30172
rect 2280 30132 2286 30144
rect 2409 30141 2421 30144
rect 2455 30141 2467 30175
rect 2409 30135 2467 30141
rect 2547 30175 2596 30181
rect 2547 30141 2559 30175
rect 2593 30141 2596 30175
rect 2547 30135 2596 30141
rect 2590 30132 2596 30135
rect 2648 30132 2654 30184
rect 4154 30132 4160 30184
rect 4212 30132 4218 30184
rect 5074 30132 5080 30184
rect 5132 30172 5138 30184
rect 5442 30172 5448 30184
rect 5132 30144 5448 30172
rect 5132 30132 5138 30144
rect 5442 30132 5448 30144
rect 5500 30132 5506 30184
rect 5534 30132 5540 30184
rect 5592 30172 5598 30184
rect 5902 30172 5908 30184
rect 5592 30144 5908 30172
rect 5592 30132 5598 30144
rect 5902 30132 5908 30144
rect 5960 30172 5966 30184
rect 6730 30172 6736 30184
rect 5960 30144 6736 30172
rect 5960 30132 5966 30144
rect 6730 30132 6736 30144
rect 6788 30132 6794 30184
rect 6825 30175 6883 30181
rect 6825 30141 6837 30175
rect 6871 30141 6883 30175
rect 6825 30135 6883 30141
rect 9953 30175 10011 30181
rect 9953 30141 9965 30175
rect 9999 30141 10011 30175
rect 10796 30172 10824 30280
rect 13998 30268 14004 30280
rect 14056 30308 14062 30320
rect 14826 30308 14832 30320
rect 14056 30280 14832 30308
rect 14056 30268 14062 30280
rect 14826 30268 14832 30280
rect 14884 30268 14890 30320
rect 15010 30268 15016 30320
rect 15068 30308 15074 30320
rect 17954 30308 17960 30320
rect 15068 30280 17960 30308
rect 15068 30268 15074 30280
rect 17954 30268 17960 30280
rect 18012 30268 18018 30320
rect 11238 30200 11244 30252
rect 11296 30240 11302 30252
rect 14183 30243 14241 30249
rect 14183 30240 14195 30243
rect 11296 30212 14195 30240
rect 11296 30200 11302 30212
rect 14183 30209 14195 30212
rect 14229 30240 14241 30243
rect 14229 30212 16252 30240
rect 14229 30209 14241 30212
rect 14183 30203 14241 30209
rect 10796 30144 13860 30172
rect 9953 30135 10011 30141
rect 1946 30104 1952 30116
rect 1504 30076 1952 30104
rect 1946 30064 1952 30076
rect 2004 30064 2010 30116
rect 5994 30104 6000 30116
rect 5092 30076 6000 30104
rect 3605 30039 3663 30045
rect 3605 30005 3617 30039
rect 3651 30036 3663 30039
rect 5092 30036 5120 30076
rect 5994 30064 6000 30076
rect 6052 30064 6058 30116
rect 6362 30064 6368 30116
rect 6420 30064 6426 30116
rect 6454 30064 6460 30116
rect 6512 30104 6518 30116
rect 6840 30104 6868 30135
rect 9030 30104 9036 30116
rect 6512 30076 6868 30104
rect 7760 30076 9036 30104
rect 6512 30064 6518 30076
rect 3651 30008 5120 30036
rect 3651 30005 3663 30008
rect 3605 29999 3663 30005
rect 5166 29996 5172 30048
rect 5224 29996 5230 30048
rect 6380 30036 6408 30064
rect 7760 30036 7788 30076
rect 9030 30064 9036 30076
rect 9088 30064 9094 30116
rect 6380 30008 7788 30036
rect 7834 29996 7840 30048
rect 7892 29996 7898 30048
rect 9968 30036 9996 30135
rect 13832 30104 13860 30144
rect 13906 30132 13912 30184
rect 13964 30132 13970 30184
rect 16224 30104 16252 30212
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 18156 30240 18184 30348
rect 18340 30308 18368 30348
rect 18969 30345 18981 30379
rect 19015 30376 19027 30379
rect 19242 30376 19248 30388
rect 19015 30348 19248 30376
rect 19015 30345 19027 30348
rect 18969 30339 19027 30345
rect 19242 30336 19248 30348
rect 19300 30336 19306 30388
rect 23753 30379 23811 30385
rect 23753 30345 23765 30379
rect 23799 30376 23811 30379
rect 23842 30376 23848 30388
rect 23799 30348 23848 30376
rect 23799 30345 23811 30348
rect 23753 30339 23811 30345
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 23992 30348 24164 30376
rect 23992 30336 23998 30348
rect 24136 30317 24164 30348
rect 24121 30311 24179 30317
rect 18340 30280 23704 30308
rect 16540 30212 18184 30240
rect 18231 30243 18289 30249
rect 16540 30200 16546 30212
rect 18231 30209 18243 30243
rect 18277 30240 18289 30243
rect 19058 30240 19064 30252
rect 18277 30212 19064 30240
rect 18277 30209 18289 30212
rect 18231 30203 18289 30209
rect 19058 30200 19064 30212
rect 19116 30200 19122 30252
rect 20530 30249 20536 30252
rect 20513 30243 20536 30249
rect 20513 30240 20525 30243
rect 19168 30212 20525 30240
rect 17586 30132 17592 30184
rect 17644 30172 17650 30184
rect 17862 30172 17868 30184
rect 17644 30144 17868 30172
rect 17644 30132 17650 30144
rect 17862 30132 17868 30144
rect 17920 30172 17926 30184
rect 17957 30175 18015 30181
rect 17957 30172 17969 30175
rect 17920 30144 17969 30172
rect 17920 30132 17926 30144
rect 17957 30141 17969 30144
rect 18003 30141 18015 30175
rect 17957 30135 18015 30141
rect 13832 30076 14044 30104
rect 16224 30076 17816 30104
rect 12434 30036 12440 30048
rect 9968 30008 12440 30036
rect 12434 29996 12440 30008
rect 12492 30036 12498 30048
rect 13814 30036 13820 30048
rect 12492 30008 13820 30036
rect 12492 29996 12498 30008
rect 13814 29996 13820 30008
rect 13872 29996 13878 30048
rect 14016 30036 14044 30076
rect 17788 30048 17816 30076
rect 14826 30036 14832 30048
rect 14016 30008 14832 30036
rect 14826 29996 14832 30008
rect 14884 29996 14890 30048
rect 14918 29996 14924 30048
rect 14976 29996 14982 30048
rect 17770 29996 17776 30048
rect 17828 29996 17834 30048
rect 18230 29996 18236 30048
rect 18288 30036 18294 30048
rect 19168 30036 19196 30212
rect 20513 30209 20525 30212
rect 20513 30203 20536 30209
rect 20530 30200 20536 30203
rect 20588 30200 20594 30252
rect 22094 30200 22100 30252
rect 22152 30200 22158 30252
rect 23290 30200 23296 30252
rect 23348 30240 23354 30252
rect 23676 30249 23704 30280
rect 24121 30277 24133 30311
rect 24167 30277 24179 30311
rect 24121 30271 24179 30277
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 23348 30212 23397 30240
rect 23348 30200 23354 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 23661 30243 23719 30249
rect 23661 30209 23673 30243
rect 23707 30209 23719 30243
rect 23661 30203 23719 30209
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 19426 30132 19432 30184
rect 19484 30172 19490 30184
rect 20257 30175 20315 30181
rect 20257 30172 20269 30175
rect 19484 30144 20269 30172
rect 19484 30132 19490 30144
rect 20257 30141 20269 30144
rect 20303 30141 20315 30175
rect 21821 30175 21879 30181
rect 21821 30172 21833 30175
rect 20257 30135 20315 30141
rect 21284 30144 21833 30172
rect 18288 30008 19196 30036
rect 18288 29996 18294 30008
rect 19978 29996 19984 30048
rect 20036 30036 20042 30048
rect 21284 30036 21312 30144
rect 21821 30141 21833 30144
rect 21867 30141 21879 30175
rect 23952 30172 23980 30203
rect 21821 30135 21879 30141
rect 23492 30144 23980 30172
rect 23492 30113 23520 30144
rect 23477 30107 23535 30113
rect 23477 30073 23489 30107
rect 23523 30073 23535 30107
rect 23477 30067 23535 30073
rect 20036 30008 21312 30036
rect 21637 30039 21695 30045
rect 20036 29996 20042 30008
rect 21637 30005 21649 30039
rect 21683 30036 21695 30039
rect 22278 30036 22284 30048
rect 21683 30008 22284 30036
rect 21683 30005 21695 30008
rect 21637 29999 21695 30005
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 22830 29996 22836 30048
rect 22888 29996 22894 30048
rect 23198 29996 23204 30048
rect 23256 29996 23262 30048
rect 24394 29996 24400 30048
rect 24452 29996 24458 30048
rect 1104 29946 24840 29968
rect 1104 29894 3917 29946
rect 3969 29894 3981 29946
rect 4033 29894 4045 29946
rect 4097 29894 4109 29946
rect 4161 29894 4173 29946
rect 4225 29894 9851 29946
rect 9903 29894 9915 29946
rect 9967 29894 9979 29946
rect 10031 29894 10043 29946
rect 10095 29894 10107 29946
rect 10159 29894 15785 29946
rect 15837 29894 15849 29946
rect 15901 29894 15913 29946
rect 15965 29894 15977 29946
rect 16029 29894 16041 29946
rect 16093 29894 21719 29946
rect 21771 29894 21783 29946
rect 21835 29894 21847 29946
rect 21899 29894 21911 29946
rect 21963 29894 21975 29946
rect 22027 29894 24840 29946
rect 1104 29872 24840 29894
rect 1118 29792 1124 29844
rect 1176 29832 1182 29844
rect 1176 29804 2360 29832
rect 1176 29792 1182 29804
rect 1578 29724 1584 29776
rect 1636 29724 1642 29776
rect 2332 29764 2360 29804
rect 2682 29792 2688 29844
rect 2740 29792 2746 29844
rect 2774 29792 2780 29844
rect 2832 29832 2838 29844
rect 2832 29804 2912 29832
rect 2832 29792 2838 29804
rect 2884 29764 2912 29804
rect 3050 29792 3056 29844
rect 3108 29832 3114 29844
rect 3237 29835 3295 29841
rect 3237 29832 3249 29835
rect 3108 29804 3249 29832
rect 3108 29792 3114 29804
rect 3237 29801 3249 29804
rect 3283 29801 3295 29835
rect 3237 29795 3295 29801
rect 3602 29792 3608 29844
rect 3660 29792 3666 29844
rect 6178 29792 6184 29844
rect 6236 29832 6242 29844
rect 6273 29835 6331 29841
rect 6273 29832 6285 29835
rect 6236 29804 6285 29832
rect 6236 29792 6242 29804
rect 6273 29801 6285 29804
rect 6319 29801 6331 29835
rect 6273 29795 6331 29801
rect 7466 29792 7472 29844
rect 7524 29792 7530 29844
rect 7834 29832 7840 29844
rect 7576 29804 7840 29832
rect 7098 29764 7104 29776
rect 2332 29736 2774 29764
rect 2884 29736 4108 29764
rect 2746 29696 2774 29736
rect 3789 29699 3847 29705
rect 3789 29696 3801 29699
rect 2746 29668 3801 29696
rect 3789 29665 3801 29668
rect 3835 29665 3847 29699
rect 3789 29659 3847 29665
rect 1394 29588 1400 29640
rect 1452 29588 1458 29640
rect 1486 29588 1492 29640
rect 1544 29628 1550 29640
rect 1673 29631 1731 29637
rect 1673 29628 1685 29631
rect 1544 29600 1685 29628
rect 1544 29588 1550 29600
rect 1673 29597 1685 29600
rect 1719 29628 1731 29631
rect 1854 29628 1860 29640
rect 1719 29600 1860 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 1854 29588 1860 29600
rect 1912 29588 1918 29640
rect 1947 29631 2005 29637
rect 1947 29597 1959 29631
rect 1993 29628 2005 29631
rect 2406 29628 2412 29640
rect 1993 29600 2412 29628
rect 1993 29597 2005 29600
rect 1947 29591 2005 29597
rect 2406 29588 2412 29600
rect 2464 29588 2470 29640
rect 3053 29631 3111 29637
rect 3053 29628 3065 29631
rect 2746 29600 3065 29628
rect 1302 29520 1308 29572
rect 1360 29560 1366 29572
rect 2746 29560 2774 29600
rect 3053 29597 3065 29600
rect 3099 29597 3111 29631
rect 3053 29591 3111 29597
rect 3421 29631 3479 29637
rect 3421 29597 3433 29631
rect 3467 29628 3479 29631
rect 3602 29628 3608 29640
rect 3467 29600 3608 29628
rect 3467 29597 3479 29600
rect 3421 29591 3479 29597
rect 3602 29588 3608 29600
rect 3660 29588 3666 29640
rect 4080 29637 4108 29736
rect 6104 29736 7104 29764
rect 6104 29708 6132 29736
rect 7098 29724 7104 29736
rect 7156 29724 7162 29776
rect 5166 29656 5172 29708
rect 5224 29656 5230 29708
rect 6086 29656 6092 29708
rect 6144 29656 6150 29708
rect 7484 29696 7512 29792
rect 7576 29773 7604 29804
rect 7834 29792 7840 29804
rect 7892 29792 7898 29844
rect 8754 29792 8760 29844
rect 8812 29792 8818 29844
rect 9030 29792 9036 29844
rect 9088 29832 9094 29844
rect 9088 29804 12112 29832
rect 9088 29792 9094 29804
rect 7561 29767 7619 29773
rect 7561 29733 7573 29767
rect 7607 29733 7619 29767
rect 7561 29727 7619 29733
rect 10502 29724 10508 29776
rect 10560 29764 10566 29776
rect 10778 29764 10784 29776
rect 10560 29736 10784 29764
rect 10560 29724 10566 29736
rect 10778 29724 10784 29736
rect 10836 29724 10842 29776
rect 11146 29724 11152 29776
rect 11204 29724 11210 29776
rect 12084 29764 12112 29804
rect 12544 29804 13952 29832
rect 12544 29764 12572 29804
rect 12084 29736 12572 29764
rect 13924 29708 13952 29804
rect 14642 29792 14648 29844
rect 14700 29832 14706 29844
rect 17405 29835 17463 29841
rect 14700 29804 15884 29832
rect 14700 29792 14706 29804
rect 10134 29696 10140 29708
rect 6196 29668 7512 29696
rect 7852 29668 10140 29696
rect 4065 29631 4123 29637
rect 4065 29597 4077 29631
rect 4111 29628 4123 29631
rect 6196 29628 6224 29668
rect 4111 29600 6224 29628
rect 4111 29597 4123 29600
rect 4065 29591 4123 29597
rect 6914 29588 6920 29640
rect 6972 29588 6978 29640
rect 7101 29631 7159 29637
rect 7101 29597 7113 29631
rect 7147 29628 7159 29631
rect 7282 29628 7288 29640
rect 7147 29600 7288 29628
rect 7147 29597 7159 29600
rect 7101 29591 7159 29597
rect 7282 29588 7288 29600
rect 7340 29588 7346 29640
rect 7852 29637 7880 29668
rect 10134 29656 10140 29668
rect 10192 29656 10198 29708
rect 10318 29696 10324 29708
rect 10244 29668 10324 29696
rect 7837 29631 7895 29637
rect 7837 29597 7849 29631
rect 7883 29597 7895 29631
rect 7837 29591 7895 29597
rect 7926 29588 7932 29640
rect 7984 29637 7990 29640
rect 7984 29631 8012 29637
rect 8000 29597 8012 29631
rect 7984 29591 8012 29597
rect 7984 29588 7990 29591
rect 8110 29588 8116 29640
rect 8168 29588 8174 29640
rect 9674 29588 9680 29640
rect 9732 29628 9738 29640
rect 10244 29628 10272 29668
rect 10318 29656 10324 29668
rect 10376 29696 10382 29708
rect 11606 29705 11612 29708
rect 11425 29699 11483 29705
rect 11425 29696 11437 29699
rect 10376 29668 11437 29696
rect 10376 29656 10382 29668
rect 11425 29665 11437 29668
rect 11471 29665 11483 29699
rect 11425 29659 11483 29665
rect 11563 29699 11612 29705
rect 11563 29665 11575 29699
rect 11609 29665 11612 29699
rect 11563 29659 11612 29665
rect 11606 29656 11612 29659
rect 11664 29656 11670 29708
rect 11701 29699 11759 29705
rect 11701 29665 11713 29699
rect 11747 29696 11759 29699
rect 12066 29696 12072 29708
rect 11747 29668 12072 29696
rect 11747 29665 11759 29668
rect 11701 29659 11759 29665
rect 12066 29656 12072 29668
rect 12124 29656 12130 29708
rect 12342 29656 12348 29708
rect 12400 29656 12406 29708
rect 13906 29656 13912 29708
rect 13964 29696 13970 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 13964 29668 14197 29696
rect 13964 29656 13970 29668
rect 14185 29665 14197 29668
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 15746 29656 15752 29708
rect 15804 29656 15810 29708
rect 15856 29696 15884 29804
rect 17405 29801 17417 29835
rect 17451 29832 17463 29835
rect 17494 29832 17500 29844
rect 17451 29804 17500 29832
rect 17451 29801 17463 29804
rect 17405 29795 17463 29801
rect 17494 29792 17500 29804
rect 17552 29792 17558 29844
rect 20530 29792 20536 29844
rect 20588 29792 20594 29844
rect 22830 29832 22836 29844
rect 22204 29804 22836 29832
rect 16206 29724 16212 29776
rect 16264 29724 16270 29776
rect 17770 29724 17776 29776
rect 17828 29764 17834 29776
rect 19886 29764 19892 29776
rect 17828 29736 19892 29764
rect 17828 29724 17834 29736
rect 19886 29724 19892 29736
rect 19944 29724 19950 29776
rect 16485 29699 16543 29705
rect 16485 29696 16497 29699
rect 15856 29668 16497 29696
rect 16485 29665 16497 29668
rect 16531 29665 16543 29699
rect 16485 29659 16543 29665
rect 16761 29699 16819 29705
rect 16761 29665 16773 29699
rect 16807 29696 16819 29699
rect 16942 29696 16948 29708
rect 16807 29668 16948 29696
rect 16807 29665 16819 29668
rect 16761 29659 16819 29665
rect 16942 29656 16948 29668
rect 17000 29656 17006 29708
rect 17126 29656 17132 29708
rect 17184 29696 17190 29708
rect 17184 29668 17816 29696
rect 17184 29656 17190 29668
rect 17788 29640 17816 29668
rect 9732 29600 10272 29628
rect 9732 29588 9738 29600
rect 10410 29588 10416 29640
rect 10468 29588 10474 29640
rect 10505 29631 10563 29637
rect 10505 29597 10517 29631
rect 10551 29628 10563 29631
rect 10594 29628 10600 29640
rect 10551 29600 10600 29628
rect 10551 29597 10563 29600
rect 10505 29591 10563 29597
rect 10594 29588 10600 29600
rect 10652 29588 10658 29640
rect 10689 29631 10747 29637
rect 10689 29597 10701 29631
rect 10735 29597 10747 29631
rect 10689 29591 10747 29597
rect 12437 29631 12495 29637
rect 12437 29597 12449 29631
rect 12483 29597 12495 29631
rect 12710 29627 12716 29640
rect 12437 29591 12495 29597
rect 12679 29621 12716 29627
rect 1360 29532 2774 29560
rect 1360 29520 1366 29532
rect 3326 29520 3332 29572
rect 3384 29560 3390 29572
rect 3384 29532 5120 29560
rect 3384 29520 3390 29532
rect 4982 29452 4988 29504
rect 5040 29452 5046 29504
rect 5092 29492 5120 29532
rect 5258 29520 5264 29572
rect 5316 29520 5322 29572
rect 5350 29520 5356 29572
rect 5408 29520 5414 29572
rect 5718 29520 5724 29572
rect 5776 29520 5782 29572
rect 10428 29560 10456 29588
rect 10704 29560 10732 29591
rect 5828 29532 6224 29560
rect 5828 29492 5856 29532
rect 5092 29464 5856 29492
rect 6086 29452 6092 29504
rect 6144 29452 6150 29504
rect 6196 29492 6224 29532
rect 9646 29532 10732 29560
rect 9646 29492 9674 29532
rect 6196 29464 9674 29492
rect 11974 29452 11980 29504
rect 12032 29492 12038 29504
rect 12452 29492 12480 29591
rect 12679 29587 12691 29621
rect 12768 29588 12774 29640
rect 14459 29631 14517 29637
rect 14459 29597 14471 29631
rect 14505 29628 14517 29631
rect 14550 29628 14556 29640
rect 14505 29600 14556 29628
rect 14505 29597 14517 29600
rect 14459 29591 14517 29597
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 15565 29631 15623 29637
rect 15565 29597 15577 29631
rect 15611 29628 15623 29631
rect 15930 29628 15936 29640
rect 15611 29600 15936 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 15930 29588 15936 29600
rect 15988 29588 15994 29640
rect 16574 29588 16580 29640
rect 16632 29637 16638 29640
rect 16632 29631 16660 29637
rect 16648 29597 16660 29631
rect 16632 29591 16660 29597
rect 16632 29588 16638 29591
rect 17770 29588 17776 29640
rect 17828 29588 17834 29640
rect 20548 29628 20576 29792
rect 21729 29699 21787 29705
rect 21729 29665 21741 29699
rect 21775 29696 21787 29699
rect 22097 29699 22155 29705
rect 22097 29696 22109 29699
rect 21775 29668 22109 29696
rect 21775 29665 21787 29668
rect 21729 29659 21787 29665
rect 22097 29665 22109 29668
rect 22143 29665 22155 29699
rect 22097 29659 22155 29665
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 20548 29600 21189 29628
rect 21177 29597 21189 29600
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 21637 29631 21695 29637
rect 21637 29597 21649 29631
rect 21683 29597 21695 29631
rect 21637 29591 21695 29597
rect 22005 29631 22063 29637
rect 22005 29597 22017 29631
rect 22051 29628 22063 29631
rect 22204 29628 22232 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 23198 29792 23204 29844
rect 23256 29832 23262 29844
rect 23256 29804 23704 29832
rect 23256 29792 23262 29804
rect 23293 29767 23351 29773
rect 23293 29733 23305 29767
rect 23339 29733 23351 29767
rect 23293 29727 23351 29733
rect 23569 29767 23627 29773
rect 23569 29733 23581 29767
rect 23615 29733 23627 29767
rect 23569 29727 23627 29733
rect 22281 29699 22339 29705
rect 22281 29665 22293 29699
rect 22327 29696 22339 29699
rect 22465 29699 22523 29705
rect 22465 29696 22477 29699
rect 22327 29668 22477 29696
rect 22327 29665 22339 29668
rect 22281 29659 22339 29665
rect 22465 29665 22477 29668
rect 22511 29665 22523 29699
rect 22465 29659 22523 29665
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22051 29600 22385 29628
rect 22051 29597 22063 29600
rect 22005 29591 22063 29597
rect 22373 29597 22385 29600
rect 22419 29597 22431 29631
rect 22373 29591 22431 29597
rect 12725 29587 12737 29588
rect 12679 29581 12737 29587
rect 21652 29560 21680 29591
rect 22554 29588 22560 29640
rect 22612 29588 22618 29640
rect 21008 29532 21680 29560
rect 22281 29563 22339 29569
rect 12032 29464 12480 29492
rect 12032 29452 12038 29464
rect 13446 29452 13452 29504
rect 13504 29452 13510 29504
rect 14458 29452 14464 29504
rect 14516 29492 14522 29504
rect 15197 29495 15255 29501
rect 15197 29492 15209 29495
rect 14516 29464 15209 29492
rect 14516 29452 14522 29464
rect 15197 29461 15209 29464
rect 15243 29461 15255 29495
rect 15197 29455 15255 29461
rect 15930 29452 15936 29504
rect 15988 29492 15994 29504
rect 16666 29492 16672 29504
rect 15988 29464 16672 29492
rect 15988 29452 15994 29464
rect 16666 29452 16672 29464
rect 16724 29492 16730 29504
rect 17034 29492 17040 29504
rect 16724 29464 17040 29492
rect 16724 29452 16730 29464
rect 17034 29452 17040 29464
rect 17092 29452 17098 29504
rect 17862 29452 17868 29504
rect 17920 29492 17926 29504
rect 19978 29492 19984 29504
rect 17920 29464 19984 29492
rect 17920 29452 17926 29464
rect 19978 29452 19984 29464
rect 20036 29452 20042 29504
rect 21008 29501 21036 29532
rect 22281 29529 22293 29563
rect 22327 29529 22339 29563
rect 23308 29560 23336 29727
rect 23485 29631 23543 29637
rect 23485 29597 23497 29631
rect 23531 29628 23543 29631
rect 23584 29628 23612 29727
rect 23531 29600 23612 29628
rect 23676 29628 23704 29804
rect 23753 29631 23811 29637
rect 23753 29628 23765 29631
rect 23676 29600 23765 29628
rect 23531 29597 23543 29600
rect 23485 29591 23543 29597
rect 23753 29597 23765 29600
rect 23799 29597 23811 29631
rect 23753 29591 23811 29597
rect 23937 29631 23995 29637
rect 23937 29597 23949 29631
rect 23983 29597 23995 29631
rect 23937 29591 23995 29597
rect 23952 29560 23980 29591
rect 24302 29560 24308 29572
rect 23308 29532 23980 29560
rect 24044 29532 24308 29560
rect 22281 29523 22339 29529
rect 20993 29495 21051 29501
rect 20993 29461 21005 29495
rect 21039 29461 21051 29495
rect 22296 29492 22324 29523
rect 24044 29492 24072 29532
rect 24302 29520 24308 29532
rect 24360 29520 24366 29572
rect 22296 29464 24072 29492
rect 24121 29495 24179 29501
rect 20993 29455 21051 29461
rect 24121 29461 24133 29495
rect 24167 29492 24179 29495
rect 25130 29492 25136 29504
rect 24167 29464 25136 29492
rect 24167 29461 24179 29464
rect 24121 29455 24179 29461
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 1104 29402 25000 29424
rect 1104 29350 6884 29402
rect 6936 29350 6948 29402
rect 7000 29350 7012 29402
rect 7064 29350 7076 29402
rect 7128 29350 7140 29402
rect 7192 29350 12818 29402
rect 12870 29350 12882 29402
rect 12934 29350 12946 29402
rect 12998 29350 13010 29402
rect 13062 29350 13074 29402
rect 13126 29350 18752 29402
rect 18804 29350 18816 29402
rect 18868 29350 18880 29402
rect 18932 29350 18944 29402
rect 18996 29350 19008 29402
rect 19060 29350 24686 29402
rect 24738 29350 24750 29402
rect 24802 29350 24814 29402
rect 24866 29350 24878 29402
rect 24930 29350 24942 29402
rect 24994 29350 25000 29402
rect 1104 29328 25000 29350
rect 1578 29248 1584 29300
rect 1636 29288 1642 29300
rect 3789 29291 3847 29297
rect 1636 29260 3464 29288
rect 1636 29248 1642 29260
rect 934 29180 940 29232
rect 992 29220 998 29232
rect 1857 29223 1915 29229
rect 1857 29220 1869 29223
rect 992 29192 1869 29220
rect 992 29180 998 29192
rect 1857 29189 1869 29192
rect 1903 29189 1915 29223
rect 3326 29220 3332 29232
rect 1857 29183 1915 29189
rect 1962 29192 3332 29220
rect 1486 29112 1492 29164
rect 1544 29112 1550 29164
rect 1962 29084 1990 29192
rect 3326 29180 3332 29192
rect 3384 29180 3390 29232
rect 2498 29152 2504 29164
rect 2459 29124 2504 29152
rect 2498 29112 2504 29124
rect 2556 29112 2562 29164
rect 1780 29056 1990 29084
rect 1302 28908 1308 28960
rect 1360 28948 1366 28960
rect 1780 28948 1808 29056
rect 2222 29044 2228 29096
rect 2280 29044 2286 29096
rect 1946 28976 1952 29028
rect 2004 28976 2010 29028
rect 2038 28976 2044 29028
rect 2096 28976 2102 29028
rect 3436 29016 3464 29260
rect 3789 29257 3801 29291
rect 3835 29257 3847 29291
rect 3789 29251 3847 29257
rect 3804 29220 3832 29251
rect 5350 29248 5356 29300
rect 5408 29288 5414 29300
rect 5905 29291 5963 29297
rect 5905 29288 5917 29291
rect 5408 29260 5917 29288
rect 5408 29248 5414 29260
rect 5905 29257 5917 29260
rect 5951 29257 5963 29291
rect 5905 29251 5963 29257
rect 6086 29248 6092 29300
rect 6144 29288 6150 29300
rect 6144 29260 8064 29288
rect 6144 29248 6150 29260
rect 7926 29220 7932 29232
rect 3804 29192 7932 29220
rect 7926 29180 7932 29192
rect 7984 29180 7990 29232
rect 3602 29112 3608 29164
rect 3660 29112 3666 29164
rect 4246 29112 4252 29164
rect 4304 29152 4310 29164
rect 4893 29155 4951 29161
rect 4893 29152 4905 29155
rect 4304 29124 4905 29152
rect 4304 29112 4310 29124
rect 4893 29121 4905 29124
rect 4939 29121 4951 29155
rect 4893 29115 4951 29121
rect 5074 29112 5080 29164
rect 5132 29152 5138 29164
rect 5167 29155 5225 29161
rect 5167 29152 5179 29155
rect 5132 29124 5179 29152
rect 5132 29112 5138 29124
rect 5167 29121 5179 29124
rect 5213 29121 5225 29155
rect 5167 29115 5225 29121
rect 7558 29112 7564 29164
rect 7616 29152 7622 29164
rect 7651 29155 7709 29161
rect 7651 29152 7663 29155
rect 7616 29124 7663 29152
rect 7616 29112 7622 29124
rect 7651 29121 7663 29124
rect 7697 29121 7709 29155
rect 8036 29156 8064 29260
rect 8110 29248 8116 29300
rect 8168 29288 8174 29300
rect 8389 29291 8447 29297
rect 8389 29288 8401 29291
rect 8168 29260 8401 29288
rect 8168 29248 8174 29260
rect 8389 29257 8401 29260
rect 8435 29257 8447 29291
rect 8389 29251 8447 29257
rect 10870 29248 10876 29300
rect 10928 29248 10934 29300
rect 11330 29288 11336 29300
rect 10980 29260 11336 29288
rect 8754 29180 8760 29232
rect 8812 29220 8818 29232
rect 10980 29220 11008 29260
rect 11330 29248 11336 29260
rect 11388 29248 11394 29300
rect 13998 29248 14004 29300
rect 14056 29288 14062 29300
rect 14277 29291 14335 29297
rect 14277 29288 14289 29291
rect 14056 29260 14289 29288
rect 14056 29248 14062 29260
rect 14277 29257 14289 29260
rect 14323 29257 14335 29291
rect 14277 29251 14335 29257
rect 14458 29248 14464 29300
rect 14516 29288 14522 29300
rect 14516 29260 14688 29288
rect 14516 29248 14522 29260
rect 8812 29192 11008 29220
rect 8812 29180 8818 29192
rect 11054 29180 11060 29232
rect 11112 29220 11118 29232
rect 11609 29223 11667 29229
rect 11609 29220 11621 29223
rect 11112 29192 11621 29220
rect 11112 29180 11118 29192
rect 11609 29189 11621 29192
rect 11655 29220 11667 29223
rect 11790 29220 11796 29232
rect 11655 29192 11796 29220
rect 11655 29189 11667 29192
rect 11609 29183 11667 29189
rect 11790 29180 11796 29192
rect 11848 29180 11854 29232
rect 12158 29180 12164 29232
rect 12216 29220 12222 29232
rect 12216 29192 12756 29220
rect 12216 29180 12222 29192
rect 8036 29128 8322 29156
rect 7651 29115 7709 29121
rect 6454 29044 6460 29096
rect 6512 29084 6518 29096
rect 7282 29084 7288 29096
rect 6512 29056 7288 29084
rect 6512 29044 6518 29056
rect 7282 29044 7288 29056
rect 7340 29084 7346 29096
rect 7377 29087 7435 29093
rect 7377 29084 7389 29087
rect 7340 29056 7389 29084
rect 7340 29044 7346 29056
rect 7377 29053 7389 29056
rect 7423 29053 7435 29087
rect 7377 29047 7435 29053
rect 8110 29016 8116 29028
rect 3436 28988 5028 29016
rect 1360 28920 1808 28948
rect 1964 28948 1992 28976
rect 2590 28948 2596 28960
rect 1964 28920 2596 28948
rect 1360 28908 1366 28920
rect 2590 28908 2596 28920
rect 2648 28908 2654 28960
rect 3234 28908 3240 28960
rect 3292 28908 3298 28960
rect 5000 28948 5028 28988
rect 5552 28988 7512 29016
rect 5552 28948 5580 28988
rect 5000 28920 5580 28948
rect 7484 28948 7512 28988
rect 8036 28988 8116 29016
rect 8036 28948 8064 28988
rect 8110 28976 8116 28988
rect 8168 28976 8174 29028
rect 8294 29016 8322 29128
rect 9030 29112 9036 29164
rect 9088 29152 9094 29164
rect 9217 29155 9275 29161
rect 9217 29152 9229 29155
rect 9088 29124 9229 29152
rect 9088 29112 9094 29124
rect 9217 29121 9229 29124
rect 9263 29121 9275 29155
rect 9490 29152 9496 29164
rect 9451 29124 9496 29152
rect 9217 29115 9275 29121
rect 9490 29112 9496 29124
rect 9548 29112 9554 29164
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29152 10655 29155
rect 11330 29152 11336 29164
rect 10643 29124 11336 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 10229 29019 10287 29025
rect 8294 28994 8340 29016
rect 8404 28994 9352 29016
rect 8294 28988 9352 28994
rect 8312 28966 8432 28988
rect 7484 28920 8064 28948
rect 9324 28948 9352 28988
rect 10229 28985 10241 29019
rect 10275 29016 10287 29019
rect 10612 29016 10640 29115
rect 11330 29112 11336 29124
rect 11388 29112 11394 29164
rect 12434 29112 12440 29164
rect 12492 29152 12498 29164
rect 12529 29155 12587 29161
rect 12529 29152 12541 29155
rect 12492 29124 12541 29152
rect 12492 29112 12498 29124
rect 12529 29121 12541 29124
rect 12575 29121 12587 29155
rect 12728 29150 12756 29192
rect 13814 29180 13820 29232
rect 13872 29220 13878 29232
rect 14550 29220 14556 29232
rect 13872 29192 14556 29220
rect 13872 29180 13878 29192
rect 14550 29180 14556 29192
rect 14608 29180 14614 29232
rect 14660 29229 14688 29260
rect 14826 29248 14832 29300
rect 14884 29288 14890 29300
rect 23109 29291 23167 29297
rect 14884 29260 15056 29288
rect 14884 29248 14890 29260
rect 15028 29229 15056 29260
rect 15304 29260 22094 29288
rect 14645 29223 14703 29229
rect 14645 29189 14657 29223
rect 14691 29189 14703 29223
rect 14645 29183 14703 29189
rect 15013 29223 15071 29229
rect 15013 29189 15025 29223
rect 15059 29189 15071 29223
rect 15013 29183 15071 29189
rect 12803 29155 12861 29161
rect 12803 29150 12815 29155
rect 12728 29122 12815 29150
rect 12529 29115 12587 29121
rect 12803 29121 12815 29122
rect 12849 29150 12861 29155
rect 15304 29152 15332 29260
rect 15381 29223 15439 29229
rect 15381 29189 15393 29223
rect 15427 29189 15439 29223
rect 15381 29183 15439 29189
rect 16786 29192 19555 29220
rect 12912 29150 15332 29152
rect 12849 29124 15332 29150
rect 15396 29152 15424 29183
rect 15470 29152 15476 29164
rect 15396 29124 15476 29152
rect 12849 29122 12940 29124
rect 12849 29121 12861 29122
rect 12803 29115 12861 29121
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 16786 29152 16814 29192
rect 15580 29124 16814 29152
rect 10873 29087 10931 29093
rect 10873 29053 10885 29087
rect 10919 29084 10931 29087
rect 10919 29056 11468 29084
rect 10919 29053 10931 29056
rect 10873 29047 10931 29053
rect 10275 28988 10640 29016
rect 10689 29019 10747 29025
rect 10275 28985 10287 28988
rect 10229 28979 10287 28985
rect 10689 28985 10701 29019
rect 10735 29016 10747 29019
rect 11146 29016 11152 29028
rect 10735 28988 11152 29016
rect 10735 28985 10747 28988
rect 10689 28979 10747 28985
rect 11146 28976 11152 28988
rect 11204 28976 11210 29028
rect 11440 28960 11468 29056
rect 11974 29044 11980 29096
rect 12032 29084 12038 29096
rect 12032 29056 12572 29084
rect 12032 29044 12038 29056
rect 11790 28976 11796 29028
rect 11848 28976 11854 29028
rect 11882 28976 11888 29028
rect 11940 29016 11946 29028
rect 12434 29016 12440 29028
rect 11940 28988 12440 29016
rect 11940 28976 11946 28988
rect 12434 28976 12440 28988
rect 12492 28976 12498 29028
rect 12544 29016 12572 29056
rect 14918 29044 14924 29096
rect 14976 29044 14982 29096
rect 15580 29025 15608 29124
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 16943 29155 17001 29161
rect 16943 29152 16955 29155
rect 16908 29124 16955 29152
rect 16908 29112 16914 29124
rect 16943 29121 16955 29124
rect 16989 29121 17001 29155
rect 16943 29115 17001 29121
rect 17862 29112 17868 29164
rect 17920 29112 17926 29164
rect 18598 29112 18604 29164
rect 18656 29152 18662 29164
rect 19151 29155 19209 29161
rect 19151 29152 19163 29155
rect 18656 29124 19163 29152
rect 18656 29112 18662 29124
rect 19151 29121 19163 29124
rect 19197 29121 19209 29155
rect 19151 29115 19209 29121
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 16224 29056 16681 29084
rect 15565 29019 15623 29025
rect 12544 29006 12664 29016
rect 12544 28988 12624 29006
rect 9582 28948 9588 28960
rect 9324 28920 9588 28948
rect 9582 28908 9588 28920
rect 9640 28908 9646 28960
rect 11422 28908 11428 28960
rect 11480 28908 11486 28960
rect 12618 28954 12624 28988
rect 12676 28954 12682 29006
rect 15565 28985 15577 29019
rect 15611 28985 15623 29019
rect 15565 28979 15623 28985
rect 16224 28960 16252 29056
rect 16669 29053 16681 29056
rect 16715 29053 16727 29087
rect 17880 29084 17908 29112
rect 18877 29087 18935 29093
rect 18877 29084 18889 29087
rect 17880 29056 18889 29084
rect 16669 29047 16727 29053
rect 18877 29053 18889 29056
rect 18923 29053 18935 29087
rect 18877 29047 18935 29053
rect 17954 28976 17960 29028
rect 18012 29016 18018 29028
rect 18598 29016 18604 29028
rect 18012 28988 18604 29016
rect 18012 28976 18018 28988
rect 18598 28976 18604 28988
rect 18656 28976 18662 29028
rect 19527 29016 19555 29192
rect 20257 29155 20315 29161
rect 20257 29152 20269 29155
rect 19628 29124 20269 29152
rect 19628 29096 19656 29124
rect 20257 29121 20269 29124
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29121 20499 29155
rect 22066 29152 22094 29260
rect 23109 29257 23121 29291
rect 23155 29257 23167 29291
rect 23109 29251 23167 29257
rect 23124 29220 23152 29251
rect 23124 29192 23888 29220
rect 23860 29161 23888 29192
rect 23293 29155 23351 29161
rect 23293 29152 23305 29155
rect 22066 29124 23305 29152
rect 20441 29115 20499 29121
rect 23293 29121 23305 29124
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 23569 29155 23627 29161
rect 23569 29121 23581 29155
rect 23615 29121 23627 29155
rect 23569 29115 23627 29121
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29121 23903 29155
rect 23845 29115 23903 29121
rect 24121 29155 24179 29161
rect 24121 29121 24133 29155
rect 24167 29121 24179 29155
rect 24121 29115 24179 29121
rect 19610 29044 19616 29096
rect 19668 29044 19674 29096
rect 19702 29044 19708 29096
rect 19760 29084 19766 29096
rect 20456 29084 20484 29115
rect 19760 29056 20484 29084
rect 19760 29044 19766 29056
rect 23106 29016 23112 29028
rect 19527 28988 23112 29016
rect 23106 28976 23112 28988
rect 23164 28976 23170 29028
rect 23385 29019 23443 29025
rect 23385 28985 23397 29019
rect 23431 29016 23443 29019
rect 23584 29016 23612 29115
rect 24136 29084 24164 29115
rect 23768 29056 24164 29084
rect 23661 29019 23719 29025
rect 23661 29016 23673 29019
rect 23431 28988 23520 29016
rect 23584 28988 23673 29016
rect 23431 28985 23443 28988
rect 23385 28979 23443 28985
rect 13541 28951 13599 28957
rect 13541 28917 13553 28951
rect 13587 28948 13599 28951
rect 13722 28948 13728 28960
rect 13587 28920 13728 28948
rect 13587 28917 13599 28920
rect 13541 28911 13599 28917
rect 13722 28908 13728 28920
rect 13780 28908 13786 28960
rect 13814 28908 13820 28960
rect 13872 28948 13878 28960
rect 14274 28948 14280 28960
rect 13872 28920 14280 28948
rect 13872 28908 13878 28920
rect 14274 28908 14280 28920
rect 14332 28908 14338 28960
rect 16206 28908 16212 28960
rect 16264 28908 16270 28960
rect 17402 28908 17408 28960
rect 17460 28948 17466 28960
rect 17681 28951 17739 28957
rect 17681 28948 17693 28951
rect 17460 28920 17693 28948
rect 17460 28908 17466 28920
rect 17681 28917 17693 28920
rect 17727 28917 17739 28951
rect 17681 28911 17739 28917
rect 19610 28908 19616 28960
rect 19668 28948 19674 28960
rect 19889 28951 19947 28957
rect 19889 28948 19901 28951
rect 19668 28920 19901 28948
rect 19668 28908 19674 28920
rect 19889 28917 19901 28920
rect 19935 28917 19947 28951
rect 19889 28911 19947 28917
rect 20346 28908 20352 28960
rect 20404 28908 20410 28960
rect 20530 28908 20536 28960
rect 20588 28948 20594 28960
rect 21174 28948 21180 28960
rect 20588 28920 21180 28948
rect 20588 28908 20594 28920
rect 21174 28908 21180 28920
rect 21232 28908 21238 28960
rect 23492 28948 23520 28988
rect 23661 28985 23673 28988
rect 23707 28985 23719 29019
rect 23661 28979 23719 28985
rect 23768 28948 23796 29056
rect 24394 28976 24400 29028
rect 24452 28976 24458 29028
rect 23492 28920 23796 28948
rect 1104 28858 24840 28880
rect 1104 28806 3917 28858
rect 3969 28806 3981 28858
rect 4033 28806 4045 28858
rect 4097 28806 4109 28858
rect 4161 28806 4173 28858
rect 4225 28806 9851 28858
rect 9903 28806 9915 28858
rect 9967 28806 9979 28858
rect 10031 28806 10043 28858
rect 10095 28806 10107 28858
rect 10159 28806 15785 28858
rect 15837 28806 15849 28858
rect 15901 28806 15913 28858
rect 15965 28806 15977 28858
rect 16029 28806 16041 28858
rect 16093 28806 21719 28858
rect 21771 28806 21783 28858
rect 21835 28806 21847 28858
rect 21899 28806 21911 28858
rect 21963 28806 21975 28858
rect 22027 28806 24840 28858
rect 1104 28784 24840 28806
rect 2774 28744 2780 28756
rect 1688 28716 2780 28744
rect 1688 28617 1716 28716
rect 2774 28704 2780 28716
rect 2832 28704 2838 28756
rect 9766 28744 9772 28756
rect 2976 28716 9772 28744
rect 1673 28611 1731 28617
rect 1673 28577 1685 28611
rect 1719 28577 1731 28611
rect 1673 28571 1731 28577
rect 2222 28568 2228 28620
rect 2280 28608 2286 28620
rect 2317 28611 2375 28617
rect 2317 28608 2329 28611
rect 2280 28580 2329 28608
rect 2280 28568 2286 28580
rect 2317 28577 2329 28580
rect 2363 28577 2375 28611
rect 2317 28571 2375 28577
rect 2976 28552 3004 28716
rect 9766 28704 9772 28716
rect 9824 28704 9830 28756
rect 11146 28704 11152 28756
rect 11204 28704 11210 28756
rect 11422 28704 11428 28756
rect 11480 28704 11486 28756
rect 11606 28704 11612 28756
rect 11664 28744 11670 28756
rect 13814 28744 13820 28756
rect 11664 28716 13820 28744
rect 11664 28704 11670 28716
rect 13814 28704 13820 28716
rect 13872 28704 13878 28756
rect 18877 28747 18935 28753
rect 13924 28716 18552 28744
rect 10781 28679 10839 28685
rect 10781 28645 10793 28679
rect 10827 28645 10839 28679
rect 10781 28639 10839 28645
rect 7282 28568 7288 28620
rect 7340 28608 7346 28620
rect 7742 28608 7748 28620
rect 7340 28580 7748 28608
rect 7340 28568 7346 28580
rect 7742 28568 7748 28580
rect 7800 28608 7806 28620
rect 8941 28611 8999 28617
rect 8941 28608 8953 28611
rect 7800 28580 8953 28608
rect 7800 28568 7806 28580
rect 8941 28577 8953 28580
rect 8987 28577 8999 28611
rect 8941 28571 8999 28577
rect 9674 28568 9680 28620
rect 9732 28568 9738 28620
rect 10796 28608 10824 28639
rect 13924 28608 13952 28716
rect 18417 28679 18475 28685
rect 18417 28645 18429 28679
rect 18463 28645 18475 28679
rect 18524 28676 18552 28716
rect 18877 28713 18889 28747
rect 18923 28744 18935 28747
rect 19702 28744 19708 28756
rect 18923 28716 19708 28744
rect 18923 28713 18935 28716
rect 18877 28707 18935 28713
rect 19702 28704 19708 28716
rect 19760 28704 19766 28756
rect 20346 28744 20352 28756
rect 19904 28716 20352 28744
rect 19518 28676 19524 28688
rect 18524 28648 19524 28676
rect 18417 28639 18475 28645
rect 10796 28580 11560 28608
rect 842 28500 848 28552
rect 900 28540 906 28552
rect 1397 28543 1455 28549
rect 1397 28540 1409 28543
rect 900 28512 1409 28540
rect 900 28500 906 28512
rect 1397 28509 1409 28512
rect 1443 28509 1455 28543
rect 2575 28513 2633 28519
rect 2575 28510 2587 28513
rect 1397 28503 1455 28509
rect 2406 28432 2412 28484
rect 2464 28472 2470 28484
rect 2516 28482 2587 28510
rect 2516 28472 2544 28482
rect 2575 28479 2587 28482
rect 2621 28479 2633 28513
rect 2958 28500 2964 28552
rect 3016 28500 3022 28552
rect 3602 28500 3608 28552
rect 3660 28540 3666 28552
rect 3881 28543 3939 28549
rect 3881 28540 3893 28543
rect 3660 28512 3893 28540
rect 3660 28500 3666 28512
rect 3881 28509 3893 28512
rect 3927 28509 3939 28543
rect 3881 28503 3939 28509
rect 4155 28543 4213 28549
rect 4155 28509 4167 28543
rect 4201 28540 4213 28543
rect 4890 28540 4896 28552
rect 4201 28512 4896 28540
rect 4201 28509 4213 28512
rect 4155 28503 4213 28509
rect 2575 28473 2633 28479
rect 2464 28444 2544 28472
rect 2464 28432 2470 28444
rect 3326 28364 3332 28416
rect 3384 28364 3390 28416
rect 3510 28364 3516 28416
rect 3568 28404 3574 28416
rect 4170 28404 4198 28503
rect 4890 28500 4896 28512
rect 4948 28500 4954 28552
rect 5074 28500 5080 28552
rect 5132 28540 5138 28552
rect 8110 28540 8116 28552
rect 5132 28512 8116 28540
rect 5132 28500 5138 28512
rect 8110 28500 8116 28512
rect 8168 28500 8174 28552
rect 8846 28500 8852 28552
rect 8904 28540 8910 28552
rect 8904 28519 9242 28540
rect 8904 28513 9257 28519
rect 8904 28512 9211 28513
rect 8904 28500 8910 28512
rect 5350 28472 5356 28484
rect 4356 28444 5356 28472
rect 4356 28416 4384 28444
rect 5350 28432 5356 28444
rect 5408 28432 5414 28484
rect 9199 28479 9211 28512
rect 9245 28510 9257 28513
rect 9245 28479 9258 28510
rect 9199 28473 9258 28479
rect 9230 28472 9258 28473
rect 9230 28444 9536 28472
rect 9508 28416 9536 28444
rect 9692 28416 9720 28568
rect 10686 28500 10692 28552
rect 10744 28500 10750 28552
rect 10962 28500 10968 28552
rect 11020 28500 11026 28552
rect 11057 28543 11115 28549
rect 11057 28509 11069 28543
rect 11103 28509 11115 28543
rect 11057 28503 11115 28509
rect 11072 28472 11100 28503
rect 11330 28500 11336 28552
rect 11388 28500 11394 28552
rect 11532 28549 11560 28580
rect 12360 28580 13952 28608
rect 11517 28543 11575 28549
rect 11517 28509 11529 28543
rect 11563 28509 11575 28543
rect 11517 28503 11575 28509
rect 11606 28500 11612 28552
rect 11664 28540 11670 28552
rect 11701 28543 11759 28549
rect 11701 28540 11713 28543
rect 11664 28512 11713 28540
rect 11664 28500 11670 28512
rect 11701 28509 11713 28512
rect 11747 28509 11759 28543
rect 11975 28543 12033 28549
rect 11975 28540 11987 28543
rect 11701 28503 11759 28509
rect 11790 28512 11987 28540
rect 10520 28444 11100 28472
rect 3568 28376 4198 28404
rect 3568 28364 3574 28376
rect 4338 28364 4344 28416
rect 4396 28364 4402 28416
rect 4890 28364 4896 28416
rect 4948 28364 4954 28416
rect 5718 28364 5724 28416
rect 5776 28404 5782 28416
rect 7466 28404 7472 28416
rect 5776 28376 7472 28404
rect 5776 28364 5782 28376
rect 7466 28364 7472 28376
rect 7524 28364 7530 28416
rect 9490 28364 9496 28416
rect 9548 28364 9554 28416
rect 9674 28364 9680 28416
rect 9732 28364 9738 28416
rect 9953 28407 10011 28413
rect 9953 28373 9965 28407
rect 9999 28404 10011 28407
rect 10318 28404 10324 28416
rect 9999 28376 10324 28404
rect 9999 28373 10011 28376
rect 9953 28367 10011 28373
rect 10318 28364 10324 28376
rect 10376 28364 10382 28416
rect 10520 28413 10548 28444
rect 10505 28407 10563 28413
rect 10505 28373 10517 28407
rect 10551 28373 10563 28407
rect 10505 28367 10563 28373
rect 10870 28364 10876 28416
rect 10928 28404 10934 28416
rect 11790 28404 11818 28512
rect 11975 28509 11987 28512
rect 12021 28540 12033 28543
rect 12360 28540 12388 28580
rect 16666 28568 16672 28620
rect 16724 28568 16730 28620
rect 17221 28611 17279 28617
rect 17221 28577 17233 28611
rect 17267 28608 17279 28611
rect 17402 28608 17408 28620
rect 17267 28580 17408 28608
rect 17267 28577 17279 28580
rect 17221 28571 17279 28577
rect 17402 28568 17408 28580
rect 17460 28568 17466 28620
rect 18432 28608 18460 28639
rect 19518 28636 19524 28648
rect 19576 28636 19582 28688
rect 19904 28617 19932 28716
rect 20346 28704 20352 28716
rect 20404 28704 20410 28756
rect 22649 28747 22707 28753
rect 22649 28713 22661 28747
rect 22695 28744 22707 28747
rect 22695 28716 23152 28744
rect 22695 28713 22707 28716
rect 22649 28707 22707 28713
rect 20714 28636 20720 28688
rect 20772 28676 20778 28688
rect 22922 28676 22928 28688
rect 20772 28648 22928 28676
rect 20772 28636 20778 28648
rect 22922 28636 22928 28648
rect 22980 28636 22986 28688
rect 19337 28611 19395 28617
rect 18432 28580 19288 28608
rect 12021 28512 12388 28540
rect 12450 28512 13216 28540
rect 12021 28509 12033 28512
rect 11975 28503 12033 28509
rect 12066 28432 12072 28484
rect 12124 28472 12130 28484
rect 12450 28472 12478 28512
rect 12124 28444 12478 28472
rect 13188 28472 13216 28512
rect 13906 28500 13912 28552
rect 13964 28540 13970 28552
rect 14093 28543 14151 28549
rect 14093 28540 14105 28543
rect 13964 28512 14105 28540
rect 13964 28500 13970 28512
rect 14093 28509 14105 28512
rect 14139 28509 14151 28543
rect 14093 28503 14151 28509
rect 14367 28543 14425 28549
rect 14367 28509 14379 28543
rect 14413 28540 14425 28543
rect 15102 28540 15108 28552
rect 14413 28512 15108 28540
rect 14413 28509 14425 28512
rect 14367 28503 14425 28509
rect 15102 28500 15108 28512
rect 15160 28500 15166 28552
rect 15194 28500 15200 28552
rect 15252 28540 15258 28552
rect 15562 28540 15568 28552
rect 15252 28512 15568 28540
rect 15252 28500 15258 28512
rect 15562 28500 15568 28512
rect 15620 28540 15626 28552
rect 16025 28543 16083 28549
rect 16025 28540 16037 28543
rect 15620 28512 16037 28540
rect 15620 28500 15626 28512
rect 16025 28509 16037 28512
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 16114 28500 16120 28552
rect 16172 28540 16178 28552
rect 16209 28543 16267 28549
rect 16209 28540 16221 28543
rect 16172 28512 16221 28540
rect 16172 28500 16178 28512
rect 16209 28509 16221 28512
rect 16255 28509 16267 28543
rect 16209 28503 16267 28509
rect 16942 28500 16948 28552
rect 17000 28500 17006 28552
rect 17126 28549 17132 28552
rect 17083 28543 17132 28549
rect 17083 28509 17095 28543
rect 17129 28509 17132 28543
rect 17083 28503 17132 28509
rect 17126 28500 17132 28503
rect 17184 28500 17190 28552
rect 17865 28543 17923 28549
rect 17865 28509 17877 28543
rect 17911 28540 17923 28543
rect 17954 28540 17960 28552
rect 17911 28512 17960 28540
rect 17911 28509 17923 28512
rect 17865 28503 17923 28509
rect 17954 28500 17960 28512
rect 18012 28540 18018 28552
rect 18601 28543 18659 28549
rect 18601 28540 18613 28543
rect 18012 28512 18613 28540
rect 18012 28500 18018 28512
rect 18601 28509 18613 28512
rect 18647 28509 18659 28543
rect 18601 28503 18659 28509
rect 19061 28543 19119 28549
rect 19061 28509 19073 28543
rect 19107 28540 19119 28543
rect 19150 28540 19156 28552
rect 19107 28512 19156 28540
rect 19107 28509 19119 28512
rect 19061 28503 19119 28509
rect 19150 28500 19156 28512
rect 19208 28500 19214 28552
rect 19260 28549 19288 28580
rect 19337 28577 19349 28611
rect 19383 28608 19395 28611
rect 19705 28611 19763 28617
rect 19705 28608 19717 28611
rect 19383 28580 19717 28608
rect 19383 28577 19395 28580
rect 19337 28571 19395 28577
rect 19705 28577 19717 28580
rect 19751 28577 19763 28611
rect 19705 28571 19763 28577
rect 19889 28611 19947 28617
rect 19889 28577 19901 28611
rect 19935 28577 19947 28611
rect 19889 28571 19947 28577
rect 19978 28568 19984 28620
rect 20036 28568 20042 28620
rect 22738 28568 22744 28620
rect 22796 28608 22802 28620
rect 23124 28608 23152 28716
rect 23216 28716 23980 28744
rect 23216 28685 23244 28716
rect 23201 28679 23259 28685
rect 23201 28645 23213 28679
rect 23247 28645 23259 28679
rect 23201 28639 23259 28645
rect 22796 28580 22968 28608
rect 23124 28580 23704 28608
rect 22796 28568 22802 28580
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 19610 28500 19616 28552
rect 19668 28500 19674 28552
rect 20255 28543 20313 28549
rect 20255 28509 20267 28543
rect 20301 28540 20313 28543
rect 20346 28540 20352 28552
rect 20301 28512 20352 28540
rect 20301 28509 20313 28512
rect 20255 28503 20313 28509
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 22833 28543 22891 28549
rect 22833 28540 22845 28543
rect 20916 28512 22845 28540
rect 19889 28475 19947 28481
rect 13188 28444 15238 28472
rect 12124 28432 12130 28444
rect 10928 28376 11818 28404
rect 10928 28364 10934 28376
rect 11882 28364 11888 28416
rect 11940 28404 11946 28416
rect 12713 28407 12771 28413
rect 12713 28404 12725 28407
rect 11940 28376 12725 28404
rect 11940 28364 11946 28376
rect 12713 28373 12725 28376
rect 12759 28373 12771 28407
rect 12713 28367 12771 28373
rect 13078 28364 13084 28416
rect 13136 28404 13142 28416
rect 13262 28404 13268 28416
rect 13136 28376 13268 28404
rect 13136 28364 13142 28376
rect 13262 28364 13268 28376
rect 13320 28364 13326 28416
rect 13998 28364 14004 28416
rect 14056 28404 14062 28416
rect 14274 28404 14280 28416
rect 14056 28376 14280 28404
rect 14056 28364 14062 28376
rect 14274 28364 14280 28376
rect 14332 28404 14338 28416
rect 15105 28407 15163 28413
rect 15105 28404 15117 28407
rect 14332 28376 15117 28404
rect 14332 28364 14338 28376
rect 15105 28373 15117 28376
rect 15151 28373 15163 28407
rect 15210 28404 15238 28444
rect 19889 28441 19901 28475
rect 19935 28472 19947 28475
rect 20438 28472 20444 28484
rect 19935 28444 20444 28472
rect 19935 28441 19947 28444
rect 19889 28435 19947 28441
rect 20438 28432 20444 28444
rect 20496 28432 20502 28484
rect 20916 28404 20944 28512
rect 22833 28509 22845 28512
rect 22879 28509 22891 28543
rect 22940 28540 22968 28580
rect 23290 28540 23296 28552
rect 22940 28512 23296 28540
rect 22833 28503 22891 28509
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 23676 28549 23704 28580
rect 23952 28549 23980 28716
rect 23385 28543 23443 28549
rect 23385 28509 23397 28543
rect 23431 28540 23443 28543
rect 23661 28543 23719 28549
rect 23431 28512 23612 28540
rect 23431 28509 23443 28512
rect 23385 28503 23443 28509
rect 15210 28376 20944 28404
rect 15105 28367 15163 28373
rect 20990 28364 20996 28416
rect 21048 28364 21054 28416
rect 23477 28407 23535 28413
rect 23477 28373 23489 28407
rect 23523 28404 23535 28407
rect 23584 28404 23612 28512
rect 23661 28509 23673 28543
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28509 23995 28543
rect 23937 28503 23995 28509
rect 23523 28376 23612 28404
rect 24121 28407 24179 28413
rect 23523 28373 23535 28376
rect 23477 28367 23535 28373
rect 24121 28373 24133 28407
rect 24167 28404 24179 28407
rect 25130 28404 25136 28416
rect 24167 28376 25136 28404
rect 24167 28373 24179 28376
rect 24121 28367 24179 28373
rect 25130 28364 25136 28376
rect 25188 28364 25194 28416
rect 1104 28314 25000 28336
rect 1104 28262 6884 28314
rect 6936 28262 6948 28314
rect 7000 28262 7012 28314
rect 7064 28262 7076 28314
rect 7128 28262 7140 28314
rect 7192 28262 12818 28314
rect 12870 28262 12882 28314
rect 12934 28262 12946 28314
rect 12998 28262 13010 28314
rect 13062 28262 13074 28314
rect 13126 28262 18752 28314
rect 18804 28262 18816 28314
rect 18868 28262 18880 28314
rect 18932 28262 18944 28314
rect 18996 28262 19008 28314
rect 19060 28262 24686 28314
rect 24738 28262 24750 28314
rect 24802 28262 24814 28314
rect 24866 28262 24878 28314
rect 24930 28262 24942 28314
rect 24994 28262 25000 28314
rect 1104 28240 25000 28262
rect 2501 28203 2559 28209
rect 2501 28169 2513 28203
rect 2547 28200 2559 28203
rect 2958 28200 2964 28212
rect 2547 28172 2964 28200
rect 2547 28169 2559 28172
rect 2501 28163 2559 28169
rect 2958 28160 2964 28172
rect 3016 28160 3022 28212
rect 3326 28160 3332 28212
rect 3384 28160 3390 28212
rect 3786 28160 3792 28212
rect 3844 28160 3850 28212
rect 3878 28160 3884 28212
rect 3936 28160 3942 28212
rect 4065 28203 4123 28209
rect 4065 28169 4077 28203
rect 4111 28200 4123 28203
rect 5813 28203 5871 28209
rect 4111 28172 5764 28200
rect 4111 28169 4123 28172
rect 4065 28163 4123 28169
rect 934 28092 940 28144
rect 992 28132 998 28144
rect 992 28104 1808 28132
rect 992 28092 998 28104
rect 750 28024 756 28076
rect 808 28064 814 28076
rect 1780 28073 1808 28104
rect 2038 28092 2044 28144
rect 2096 28132 2102 28144
rect 2774 28132 2780 28144
rect 2096 28104 2780 28132
rect 2096 28092 2102 28104
rect 2774 28092 2780 28104
rect 2832 28132 2838 28144
rect 3145 28135 3203 28141
rect 2832 28104 2877 28132
rect 2832 28092 2838 28104
rect 3145 28101 3157 28135
rect 3191 28132 3203 28135
rect 3344 28132 3372 28160
rect 3804 28132 3832 28160
rect 3191 28104 3372 28132
rect 3436 28104 3832 28132
rect 3896 28132 3924 28160
rect 4338 28132 4344 28144
rect 3896 28104 4344 28132
rect 3191 28101 3203 28104
rect 3145 28095 3203 28101
rect 1489 28067 1547 28073
rect 1489 28064 1501 28067
rect 808 28036 1501 28064
rect 808 28024 814 28036
rect 1489 28033 1501 28036
rect 1535 28033 1547 28067
rect 1489 28027 1547 28033
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28033 1823 28067
rect 1765 28027 1823 28033
rect 2314 28024 2320 28076
rect 2372 28024 2378 28076
rect 3053 28067 3111 28073
rect 3053 28033 3065 28067
rect 3099 28064 3111 28067
rect 3436 28064 3464 28104
rect 4338 28092 4344 28104
rect 4396 28092 4402 28144
rect 4522 28092 4528 28144
rect 4580 28092 4586 28144
rect 4798 28092 4804 28144
rect 4856 28092 4862 28144
rect 4893 28135 4951 28141
rect 4893 28101 4905 28135
rect 4939 28132 4951 28135
rect 5534 28132 5540 28144
rect 4939 28104 5540 28132
rect 4939 28101 4951 28104
rect 4893 28095 4951 28101
rect 5534 28092 5540 28104
rect 5592 28092 5598 28144
rect 5629 28135 5687 28141
rect 5629 28101 5641 28135
rect 5675 28101 5687 28135
rect 5736 28132 5764 28172
rect 5813 28169 5825 28203
rect 5859 28200 5871 28203
rect 9122 28200 9128 28212
rect 5859 28172 9128 28200
rect 5859 28169 5871 28172
rect 5813 28163 5871 28169
rect 9122 28160 9128 28172
rect 9180 28160 9186 28212
rect 16209 28203 16267 28209
rect 9646 28172 14780 28200
rect 9646 28132 9674 28172
rect 5736 28104 9674 28132
rect 10060 28104 11652 28132
rect 5629 28095 5687 28101
rect 3099 28036 3464 28064
rect 3099 28033 3111 28036
rect 3053 28027 3111 28033
rect 3510 28024 3516 28076
rect 3568 28064 3574 28076
rect 5261 28067 5319 28073
rect 5261 28064 5273 28067
rect 3568 28036 5273 28064
rect 3568 28024 3574 28036
rect 5261 28033 5273 28036
rect 5307 28033 5319 28067
rect 5261 28027 5319 28033
rect 5350 28024 5356 28076
rect 5408 28064 5414 28076
rect 5644 28064 5672 28095
rect 5408 28036 5672 28064
rect 6639 28067 6697 28073
rect 5408 28024 5414 28036
rect 6639 28033 6651 28067
rect 6685 28064 6697 28067
rect 7558 28064 7564 28076
rect 6685 28036 7564 28064
rect 6685 28033 6697 28036
rect 6639 28027 6697 28033
rect 7558 28024 7564 28036
rect 7616 28024 7622 28076
rect 8110 28024 8116 28076
rect 8168 28064 8174 28076
rect 9950 28064 9956 28076
rect 8168 28036 9956 28064
rect 8168 28024 8174 28036
rect 9950 28024 9956 28036
rect 10008 28024 10014 28076
rect 3234 27956 3240 28008
rect 3292 27956 3298 28008
rect 4890 27956 4896 28008
rect 4948 27956 4954 28008
rect 6086 27956 6092 28008
rect 6144 27996 6150 28008
rect 6362 27996 6368 28008
rect 6144 27968 6368 27996
rect 6144 27956 6150 27968
rect 6362 27956 6368 27968
rect 6420 27956 6426 28008
rect 10060 28005 10088 28104
rect 11624 28076 11652 28104
rect 10319 28067 10377 28073
rect 10319 28033 10331 28067
rect 10365 28064 10377 28067
rect 11330 28064 11336 28076
rect 10365 28036 11336 28064
rect 10365 28033 10377 28036
rect 10319 28027 10377 28033
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 11606 28024 11612 28076
rect 11664 28064 11670 28076
rect 11790 28064 11796 28076
rect 11664 28036 11796 28064
rect 11664 28024 11670 28036
rect 11790 28024 11796 28036
rect 11848 28024 11854 28076
rect 12084 28036 13124 28064
rect 12084 28008 12112 28036
rect 10045 27999 10103 28005
rect 10045 27965 10057 27999
rect 10091 27965 10103 27999
rect 10045 27959 10103 27965
rect 12066 27956 12072 28008
rect 12124 27956 12130 28008
rect 12618 27956 12624 28008
rect 12676 27996 12682 28008
rect 12805 27999 12863 28005
rect 12805 27996 12817 27999
rect 12676 27968 12817 27996
rect 12676 27956 12682 27968
rect 12805 27965 12817 27968
rect 12851 27965 12863 27999
rect 12805 27959 12863 27965
rect 12989 27999 13047 28005
rect 12989 27965 13001 27999
rect 13035 27965 13047 27999
rect 13096 27996 13124 28036
rect 13998 28024 14004 28076
rect 14056 28024 14062 28076
rect 13725 27999 13783 28005
rect 13725 27996 13737 27999
rect 13096 27968 13737 27996
rect 12989 27959 13047 27965
rect 13725 27965 13737 27968
rect 13771 27965 13783 27999
rect 13725 27959 13783 27965
rect 1673 27931 1731 27937
rect 1673 27897 1685 27931
rect 1719 27928 1731 27931
rect 1854 27928 1860 27940
rect 1719 27900 1860 27928
rect 1719 27897 1731 27900
rect 1673 27891 1731 27897
rect 1854 27888 1860 27900
rect 1912 27888 1918 27940
rect 2682 27928 2688 27940
rect 1964 27900 2688 27928
rect 1964 27869 1992 27900
rect 2682 27888 2688 27900
rect 2740 27928 2746 27940
rect 2740 27888 2774 27928
rect 12158 27888 12164 27940
rect 12216 27928 12222 27940
rect 13004 27928 13032 27959
rect 13814 27956 13820 28008
rect 13872 28005 13878 28008
rect 13872 27999 13900 28005
rect 13888 27965 13900 27999
rect 13872 27959 13900 27965
rect 13872 27956 13878 27959
rect 12216 27900 13032 27928
rect 13449 27931 13507 27937
rect 12216 27888 12222 27900
rect 13449 27897 13461 27931
rect 13495 27897 13507 27931
rect 13449 27891 13507 27897
rect 2746 27872 2774 27888
rect 1949 27863 2007 27869
rect 1949 27829 1961 27863
rect 1995 27829 2007 27863
rect 2746 27832 2780 27872
rect 1949 27823 2007 27829
rect 2774 27820 2780 27832
rect 2832 27820 2838 27872
rect 6730 27820 6736 27872
rect 6788 27860 6794 27872
rect 7377 27863 7435 27869
rect 7377 27860 7389 27863
rect 6788 27832 7389 27860
rect 6788 27820 6794 27832
rect 7377 27829 7389 27832
rect 7423 27829 7435 27863
rect 7377 27823 7435 27829
rect 11054 27820 11060 27872
rect 11112 27820 11118 27872
rect 13464 27860 13492 27891
rect 13722 27860 13728 27872
rect 13464 27832 13728 27860
rect 13722 27820 13728 27832
rect 13780 27820 13786 27872
rect 14642 27820 14648 27872
rect 14700 27820 14706 27872
rect 14752 27860 14780 28172
rect 16209 28169 16221 28203
rect 16255 28200 16267 28203
rect 16666 28200 16672 28212
rect 16255 28172 16672 28200
rect 16255 28169 16267 28172
rect 16209 28163 16267 28169
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 19150 28160 19156 28212
rect 19208 28200 19214 28212
rect 19245 28203 19303 28209
rect 19245 28200 19257 28203
rect 19208 28172 19257 28200
rect 19208 28160 19214 28172
rect 19245 28169 19257 28172
rect 19291 28169 19303 28203
rect 19245 28163 19303 28169
rect 19518 28160 19524 28212
rect 19576 28200 19582 28212
rect 20714 28200 20720 28212
rect 19576 28172 20720 28200
rect 19576 28160 19582 28172
rect 20714 28160 20720 28172
rect 20772 28160 20778 28212
rect 20990 28160 20996 28212
rect 21048 28160 21054 28212
rect 21450 28160 21456 28212
rect 21508 28200 21514 28212
rect 22097 28203 22155 28209
rect 21508 28172 22023 28200
rect 21508 28160 21514 28172
rect 21008 28132 21036 28160
rect 17880 28104 19334 28132
rect 14918 28024 14924 28076
rect 14976 28064 14982 28076
rect 15439 28067 15497 28073
rect 15439 28064 15451 28067
rect 14976 28036 15451 28064
rect 14976 28024 14982 28036
rect 15439 28033 15451 28036
rect 15485 28033 15497 28067
rect 15439 28027 15497 28033
rect 15102 27956 15108 28008
rect 15160 27996 15166 28008
rect 15197 27999 15255 28005
rect 15197 27996 15209 27999
rect 15160 27968 15209 27996
rect 15160 27956 15166 27968
rect 15197 27965 15209 27968
rect 15243 27965 15255 27999
rect 15197 27959 15255 27965
rect 17678 27956 17684 28008
rect 17736 27996 17742 28008
rect 17880 28005 17908 28104
rect 17954 28024 17960 28076
rect 18012 28064 18018 28076
rect 18121 28067 18179 28073
rect 18121 28064 18133 28067
rect 18012 28036 18133 28064
rect 18012 28024 18018 28036
rect 18121 28033 18133 28036
rect 18167 28033 18179 28067
rect 19306 28064 19334 28104
rect 21008 28104 21864 28132
rect 19426 28064 19432 28076
rect 19306 28036 19432 28064
rect 18121 28027 18179 28033
rect 19426 28024 19432 28036
rect 19484 28024 19490 28076
rect 19702 28073 19708 28076
rect 19685 28067 19708 28073
rect 19685 28064 19697 28067
rect 19527 28036 19697 28064
rect 17865 27999 17923 28005
rect 17865 27996 17877 27999
rect 17736 27968 17877 27996
rect 17736 27956 17742 27968
rect 17865 27965 17877 27968
rect 17911 27965 17923 27999
rect 19527 27996 19555 28036
rect 19685 28033 19697 28036
rect 19685 28027 19708 28033
rect 19702 28024 19708 28027
rect 19760 28024 19766 28076
rect 20901 28067 20959 28073
rect 20901 28033 20913 28067
rect 20947 28064 20959 28067
rect 21008 28064 21036 28104
rect 21836 28073 21864 28104
rect 21995 28073 22023 28172
rect 22097 28169 22109 28203
rect 22143 28200 22155 28203
rect 22738 28200 22744 28212
rect 22143 28172 22744 28200
rect 22143 28169 22155 28172
rect 22097 28163 22155 28169
rect 22738 28160 22744 28172
rect 22796 28160 22802 28212
rect 23477 28203 23535 28209
rect 23477 28169 23489 28203
rect 23523 28169 23535 28203
rect 23477 28163 23535 28169
rect 21269 28067 21327 28073
rect 21269 28064 21281 28067
rect 20947 28036 21036 28064
rect 21100 28036 21281 28064
rect 20947 28033 20959 28036
rect 20901 28027 20959 28033
rect 17865 27959 17923 27965
rect 19444 27968 19555 27996
rect 16666 27888 16672 27940
rect 16724 27928 16730 27940
rect 17310 27928 17316 27940
rect 16724 27900 17316 27928
rect 16724 27888 16730 27900
rect 17310 27888 17316 27900
rect 17368 27888 17374 27940
rect 19444 27860 19472 27968
rect 20622 27956 20628 28008
rect 20680 27996 20686 28008
rect 21100 27996 21128 28036
rect 21269 28033 21281 28036
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 21821 28067 21879 28073
rect 21821 28033 21833 28067
rect 21867 28033 21879 28067
rect 21995 28067 22063 28073
rect 21995 28036 22017 28067
rect 21821 28027 21879 28033
rect 22005 28033 22017 28036
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22281 28067 22339 28073
rect 22281 28033 22293 28067
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 20680 27968 21128 27996
rect 21177 27999 21235 28005
rect 20680 27956 20686 27968
rect 21177 27965 21189 27999
rect 21223 27996 21235 27999
rect 21913 27999 21971 28005
rect 21913 27996 21925 27999
rect 21223 27968 21925 27996
rect 21223 27965 21235 27968
rect 21177 27959 21235 27965
rect 21913 27965 21925 27968
rect 21959 27965 21971 27999
rect 21913 27959 21971 27965
rect 20993 27931 21051 27937
rect 20993 27897 21005 27931
rect 21039 27928 21051 27931
rect 21361 27931 21419 27937
rect 21361 27928 21373 27931
rect 21039 27900 21373 27928
rect 21039 27897 21051 27900
rect 20993 27891 21051 27897
rect 21361 27897 21373 27900
rect 21407 27897 21419 27931
rect 21361 27891 21419 27897
rect 21542 27888 21548 27940
rect 21600 27928 21606 27940
rect 22296 27928 22324 28027
rect 22830 28024 22836 28076
rect 22888 28024 22894 28076
rect 22922 28024 22928 28076
rect 22980 28064 22986 28076
rect 23109 28067 23167 28073
rect 23109 28064 23121 28067
rect 22980 28036 23121 28064
rect 22980 28024 22986 28036
rect 23109 28033 23121 28036
rect 23155 28033 23167 28067
rect 23109 28027 23167 28033
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28064 23443 28067
rect 23490 28064 23518 28163
rect 23431 28036 23518 28064
rect 23661 28067 23719 28073
rect 23431 28033 23443 28036
rect 23385 28027 23443 28033
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 23676 27996 23704 28027
rect 23934 28024 23940 28076
rect 23992 28024 23998 28076
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28033 24179 28067
rect 24121 28027 24179 28033
rect 22940 27968 23704 27996
rect 22940 27937 22968 27968
rect 21600 27900 22324 27928
rect 22925 27931 22983 27937
rect 21600 27888 21606 27900
rect 22925 27897 22937 27931
rect 22971 27897 22983 27931
rect 22925 27891 22983 27897
rect 23201 27931 23259 27937
rect 23201 27897 23213 27931
rect 23247 27928 23259 27931
rect 24136 27928 24164 28027
rect 23247 27900 24164 27928
rect 23247 27897 23259 27900
rect 23201 27891 23259 27897
rect 14752 27832 19472 27860
rect 20806 27820 20812 27872
rect 20864 27820 20870 27872
rect 21085 27863 21143 27869
rect 21085 27829 21097 27863
rect 21131 27860 21143 27863
rect 22554 27860 22560 27872
rect 21131 27832 22560 27860
rect 21131 27829 21143 27832
rect 21085 27823 21143 27829
rect 22554 27820 22560 27832
rect 22612 27820 22618 27872
rect 22649 27863 22707 27869
rect 22649 27829 22661 27863
rect 22695 27860 22707 27863
rect 23474 27860 23480 27872
rect 22695 27832 23480 27860
rect 22695 27829 22707 27832
rect 22649 27823 22707 27829
rect 23474 27820 23480 27832
rect 23532 27820 23538 27872
rect 23750 27820 23756 27872
rect 23808 27820 23814 27872
rect 24394 27820 24400 27872
rect 24452 27820 24458 27872
rect 1104 27770 24840 27792
rect 1104 27718 3917 27770
rect 3969 27718 3981 27770
rect 4033 27718 4045 27770
rect 4097 27718 4109 27770
rect 4161 27718 4173 27770
rect 4225 27718 9851 27770
rect 9903 27718 9915 27770
rect 9967 27718 9979 27770
rect 10031 27718 10043 27770
rect 10095 27718 10107 27770
rect 10159 27718 15785 27770
rect 15837 27718 15849 27770
rect 15901 27718 15913 27770
rect 15965 27718 15977 27770
rect 16029 27718 16041 27770
rect 16093 27718 21719 27770
rect 21771 27718 21783 27770
rect 21835 27718 21847 27770
rect 21899 27718 21911 27770
rect 21963 27718 21975 27770
rect 22027 27718 24840 27770
rect 1104 27696 24840 27718
rect 1762 27656 1768 27668
rect 1412 27628 1768 27656
rect 1412 27529 1440 27628
rect 1762 27616 1768 27628
rect 1820 27616 1826 27668
rect 3786 27616 3792 27668
rect 3844 27656 3850 27668
rect 5258 27656 5264 27668
rect 3844 27628 5264 27656
rect 3844 27616 3850 27628
rect 5258 27616 5264 27628
rect 5316 27616 5322 27668
rect 9122 27616 9128 27668
rect 9180 27656 9186 27668
rect 20622 27656 20628 27668
rect 9180 27628 19334 27656
rect 9180 27616 9186 27628
rect 5813 27591 5871 27597
rect 5813 27557 5825 27591
rect 5859 27557 5871 27591
rect 5813 27551 5871 27557
rect 1397 27523 1455 27529
rect 1397 27489 1409 27523
rect 1443 27489 1455 27523
rect 5828 27520 5856 27551
rect 5828 27492 6210 27520
rect 1397 27483 1455 27489
rect 7926 27480 7932 27532
rect 7984 27520 7990 27532
rect 8941 27523 8999 27529
rect 8941 27520 8953 27523
rect 7984 27492 8953 27520
rect 7984 27480 7990 27492
rect 8941 27489 8953 27492
rect 8987 27489 8999 27523
rect 8941 27483 8999 27489
rect 9125 27523 9183 27529
rect 9125 27489 9137 27523
rect 9171 27520 9183 27523
rect 9214 27520 9220 27532
rect 9171 27492 9220 27520
rect 9171 27489 9183 27492
rect 9125 27483 9183 27489
rect 14 27412 20 27464
rect 72 27452 78 27464
rect 1639 27455 1697 27461
rect 1639 27452 1651 27455
rect 72 27424 1651 27452
rect 72 27412 78 27424
rect 1639 27421 1651 27424
rect 1685 27452 1697 27455
rect 2777 27455 2835 27461
rect 2777 27452 2789 27455
rect 1685 27424 1900 27452
rect 1685 27421 1697 27424
rect 1639 27415 1697 27421
rect 1872 27396 1900 27424
rect 1964 27424 2789 27452
rect 1854 27344 1860 27396
rect 1912 27344 1918 27396
rect 1118 27276 1124 27328
rect 1176 27316 1182 27328
rect 1964 27316 1992 27424
rect 2777 27421 2789 27424
rect 2823 27421 2835 27455
rect 2777 27415 2835 27421
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 4801 27455 4859 27461
rect 4801 27421 4813 27455
rect 4847 27452 4859 27455
rect 4982 27452 4988 27464
rect 4847 27424 4988 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 2682 27344 2688 27396
rect 2740 27384 2746 27396
rect 3068 27384 3096 27415
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 5075 27455 5133 27461
rect 5075 27421 5087 27455
rect 5121 27452 5133 27455
rect 6086 27452 6092 27464
rect 5121 27424 6092 27452
rect 5121 27421 5133 27424
rect 5075 27415 5133 27421
rect 6086 27412 6092 27424
rect 6144 27412 6150 27464
rect 6730 27412 6736 27464
rect 6788 27412 6794 27464
rect 6546 27384 6552 27396
rect 2740 27356 3096 27384
rect 3160 27356 6552 27384
rect 2740 27344 2746 27356
rect 1176 27288 1992 27316
rect 2409 27319 2467 27325
rect 1176 27276 1182 27288
rect 2409 27285 2421 27319
rect 2455 27316 2467 27319
rect 2498 27316 2504 27328
rect 2455 27288 2504 27316
rect 2455 27285 2467 27288
rect 2409 27279 2467 27285
rect 2498 27276 2504 27288
rect 2556 27276 2562 27328
rect 2961 27319 3019 27325
rect 2961 27285 2973 27319
rect 3007 27316 3019 27319
rect 3160 27316 3188 27356
rect 6546 27344 6552 27356
rect 6604 27344 6610 27396
rect 6638 27344 6644 27396
rect 6696 27344 6702 27396
rect 7101 27387 7159 27393
rect 7101 27353 7113 27387
rect 7147 27353 7159 27387
rect 7101 27347 7159 27353
rect 7469 27387 7527 27393
rect 7469 27353 7481 27387
rect 7515 27384 7527 27387
rect 7515 27356 8248 27384
rect 7515 27353 7527 27356
rect 7469 27347 7527 27353
rect 3007 27288 3188 27316
rect 3237 27319 3295 27325
rect 3007 27285 3019 27288
rect 2961 27279 3019 27285
rect 3237 27285 3249 27319
rect 3283 27316 3295 27319
rect 3786 27316 3792 27328
rect 3283 27288 3792 27316
rect 3283 27285 3295 27288
rect 3237 27279 3295 27285
rect 3786 27276 3792 27288
rect 3844 27276 3850 27328
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 6365 27319 6423 27325
rect 6365 27316 6377 27319
rect 4580 27288 6377 27316
rect 4580 27276 4586 27288
rect 6365 27285 6377 27288
rect 6411 27285 6423 27319
rect 6365 27279 6423 27285
rect 6454 27276 6460 27328
rect 6512 27316 6518 27328
rect 7116 27316 7144 27347
rect 8220 27328 8248 27356
rect 7282 27316 7288 27328
rect 6512 27288 7288 27316
rect 6512 27276 6518 27288
rect 7282 27276 7288 27288
rect 7340 27276 7346 27328
rect 7650 27276 7656 27328
rect 7708 27276 7714 27328
rect 8202 27276 8208 27328
rect 8260 27276 8266 27328
rect 8956 27316 8984 27483
rect 9214 27480 9220 27492
rect 9272 27480 9278 27532
rect 9582 27480 9588 27532
rect 9640 27480 9646 27532
rect 10042 27529 10048 27532
rect 9999 27523 10048 27529
rect 9999 27489 10011 27523
rect 10045 27489 10048 27523
rect 9999 27483 10048 27489
rect 10042 27480 10048 27483
rect 10100 27480 10106 27532
rect 10137 27523 10195 27529
rect 10137 27489 10149 27523
rect 10183 27520 10195 27523
rect 10318 27520 10324 27532
rect 10183 27492 10324 27520
rect 10183 27489 10195 27492
rect 10137 27483 10195 27489
rect 10318 27480 10324 27492
rect 10376 27480 10382 27532
rect 12802 27480 12808 27532
rect 12860 27520 12866 27532
rect 15102 27520 15108 27532
rect 12860 27492 15108 27520
rect 12860 27480 12866 27492
rect 9858 27412 9864 27464
rect 9916 27412 9922 27464
rect 11514 27412 11520 27464
rect 11572 27412 11578 27464
rect 11775 27455 11833 27461
rect 11775 27421 11787 27455
rect 11821 27452 11833 27455
rect 12250 27452 12256 27464
rect 11821 27424 12256 27452
rect 11821 27421 11833 27424
rect 11775 27415 11833 27421
rect 10778 27344 10784 27396
rect 10836 27344 10842 27396
rect 11422 27344 11428 27396
rect 11480 27384 11486 27396
rect 11790 27384 11818 27415
rect 12250 27412 12256 27424
rect 12308 27412 12314 27464
rect 13814 27384 13820 27396
rect 11480 27356 11818 27384
rect 12360 27356 13820 27384
rect 11480 27344 11486 27356
rect 12360 27316 12388 27356
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 8956 27288 12388 27316
rect 12434 27276 12440 27328
rect 12492 27316 12498 27328
rect 12529 27319 12587 27325
rect 12529 27316 12541 27319
rect 12492 27288 12541 27316
rect 12492 27276 12498 27288
rect 12529 27285 12541 27288
rect 12575 27285 12587 27319
rect 14568 27316 14596 27492
rect 15102 27480 15108 27492
rect 15160 27520 15166 27532
rect 16206 27520 16212 27532
rect 15160 27492 16212 27520
rect 15160 27480 15166 27492
rect 16206 27480 16212 27492
rect 16264 27480 16270 27532
rect 17310 27480 17316 27532
rect 17368 27520 17374 27532
rect 17589 27523 17647 27529
rect 17589 27520 17601 27523
rect 17368 27492 17601 27520
rect 17368 27480 17374 27492
rect 17589 27489 17601 27492
rect 17635 27489 17647 27523
rect 17589 27483 17647 27489
rect 14642 27412 14648 27464
rect 14700 27452 14706 27464
rect 15197 27455 15255 27461
rect 15197 27452 15209 27455
rect 14700 27424 15209 27452
rect 14700 27412 14706 27424
rect 15197 27421 15209 27424
rect 15243 27421 15255 27455
rect 15197 27415 15255 27421
rect 16483 27445 16541 27451
rect 16483 27411 16495 27445
rect 16529 27428 16541 27445
rect 16529 27411 16620 27428
rect 17218 27412 17224 27464
rect 17276 27452 17282 27464
rect 17831 27455 17889 27461
rect 17831 27452 17843 27455
rect 17276 27424 17843 27452
rect 17276 27412 17282 27424
rect 17831 27421 17843 27424
rect 17877 27421 17889 27455
rect 19306 27452 19334 27628
rect 19996 27628 20628 27656
rect 19996 27597 20024 27628
rect 20622 27616 20628 27628
rect 20680 27616 20686 27668
rect 20901 27659 20959 27665
rect 20901 27625 20913 27659
rect 20947 27656 20959 27659
rect 21450 27656 21456 27668
rect 20947 27628 21456 27656
rect 20947 27625 20959 27628
rect 20901 27619 20959 27625
rect 21450 27616 21456 27628
rect 21508 27616 21514 27668
rect 22557 27659 22615 27665
rect 22557 27625 22569 27659
rect 22603 27656 22615 27659
rect 22830 27656 22836 27668
rect 22603 27628 22836 27656
rect 22603 27625 22615 27628
rect 22557 27619 22615 27625
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 23569 27659 23627 27665
rect 23569 27625 23581 27659
rect 23615 27656 23627 27659
rect 23934 27656 23940 27668
rect 23615 27628 23940 27656
rect 23615 27625 23627 27628
rect 23569 27619 23627 27625
rect 23934 27616 23940 27628
rect 23992 27616 23998 27668
rect 19981 27591 20039 27597
rect 19981 27557 19993 27591
rect 20027 27557 20039 27591
rect 19981 27551 20039 27557
rect 22741 27591 22799 27597
rect 22741 27557 22753 27591
rect 22787 27588 22799 27591
rect 23109 27591 23167 27597
rect 23109 27588 23121 27591
rect 22787 27560 23121 27588
rect 22787 27557 22799 27560
rect 22741 27551 22799 27557
rect 23109 27557 23121 27560
rect 23155 27557 23167 27591
rect 23109 27551 23167 27557
rect 19426 27480 19432 27532
rect 19484 27520 19490 27532
rect 22925 27523 22983 27529
rect 19484 27492 21220 27520
rect 19484 27480 19490 27492
rect 21192 27464 21220 27492
rect 22925 27489 22937 27523
rect 22971 27520 22983 27523
rect 23385 27523 23443 27529
rect 23385 27520 23397 27523
rect 22971 27492 23397 27520
rect 22971 27489 22983 27492
rect 22925 27483 22983 27489
rect 23385 27489 23397 27492
rect 23431 27489 23443 27523
rect 23385 27483 23443 27489
rect 23584 27492 23980 27520
rect 23584 27464 23612 27492
rect 19306 27424 19656 27452
rect 17831 27415 17889 27421
rect 16483 27405 16620 27411
rect 16500 27400 16620 27405
rect 14642 27316 14648 27328
rect 14568 27288 14648 27316
rect 12529 27279 12587 27285
rect 14642 27276 14648 27288
rect 14700 27276 14706 27328
rect 15010 27276 15016 27328
rect 15068 27276 15074 27328
rect 16482 27276 16488 27328
rect 16540 27316 16546 27328
rect 16592 27316 16620 27400
rect 19628 27384 19656 27424
rect 19702 27412 19708 27464
rect 19760 27452 19766 27464
rect 20165 27455 20223 27461
rect 20165 27452 20177 27455
rect 19760 27424 20177 27452
rect 19760 27412 19766 27424
rect 20165 27421 20177 27424
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 20806 27412 20812 27464
rect 20864 27452 20870 27464
rect 21085 27455 21143 27461
rect 21085 27452 21097 27455
rect 20864 27424 21097 27452
rect 20864 27412 20870 27424
rect 21085 27421 21097 27424
rect 21131 27421 21143 27455
rect 21085 27415 21143 27421
rect 21174 27412 21180 27464
rect 21232 27412 21238 27464
rect 22649 27455 22707 27461
rect 22649 27421 22661 27455
rect 22695 27421 22707 27455
rect 22649 27415 22707 27421
rect 21422 27387 21480 27393
rect 21422 27384 21434 27387
rect 19628 27356 21434 27384
rect 21422 27353 21434 27356
rect 21468 27384 21480 27387
rect 21542 27384 21548 27396
rect 21468 27356 21548 27384
rect 21468 27353 21480 27356
rect 21422 27347 21480 27353
rect 21542 27344 21548 27356
rect 21600 27344 21606 27396
rect 22664 27384 22692 27415
rect 22738 27412 22744 27464
rect 22796 27452 22802 27464
rect 23017 27455 23075 27461
rect 23017 27452 23029 27455
rect 22796 27424 23029 27452
rect 22796 27412 22802 27424
rect 23017 27421 23029 27424
rect 23063 27421 23075 27455
rect 23017 27415 23075 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 22830 27384 22836 27396
rect 22664 27356 22836 27384
rect 22830 27344 22836 27356
rect 22888 27384 22894 27396
rect 23308 27384 23336 27415
rect 23474 27412 23480 27464
rect 23532 27412 23538 27464
rect 23566 27412 23572 27464
rect 23624 27412 23630 27464
rect 23952 27461 23980 27492
rect 23753 27455 23811 27461
rect 23753 27421 23765 27455
rect 23799 27421 23811 27455
rect 23753 27415 23811 27421
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 22888 27356 23336 27384
rect 22888 27344 22894 27356
rect 16540 27288 16620 27316
rect 16540 27276 16546 27288
rect 17218 27276 17224 27328
rect 17276 27276 17282 27328
rect 17862 27276 17868 27328
rect 17920 27316 17926 27328
rect 18601 27319 18659 27325
rect 18601 27316 18613 27319
rect 17920 27288 18613 27316
rect 17920 27276 17926 27288
rect 18601 27285 18613 27288
rect 18647 27285 18659 27319
rect 18601 27279 18659 27285
rect 22738 27276 22744 27328
rect 22796 27316 22802 27328
rect 22925 27319 22983 27325
rect 22925 27316 22937 27319
rect 22796 27288 22937 27316
rect 22796 27276 22802 27288
rect 22925 27285 22937 27288
rect 22971 27285 22983 27319
rect 22925 27279 22983 27285
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 23768 27316 23796 27415
rect 23072 27288 23796 27316
rect 24121 27319 24179 27325
rect 23072 27276 23078 27288
rect 24121 27285 24133 27319
rect 24167 27316 24179 27319
rect 25130 27316 25136 27328
rect 24167 27288 25136 27316
rect 24167 27285 24179 27288
rect 24121 27279 24179 27285
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 1104 27226 25000 27248
rect 1104 27174 6884 27226
rect 6936 27174 6948 27226
rect 7000 27174 7012 27226
rect 7064 27174 7076 27226
rect 7128 27174 7140 27226
rect 7192 27174 12818 27226
rect 12870 27174 12882 27226
rect 12934 27174 12946 27226
rect 12998 27174 13010 27226
rect 13062 27174 13074 27226
rect 13126 27174 18752 27226
rect 18804 27174 18816 27226
rect 18868 27174 18880 27226
rect 18932 27174 18944 27226
rect 18996 27174 19008 27226
rect 19060 27174 24686 27226
rect 24738 27174 24750 27226
rect 24802 27174 24814 27226
rect 24866 27174 24878 27226
rect 24930 27174 24942 27226
rect 24994 27174 25000 27226
rect 1104 27152 25000 27174
rect 1210 27072 1216 27124
rect 1268 27112 1274 27124
rect 1268 27084 3556 27112
rect 1268 27072 1274 27084
rect 2038 27004 2044 27056
rect 2096 27004 2102 27056
rect 2682 27044 2688 27056
rect 2148 27016 2688 27044
rect 1302 26936 1308 26988
rect 1360 26976 1366 26988
rect 2148 26976 2176 27016
rect 2682 27004 2688 27016
rect 2740 27004 2746 27056
rect 3050 27004 3056 27056
rect 3108 27004 3114 27056
rect 3142 27004 3148 27056
rect 3200 27004 3206 27056
rect 1360 26948 2176 26976
rect 1360 26936 1366 26948
rect 2314 26936 2320 26988
rect 2372 26936 2378 26988
rect 2406 26936 2412 26988
rect 2464 26936 2470 26988
rect 2777 26979 2835 26985
rect 2777 26945 2789 26979
rect 2823 26976 2835 26979
rect 2958 26976 2964 26988
rect 2823 26948 2964 26976
rect 2823 26945 2835 26948
rect 2777 26939 2835 26945
rect 2958 26936 2964 26948
rect 3016 26936 3022 26988
rect 3068 26976 3096 27004
rect 3068 26948 3188 26976
rect 2498 26868 2504 26920
rect 2556 26868 2562 26920
rect 3160 26840 3188 26948
rect 3326 26936 3332 26988
rect 3384 26936 3390 26988
rect 3528 26985 3556 27084
rect 6546 27072 6552 27124
rect 6604 27112 6610 27124
rect 8757 27115 8815 27121
rect 6604 27084 8524 27112
rect 6604 27072 6610 27084
rect 5350 27004 5356 27056
rect 5408 27044 5414 27056
rect 8496 27044 8524 27084
rect 8757 27081 8769 27115
rect 8803 27112 8815 27115
rect 9582 27112 9588 27124
rect 8803 27084 9588 27112
rect 8803 27081 8815 27084
rect 8757 27075 8815 27081
rect 9582 27072 9588 27084
rect 9640 27072 9646 27124
rect 11514 27072 11520 27124
rect 11572 27112 11578 27124
rect 12710 27112 12716 27124
rect 11572 27084 12716 27112
rect 11572 27072 11578 27084
rect 12710 27072 12716 27084
rect 12768 27072 12774 27124
rect 15194 27112 15200 27124
rect 13004 27084 15200 27112
rect 13004 27044 13032 27084
rect 15194 27072 15200 27084
rect 15252 27072 15258 27124
rect 20714 27112 20720 27124
rect 16868 27084 20720 27112
rect 5408 27016 8432 27044
rect 8496 27016 13032 27044
rect 14645 27047 14703 27053
rect 5408 27004 5414 27016
rect 4799 26989 4857 26995
rect 3513 26979 3571 26985
rect 3513 26945 3525 26979
rect 3559 26945 3571 26979
rect 3513 26939 3571 26945
rect 3602 26936 3608 26988
rect 3660 26976 3666 26988
rect 4522 26976 4528 26988
rect 3660 26948 4528 26976
rect 3660 26936 3666 26948
rect 4522 26936 4528 26948
rect 4580 26936 4586 26988
rect 4799 26955 4811 26989
rect 4845 26986 4857 26989
rect 4890 26986 4896 26988
rect 4845 26958 4896 26986
rect 4845 26955 4857 26958
rect 4799 26949 4857 26955
rect 4890 26936 4896 26958
rect 4948 26936 4954 26988
rect 7742 26936 7748 26988
rect 7800 26936 7806 26988
rect 8019 26979 8077 26985
rect 8019 26945 8031 26979
rect 8065 26976 8077 26979
rect 8110 26976 8116 26988
rect 8065 26948 8116 26976
rect 8065 26945 8077 26948
rect 8019 26939 8077 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 3344 26908 3372 26936
rect 3620 26908 3648 26936
rect 3344 26880 3648 26908
rect 5534 26868 5540 26920
rect 5592 26868 5598 26920
rect 8404 26908 8432 27016
rect 14645 27013 14657 27047
rect 14691 27044 14703 27047
rect 16868 27044 16896 27084
rect 20714 27072 20720 27084
rect 20772 27072 20778 27124
rect 20806 27072 20812 27124
rect 20864 27112 20870 27124
rect 20864 27084 22094 27112
rect 20864 27072 20870 27084
rect 14691 27016 16896 27044
rect 14691 27013 14703 27016
rect 14645 27007 14703 27013
rect 18598 27004 18604 27056
rect 18656 27044 18662 27056
rect 19610 27044 19616 27056
rect 18656 27016 19616 27044
rect 18656 27004 18662 27016
rect 19610 27004 19616 27016
rect 19668 27004 19674 27056
rect 22066 27044 22094 27084
rect 22830 27072 22836 27124
rect 22888 27072 22894 27124
rect 23014 27072 23020 27124
rect 23072 27072 23078 27124
rect 23293 27115 23351 27121
rect 23293 27081 23305 27115
rect 23339 27112 23351 27115
rect 23566 27112 23572 27124
rect 23339 27084 23572 27112
rect 23339 27081 23351 27084
rect 23293 27075 23351 27081
rect 23566 27072 23572 27084
rect 23624 27072 23630 27124
rect 23750 27072 23756 27124
rect 23808 27072 23814 27124
rect 23937 27115 23995 27121
rect 23937 27081 23949 27115
rect 23983 27081 23995 27115
rect 23937 27075 23995 27081
rect 23032 27044 23060 27072
rect 23768 27044 23796 27072
rect 22066 27016 23060 27044
rect 23492 27016 23796 27044
rect 23952 27044 23980 27075
rect 23952 27016 24256 27044
rect 10410 26936 10416 26988
rect 10468 26976 10474 26988
rect 11606 26976 11612 26988
rect 10468 26948 11612 26976
rect 10468 26936 10474 26948
rect 11606 26936 11612 26948
rect 11664 26936 11670 26988
rect 12710 26936 12716 26988
rect 12768 26976 12774 26988
rect 12989 26979 13047 26985
rect 12989 26976 13001 26979
rect 12768 26948 13001 26976
rect 12768 26936 12774 26948
rect 12989 26945 13001 26948
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 13814 26936 13820 26988
rect 13872 26985 13878 26988
rect 13872 26979 13900 26985
rect 13888 26945 13900 26979
rect 13872 26939 13900 26945
rect 15011 26979 15069 26985
rect 15011 26945 15023 26979
rect 15057 26976 15069 26979
rect 15102 26976 15108 26988
rect 15057 26948 15108 26976
rect 15057 26945 15069 26948
rect 15011 26939 15069 26945
rect 13872 26936 13878 26939
rect 15102 26936 15108 26948
rect 15160 26936 15166 26988
rect 16669 26979 16727 26985
rect 16669 26945 16681 26979
rect 16715 26976 16727 26979
rect 16758 26976 16764 26988
rect 16715 26948 16764 26976
rect 16715 26945 16727 26948
rect 16669 26939 16727 26945
rect 12618 26908 12624 26920
rect 8404 26880 12624 26908
rect 12618 26868 12624 26880
rect 12676 26908 12682 26920
rect 12805 26911 12863 26917
rect 12805 26908 12817 26911
rect 12676 26880 12817 26908
rect 12676 26868 12682 26880
rect 12805 26877 12817 26880
rect 12851 26908 12863 26911
rect 12894 26908 12900 26920
rect 12851 26880 12900 26908
rect 12851 26877 12863 26880
rect 12805 26871 12863 26877
rect 12894 26868 12900 26880
rect 12952 26868 12958 26920
rect 13446 26868 13452 26920
rect 13504 26868 13510 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 13556 26880 13737 26908
rect 3329 26843 3387 26849
rect 3329 26840 3341 26843
rect 3160 26812 3341 26840
rect 3329 26809 3341 26812
rect 3375 26809 3387 26843
rect 3329 26803 3387 26809
rect 3697 26843 3755 26849
rect 3697 26809 3709 26843
rect 3743 26809 3755 26843
rect 3697 26803 3755 26809
rect 3712 26772 3740 26803
rect 5350 26772 5356 26784
rect 3712 26744 5356 26772
rect 5350 26732 5356 26744
rect 5408 26732 5414 26784
rect 5552 26781 5580 26868
rect 5810 26800 5816 26852
rect 5868 26840 5874 26852
rect 5868 26812 7880 26840
rect 5868 26800 5874 26812
rect 5537 26775 5595 26781
rect 5537 26741 5549 26775
rect 5583 26741 5595 26775
rect 7852 26772 7880 26812
rect 9306 26800 9312 26852
rect 9364 26840 9370 26852
rect 13262 26840 13268 26852
rect 9364 26812 13268 26840
rect 9364 26800 9370 26812
rect 13262 26800 13268 26812
rect 13320 26840 13326 26852
rect 13556 26840 13584 26880
rect 13725 26877 13737 26880
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 14001 26911 14059 26917
rect 14001 26877 14013 26911
rect 14047 26908 14059 26911
rect 14047 26880 14596 26908
rect 14047 26877 14059 26880
rect 14001 26871 14059 26877
rect 13320 26812 13584 26840
rect 13320 26800 13326 26812
rect 9766 26772 9772 26784
rect 7852 26744 9772 26772
rect 5537 26735 5595 26741
rect 9766 26732 9772 26744
rect 9824 26772 9830 26784
rect 11238 26772 11244 26784
rect 9824 26744 11244 26772
rect 9824 26732 9830 26744
rect 11238 26732 11244 26744
rect 11296 26732 11302 26784
rect 14568 26772 14596 26880
rect 14642 26868 14648 26920
rect 14700 26908 14706 26920
rect 14737 26911 14795 26917
rect 14737 26908 14749 26911
rect 14700 26880 14749 26908
rect 14700 26868 14706 26880
rect 14737 26877 14749 26880
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 15749 26775 15807 26781
rect 15749 26772 15761 26775
rect 14568 26744 15761 26772
rect 15749 26741 15761 26744
rect 15795 26741 15807 26775
rect 16684 26772 16712 26939
rect 16758 26936 16764 26948
rect 16816 26936 16822 26988
rect 17862 26936 17868 26988
rect 17920 26936 17926 26988
rect 22095 26979 22153 26985
rect 22095 26945 22107 26979
rect 22141 26976 22153 26979
rect 22186 26976 22192 26988
rect 22141 26948 22192 26976
rect 22141 26945 22153 26948
rect 22095 26939 22153 26945
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 23492 26985 23520 27016
rect 23477 26979 23535 26985
rect 23477 26945 23489 26979
rect 23523 26945 23535 26979
rect 23477 26939 23535 26945
rect 23750 26936 23756 26988
rect 23808 26936 23814 26988
rect 24228 26985 24256 27016
rect 24121 26979 24179 26985
rect 24121 26945 24133 26979
rect 24167 26945 24179 26979
rect 24121 26939 24179 26945
rect 24213 26979 24271 26985
rect 24213 26945 24225 26979
rect 24259 26945 24271 26979
rect 24213 26939 24271 26945
rect 16850 26868 16856 26920
rect 16908 26868 16914 26920
rect 17218 26868 17224 26920
rect 17276 26908 17282 26920
rect 17313 26911 17371 26917
rect 17313 26908 17325 26911
rect 17276 26880 17325 26908
rect 17276 26868 17282 26880
rect 17313 26877 17325 26880
rect 17359 26877 17371 26911
rect 17313 26871 17371 26877
rect 17586 26868 17592 26920
rect 17644 26868 17650 26920
rect 17770 26917 17776 26920
rect 17727 26911 17776 26917
rect 17727 26877 17739 26911
rect 17773 26877 17776 26911
rect 17727 26871 17776 26877
rect 17770 26868 17776 26871
rect 17828 26868 17834 26920
rect 19978 26868 19984 26920
rect 20036 26908 20042 26920
rect 21542 26908 21548 26920
rect 20036 26880 21548 26908
rect 20036 26868 20042 26880
rect 21542 26868 21548 26880
rect 21600 26908 21606 26920
rect 21821 26911 21879 26917
rect 21821 26908 21833 26911
rect 21600 26880 21833 26908
rect 21600 26868 21606 26880
rect 21821 26877 21833 26880
rect 21867 26877 21879 26911
rect 24136 26908 24164 26939
rect 21821 26871 21879 26877
rect 23584 26880 24164 26908
rect 23584 26849 23612 26880
rect 23569 26843 23627 26849
rect 23569 26809 23581 26843
rect 23615 26809 23627 26843
rect 23569 26803 23627 26809
rect 17402 26772 17408 26784
rect 16684 26744 17408 26772
rect 15749 26735 15807 26741
rect 17402 26732 17408 26744
rect 17460 26732 17466 26784
rect 18509 26775 18567 26781
rect 18509 26741 18521 26775
rect 18555 26772 18567 26775
rect 19426 26772 19432 26784
rect 18555 26744 19432 26772
rect 18555 26741 18567 26744
rect 18509 26735 18567 26741
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 22738 26732 22744 26784
rect 22796 26772 22802 26784
rect 23934 26772 23940 26784
rect 22796 26744 23940 26772
rect 22796 26732 22802 26744
rect 23934 26732 23940 26744
rect 23992 26732 23998 26784
rect 24394 26732 24400 26784
rect 24452 26732 24458 26784
rect 25314 26704 25320 26716
rect 1104 26682 24840 26704
rect 1104 26630 3917 26682
rect 3969 26630 3981 26682
rect 4033 26630 4045 26682
rect 4097 26630 4109 26682
rect 4161 26630 4173 26682
rect 4225 26630 9851 26682
rect 9903 26630 9915 26682
rect 9967 26630 9979 26682
rect 10031 26630 10043 26682
rect 10095 26630 10107 26682
rect 10159 26630 15785 26682
rect 15837 26630 15849 26682
rect 15901 26630 15913 26682
rect 15965 26630 15977 26682
rect 16029 26630 16041 26682
rect 16093 26630 21719 26682
rect 21771 26630 21783 26682
rect 21835 26630 21847 26682
rect 21899 26630 21911 26682
rect 21963 26630 21975 26682
rect 22027 26630 24840 26682
rect 1104 26608 24840 26630
rect 25240 26676 25320 26704
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 2593 26571 2651 26577
rect 2593 26568 2605 26571
rect 2464 26540 2605 26568
rect 2464 26528 2470 26540
rect 2593 26537 2605 26540
rect 2639 26537 2651 26571
rect 2593 26531 2651 26537
rect 3234 26528 3240 26580
rect 3292 26528 3298 26580
rect 3329 26571 3387 26577
rect 3329 26537 3341 26571
rect 3375 26568 3387 26571
rect 3510 26568 3516 26580
rect 3375 26540 3516 26568
rect 3375 26537 3387 26540
rect 3329 26531 3387 26537
rect 3510 26528 3516 26540
rect 3568 26528 3574 26580
rect 4249 26571 4307 26577
rect 4249 26537 4261 26571
rect 4295 26568 4307 26571
rect 4295 26540 10916 26568
rect 4295 26537 4307 26540
rect 4249 26531 4307 26537
rect 2958 26460 2964 26512
rect 3016 26500 3022 26512
rect 3602 26500 3608 26512
rect 3016 26472 3608 26500
rect 3016 26460 3022 26472
rect 3602 26460 3608 26472
rect 3660 26460 3666 26512
rect 4522 26460 4528 26512
rect 4580 26500 4586 26512
rect 4580 26472 6592 26500
rect 4580 26460 4586 26472
rect 6564 26444 6592 26472
rect 9674 26460 9680 26512
rect 9732 26500 9738 26512
rect 9861 26503 9919 26509
rect 9861 26500 9873 26503
rect 9732 26472 9873 26500
rect 9732 26460 9738 26472
rect 9861 26469 9873 26472
rect 9907 26469 9919 26503
rect 10888 26500 10916 26540
rect 10962 26528 10968 26580
rect 11020 26568 11026 26580
rect 11057 26571 11115 26577
rect 11057 26568 11069 26571
rect 11020 26540 11069 26568
rect 11020 26528 11026 26540
rect 11057 26537 11069 26540
rect 11103 26537 11115 26571
rect 11057 26531 11115 26537
rect 12894 26528 12900 26580
rect 12952 26568 12958 26580
rect 13630 26568 13636 26580
rect 12952 26540 13636 26568
rect 12952 26528 12958 26540
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 15838 26568 15844 26580
rect 15028 26540 15844 26568
rect 11146 26500 11152 26512
rect 10888 26472 11152 26500
rect 9861 26463 9919 26469
rect 11146 26460 11152 26472
rect 11204 26460 11210 26512
rect 12805 26503 12863 26509
rect 12805 26469 12817 26503
rect 12851 26500 12863 26503
rect 15028 26500 15056 26540
rect 15838 26528 15844 26540
rect 15896 26528 15902 26580
rect 15933 26571 15991 26577
rect 15933 26537 15945 26571
rect 15979 26537 15991 26571
rect 15933 26531 15991 26537
rect 15948 26500 15976 26531
rect 16022 26528 16028 26580
rect 16080 26568 16086 26580
rect 20254 26568 20260 26580
rect 16080 26540 20260 26568
rect 16080 26528 16086 26540
rect 20254 26528 20260 26540
rect 20312 26528 20318 26580
rect 20438 26528 20444 26580
rect 20496 26528 20502 26580
rect 22741 26571 22799 26577
rect 22741 26537 22753 26571
rect 22787 26568 22799 26571
rect 23750 26568 23756 26580
rect 22787 26540 23756 26568
rect 22787 26537 22799 26540
rect 22741 26531 22799 26537
rect 23750 26528 23756 26540
rect 23808 26528 23814 26580
rect 12851 26472 15056 26500
rect 15856 26472 15976 26500
rect 19061 26503 19119 26509
rect 12851 26469 12863 26472
rect 12805 26463 12863 26469
rect 2314 26392 2320 26444
rect 2372 26432 2378 26444
rect 4338 26432 4344 26444
rect 2372 26404 4344 26432
rect 2372 26392 2378 26404
rect 4338 26392 4344 26404
rect 4396 26432 4402 26444
rect 6086 26432 6092 26444
rect 4396 26404 6092 26432
rect 4396 26392 4402 26404
rect 6086 26392 6092 26404
rect 6144 26392 6150 26444
rect 6546 26392 6552 26444
rect 6604 26392 6610 26444
rect 9217 26435 9275 26441
rect 9217 26401 9229 26435
rect 9263 26432 9275 26435
rect 9950 26432 9956 26444
rect 9263 26404 9956 26432
rect 9263 26401 9275 26404
rect 9217 26395 9275 26401
rect 9950 26392 9956 26404
rect 10008 26392 10014 26444
rect 10318 26441 10324 26444
rect 10275 26435 10324 26441
rect 10275 26401 10287 26435
rect 10321 26401 10324 26435
rect 10275 26395 10324 26401
rect 10318 26392 10324 26395
rect 10376 26392 10382 26444
rect 10778 26392 10784 26444
rect 10836 26432 10842 26444
rect 10836 26404 11008 26432
rect 10836 26392 10842 26404
rect 1486 26324 1492 26376
rect 1544 26364 1550 26376
rect 1581 26367 1639 26373
rect 1581 26364 1593 26367
rect 1544 26336 1593 26364
rect 1544 26324 1550 26336
rect 1581 26333 1593 26336
rect 1627 26364 1639 26367
rect 1762 26364 1768 26376
rect 1627 26336 1768 26364
rect 1627 26333 1639 26336
rect 1581 26327 1639 26333
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 1855 26367 1913 26373
rect 1855 26333 1867 26367
rect 1901 26364 1913 26367
rect 2958 26364 2964 26376
rect 1901 26336 2964 26364
rect 1901 26333 1913 26336
rect 1855 26327 1913 26333
rect 2958 26324 2964 26336
rect 3016 26364 3022 26376
rect 3234 26364 3240 26376
rect 3016 26336 3240 26364
rect 3016 26324 3022 26336
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 3510 26324 3516 26376
rect 3568 26324 3574 26376
rect 3789 26367 3847 26373
rect 3789 26333 3801 26367
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 3804 26296 3832 26327
rect 4062 26324 4068 26376
rect 4120 26324 4126 26376
rect 4890 26324 4896 26376
rect 4948 26364 4954 26376
rect 5534 26364 5540 26376
rect 4948 26336 5540 26364
rect 4948 26324 4954 26336
rect 5534 26324 5540 26336
rect 5592 26324 5598 26376
rect 6822 26364 6828 26376
rect 6783 26336 6828 26364
rect 6822 26324 6828 26336
rect 6880 26364 6886 26376
rect 7834 26364 7840 26376
rect 6880 26336 7840 26364
rect 6880 26324 6886 26336
rect 7834 26324 7840 26336
rect 7892 26324 7898 26376
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 9364 26336 9413 26364
rect 9364 26324 9370 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 9401 26327 9459 26333
rect 10134 26324 10140 26376
rect 10192 26324 10198 26376
rect 10410 26324 10416 26376
rect 10468 26324 10474 26376
rect 10980 26364 11008 26404
rect 11054 26392 11060 26444
rect 11112 26432 11118 26444
rect 15856 26432 15884 26472
rect 19061 26469 19073 26503
rect 19107 26500 19119 26503
rect 19518 26500 19524 26512
rect 19107 26472 19524 26500
rect 19107 26469 19119 26472
rect 19061 26463 19119 26469
rect 19518 26460 19524 26472
rect 19576 26460 19582 26512
rect 20456 26500 20484 26528
rect 25240 26512 25268 26676
rect 25314 26664 25320 26676
rect 25372 26664 25378 26716
rect 20456 26472 23336 26500
rect 15930 26432 15936 26444
rect 11112 26404 11362 26432
rect 15856 26404 15936 26432
rect 11112 26392 11118 26404
rect 15930 26392 15936 26404
rect 15988 26432 15994 26444
rect 16301 26435 16359 26441
rect 16301 26432 16313 26435
rect 15988 26404 16313 26432
rect 15988 26392 15994 26404
rect 16301 26401 16313 26404
rect 16347 26401 16359 26435
rect 16301 26395 16359 26401
rect 18690 26392 18696 26444
rect 18748 26432 18754 26444
rect 23308 26432 23336 26472
rect 25222 26460 25228 26512
rect 25280 26460 25286 26512
rect 18748 26404 22094 26432
rect 23308 26404 23888 26432
rect 18748 26392 18754 26404
rect 11793 26367 11851 26373
rect 11793 26364 11805 26367
rect 10980 26336 11805 26364
rect 11793 26333 11805 26336
rect 11839 26364 11851 26367
rect 11839 26336 12388 26364
rect 11839 26333 11851 26336
rect 11793 26327 11851 26333
rect 12360 26308 12388 26336
rect 13906 26324 13912 26376
rect 13964 26364 13970 26376
rect 14734 26364 14740 26376
rect 13964 26336 14740 26364
rect 13964 26324 13970 26336
rect 14734 26324 14740 26336
rect 14792 26364 14798 26376
rect 14921 26367 14979 26373
rect 14921 26364 14933 26367
rect 14792 26336 14933 26364
rect 14792 26324 14798 26336
rect 14921 26333 14933 26336
rect 14967 26333 14979 26367
rect 14921 26327 14979 26333
rect 15179 26337 15237 26343
rect 9122 26296 9128 26308
rect 2746 26268 3832 26296
rect 3988 26268 9128 26296
rect 566 26188 572 26240
rect 624 26228 630 26240
rect 2038 26228 2044 26240
rect 624 26200 2044 26228
rect 624 26188 630 26200
rect 2038 26188 2044 26200
rect 2096 26188 2102 26240
rect 2590 26188 2596 26240
rect 2648 26228 2654 26240
rect 2746 26228 2774 26268
rect 3988 26237 4016 26268
rect 9122 26256 9128 26268
rect 9180 26256 9186 26308
rect 11238 26256 11244 26308
rect 11296 26296 11302 26308
rect 11517 26299 11575 26305
rect 11517 26296 11529 26299
rect 11296 26268 11529 26296
rect 11296 26256 11302 26268
rect 11517 26265 11529 26268
rect 11563 26265 11575 26299
rect 11517 26259 11575 26265
rect 11882 26256 11888 26308
rect 11940 26256 11946 26308
rect 12250 26256 12256 26308
rect 12308 26256 12314 26308
rect 12342 26256 12348 26308
rect 12400 26256 12406 26308
rect 15179 26303 15191 26337
rect 15225 26334 15237 26337
rect 15225 26303 15238 26334
rect 15654 26324 15660 26376
rect 15712 26364 15718 26376
rect 16485 26367 16543 26373
rect 16485 26364 16497 26367
rect 15712 26336 16497 26364
rect 15712 26324 15718 26336
rect 16485 26333 16497 26336
rect 16531 26333 16543 26367
rect 16853 26367 16911 26373
rect 16853 26364 16865 26367
rect 16485 26327 16543 26333
rect 16574 26336 16865 26364
rect 15179 26297 15238 26303
rect 15210 26296 15238 26297
rect 15838 26296 15844 26308
rect 12544 26268 12756 26296
rect 15210 26268 15844 26296
rect 2648 26200 2774 26228
rect 3973 26231 4031 26237
rect 2648 26188 2654 26200
rect 3973 26197 3985 26231
rect 4019 26197 4031 26231
rect 3973 26191 4031 26197
rect 4982 26188 4988 26240
rect 5040 26228 5046 26240
rect 6178 26228 6184 26240
rect 5040 26200 6184 26228
rect 5040 26188 5046 26200
rect 6178 26188 6184 26200
rect 6236 26188 6242 26240
rect 7558 26188 7564 26240
rect 7616 26188 7622 26240
rect 7834 26188 7840 26240
rect 7892 26228 7898 26240
rect 12544 26228 12572 26268
rect 7892 26200 12572 26228
rect 7892 26188 7898 26200
rect 12618 26188 12624 26240
rect 12676 26188 12682 26240
rect 12728 26228 12756 26268
rect 15838 26256 15844 26268
rect 15896 26256 15902 26308
rect 16022 26256 16028 26308
rect 16080 26296 16086 26308
rect 16574 26296 16602 26336
rect 16853 26333 16865 26336
rect 16899 26333 16911 26367
rect 16853 26327 16911 26333
rect 17678 26324 17684 26376
rect 17736 26324 17742 26376
rect 17948 26367 18006 26373
rect 17948 26333 17960 26367
rect 17994 26364 18006 26367
rect 19426 26364 19432 26376
rect 17994 26336 19432 26364
rect 17994 26333 18006 26336
rect 17948 26327 18006 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 22066 26364 22094 26404
rect 22925 26367 22983 26373
rect 22925 26364 22937 26367
rect 22066 26336 22937 26364
rect 22925 26333 22937 26336
rect 22971 26333 22983 26367
rect 22925 26327 22983 26333
rect 23474 26324 23480 26376
rect 23532 26324 23538 26376
rect 23566 26324 23572 26376
rect 23624 26364 23630 26376
rect 23860 26373 23888 26404
rect 23661 26367 23719 26373
rect 23661 26364 23673 26367
rect 23624 26336 23673 26364
rect 23624 26324 23630 26336
rect 23661 26333 23673 26336
rect 23707 26333 23719 26367
rect 23661 26327 23719 26333
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26333 23903 26367
rect 23845 26327 23903 26333
rect 16080 26268 16602 26296
rect 16761 26299 16819 26305
rect 16080 26256 16086 26268
rect 16761 26265 16773 26299
rect 16807 26296 16819 26299
rect 24213 26299 24271 26305
rect 16807 26268 18000 26296
rect 16807 26265 16819 26268
rect 16761 26259 16819 26265
rect 17972 26240 18000 26268
rect 24213 26265 24225 26299
rect 24259 26296 24271 26299
rect 25130 26296 25136 26308
rect 24259 26268 25136 26296
rect 24259 26265 24271 26268
rect 24213 26259 24271 26265
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 16850 26228 16856 26240
rect 12728 26200 16856 26228
rect 16850 26188 16856 26200
rect 16908 26188 16914 26240
rect 17954 26188 17960 26240
rect 18012 26188 18018 26240
rect 19242 26188 19248 26240
rect 19300 26188 19306 26240
rect 23658 26188 23664 26240
rect 23716 26188 23722 26240
rect 1104 26138 25000 26160
rect 1104 26086 6884 26138
rect 6936 26086 6948 26138
rect 7000 26086 7012 26138
rect 7064 26086 7076 26138
rect 7128 26086 7140 26138
rect 7192 26086 12818 26138
rect 12870 26086 12882 26138
rect 12934 26086 12946 26138
rect 12998 26086 13010 26138
rect 13062 26086 13074 26138
rect 13126 26086 18752 26138
rect 18804 26086 18816 26138
rect 18868 26086 18880 26138
rect 18932 26086 18944 26138
rect 18996 26086 19008 26138
rect 19060 26086 24686 26138
rect 24738 26086 24750 26138
rect 24802 26086 24814 26138
rect 24866 26086 24878 26138
rect 24930 26086 24942 26138
rect 24994 26086 25000 26138
rect 1104 26064 25000 26086
rect 1670 25984 1676 26036
rect 1728 26024 1734 26036
rect 2590 26024 2596 26036
rect 1728 25996 2596 26024
rect 1728 25984 1734 25996
rect 2590 25984 2596 25996
rect 2648 25984 2654 26036
rect 3053 26027 3111 26033
rect 3053 25993 3065 26027
rect 3099 26024 3111 26027
rect 3329 26027 3387 26033
rect 3099 25996 3280 26024
rect 3099 25993 3111 25996
rect 3053 25987 3111 25993
rect 1302 25916 1308 25968
rect 1360 25956 1366 25968
rect 3252 25956 3280 25996
rect 3329 25993 3341 26027
rect 3375 26024 3387 26027
rect 7834 26024 7840 26036
rect 3375 25996 7840 26024
rect 3375 25993 3387 25996
rect 3329 25987 3387 25993
rect 7834 25984 7840 25996
rect 7892 25984 7898 26036
rect 8205 26027 8263 26033
rect 8205 25993 8217 26027
rect 8251 25993 8263 26027
rect 8205 25987 8263 25993
rect 3970 25956 3976 25968
rect 1360 25928 3188 25956
rect 3252 25928 3976 25956
rect 1360 25916 1366 25928
rect 1026 25848 1032 25900
rect 1084 25888 1090 25900
rect 1486 25888 1492 25900
rect 1084 25860 1492 25888
rect 1084 25848 1090 25860
rect 1486 25848 1492 25860
rect 1544 25848 1550 25900
rect 1762 25888 1768 25900
rect 1723 25860 1768 25888
rect 1762 25848 1768 25860
rect 1820 25848 1826 25900
rect 1854 25848 1860 25900
rect 1912 25888 1918 25900
rect 2682 25888 2688 25900
rect 1912 25860 2688 25888
rect 1912 25848 1918 25860
rect 2682 25848 2688 25860
rect 2740 25848 2746 25900
rect 3160 25897 3188 25928
rect 3970 25916 3976 25928
rect 4028 25916 4034 25968
rect 5350 25956 5356 25968
rect 4816 25928 5356 25956
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25857 2927 25891
rect 2869 25851 2927 25857
rect 3145 25891 3203 25897
rect 3145 25857 3157 25891
rect 3191 25857 3203 25891
rect 3145 25851 3203 25857
rect 2222 25712 2228 25764
rect 2280 25752 2286 25764
rect 2884 25752 2912 25851
rect 3326 25848 3332 25900
rect 3384 25888 3390 25900
rect 3421 25891 3479 25897
rect 3421 25888 3433 25891
rect 3384 25860 3433 25888
rect 3384 25848 3390 25860
rect 3421 25857 3433 25860
rect 3467 25857 3479 25891
rect 3421 25851 3479 25857
rect 3695 25891 3753 25897
rect 3695 25857 3707 25891
rect 3741 25888 3753 25891
rect 4430 25888 4436 25900
rect 3741 25860 4436 25888
rect 3741 25857 3753 25860
rect 3695 25851 3753 25857
rect 4430 25848 4436 25860
rect 4488 25888 4494 25900
rect 4816 25897 4844 25928
rect 5350 25916 5356 25928
rect 5408 25916 5414 25968
rect 5994 25956 6000 25968
rect 5460 25928 6000 25956
rect 4801 25891 4859 25897
rect 4488 25860 4568 25888
rect 4488 25848 4494 25860
rect 2280 25724 2912 25752
rect 4540 25752 4568 25860
rect 4801 25857 4813 25891
rect 4847 25857 4859 25891
rect 4801 25851 4859 25857
rect 5075 25891 5133 25897
rect 5075 25857 5087 25891
rect 5121 25888 5133 25891
rect 5460 25888 5488 25928
rect 5994 25916 6000 25928
rect 6052 25916 6058 25968
rect 6840 25928 7052 25956
rect 6840 25897 6868 25928
rect 5121 25860 5488 25888
rect 6825 25891 6883 25897
rect 5121 25857 5133 25860
rect 5075 25851 5133 25857
rect 6825 25857 6837 25891
rect 6871 25857 6883 25891
rect 7024 25888 7052 25928
rect 7098 25916 7104 25968
rect 7156 25916 7162 25968
rect 7282 25916 7288 25968
rect 7340 25956 7346 25968
rect 7340 25928 7880 25956
rect 7340 25916 7346 25928
rect 7377 25891 7435 25897
rect 7377 25888 7389 25891
rect 7024 25860 7389 25888
rect 6825 25851 6883 25857
rect 7377 25857 7389 25860
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25888 7527 25891
rect 7650 25888 7656 25900
rect 7515 25860 7656 25888
rect 7515 25857 7527 25860
rect 7469 25851 7527 25857
rect 7650 25848 7656 25860
rect 7708 25848 7714 25900
rect 7852 25897 7880 25928
rect 8220 25900 8248 25987
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10744 25996 10885 26024
rect 10744 25984 10750 25996
rect 10873 25993 10885 25996
rect 10919 25993 10931 26027
rect 10873 25987 10931 25993
rect 11146 25984 11152 26036
rect 11204 26024 11210 26036
rect 12250 26024 12256 26036
rect 11204 25996 12256 26024
rect 11204 25984 11210 25996
rect 12250 25984 12256 25996
rect 12308 25984 12314 26036
rect 12526 25984 12532 26036
rect 12584 26024 12590 26036
rect 13446 26024 13452 26036
rect 12584 25996 13452 26024
rect 12584 25984 12590 25996
rect 13446 25984 13452 25996
rect 13504 25984 13510 26036
rect 15010 25984 15016 26036
rect 15068 25984 15074 26036
rect 15654 25984 15660 26036
rect 15712 25984 15718 26036
rect 15930 25984 15936 26036
rect 15988 25984 15994 26036
rect 16022 25984 16028 26036
rect 16080 25984 16086 26036
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 17218 26024 17224 26036
rect 16540 25996 17224 26024
rect 16540 25984 16546 25996
rect 17218 25984 17224 25996
rect 17276 25984 17282 26036
rect 19978 26024 19984 26036
rect 18524 25996 19984 26024
rect 11882 25956 11888 25968
rect 11808 25928 11888 25956
rect 11808 25927 11836 25928
rect 11775 25921 11836 25927
rect 7837 25891 7895 25897
rect 7837 25857 7849 25891
rect 7883 25857 7895 25891
rect 7837 25851 7895 25857
rect 8202 25848 8208 25900
rect 8260 25848 8266 25900
rect 10042 25848 10048 25900
rect 10100 25897 10106 25900
rect 10100 25891 10128 25897
rect 10116 25857 10128 25891
rect 10100 25851 10128 25857
rect 10100 25848 10106 25851
rect 11514 25848 11520 25900
rect 11572 25848 11578 25900
rect 11775 25887 11787 25921
rect 11821 25890 11836 25921
rect 11882 25916 11888 25928
rect 11940 25916 11946 25968
rect 15028 25956 15056 25984
rect 15028 25928 15608 25956
rect 11821 25887 11833 25890
rect 11775 25881 11833 25887
rect 13262 25848 13268 25900
rect 13320 25848 13326 25900
rect 14274 25848 14280 25900
rect 14332 25848 14338 25900
rect 15580 25897 15608 25928
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25888 14979 25891
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 14967 25860 15485 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 15565 25891 15623 25897
rect 15565 25857 15577 25891
rect 15611 25857 15623 25891
rect 15565 25851 15623 25857
rect 15841 25891 15899 25897
rect 15841 25857 15853 25891
rect 15887 25888 15899 25891
rect 15948 25888 15976 25984
rect 15887 25860 15976 25888
rect 16025 25891 16083 25897
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16025 25857 16037 25891
rect 16071 25857 16083 25891
rect 18524 25888 18552 25996
rect 19978 25984 19984 25996
rect 20036 25984 20042 26036
rect 22373 26027 22431 26033
rect 22373 25993 22385 26027
rect 22419 25993 22431 26027
rect 22373 25987 22431 25993
rect 23477 26027 23535 26033
rect 23477 25993 23489 26027
rect 23523 26024 23535 26027
rect 23566 26024 23572 26036
rect 23523 25996 23572 26024
rect 23523 25993 23535 25996
rect 23477 25987 23535 25993
rect 18690 25916 18696 25968
rect 18748 25956 18754 25968
rect 22388 25956 22416 25987
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 23937 26027 23995 26033
rect 23937 25993 23949 26027
rect 23983 26024 23995 26027
rect 24026 26024 24032 26036
rect 23983 25996 24032 26024
rect 23983 25993 23995 25996
rect 23937 25987 23995 25993
rect 24026 25984 24032 25996
rect 24084 25984 24090 26036
rect 18748 25928 18886 25956
rect 22388 25928 23060 25956
rect 18748 25916 18754 25928
rect 18858 25927 18886 25928
rect 18858 25921 18917 25927
rect 18601 25891 18659 25897
rect 18601 25888 18613 25891
rect 18524 25860 18613 25888
rect 16025 25851 16083 25857
rect 18601 25857 18613 25860
rect 18647 25857 18659 25891
rect 18858 25890 18871 25921
rect 18859 25887 18871 25890
rect 18905 25887 18917 25921
rect 19981 25891 20039 25897
rect 19981 25888 19993 25891
rect 18859 25881 18917 25887
rect 18601 25851 18659 25857
rect 19628 25860 19993 25888
rect 7558 25780 7564 25832
rect 7616 25780 7622 25832
rect 8294 25780 8300 25832
rect 8352 25820 8358 25832
rect 9033 25823 9091 25829
rect 9033 25820 9045 25823
rect 8352 25792 9045 25820
rect 8352 25780 8358 25792
rect 9033 25789 9045 25792
rect 9079 25789 9091 25823
rect 9033 25783 9091 25789
rect 9214 25780 9220 25832
rect 9272 25780 9278 25832
rect 9953 25823 10011 25829
rect 9953 25820 9965 25823
rect 9600 25792 9965 25820
rect 9600 25764 9628 25792
rect 9953 25789 9965 25792
rect 9999 25789 10011 25823
rect 9953 25783 10011 25789
rect 10229 25823 10287 25829
rect 10229 25789 10241 25823
rect 10275 25820 10287 25823
rect 10410 25820 10416 25832
rect 10275 25792 10416 25820
rect 10275 25789 10287 25792
rect 10229 25783 10287 25789
rect 10410 25780 10416 25792
rect 10468 25780 10474 25832
rect 12342 25780 12348 25832
rect 12400 25820 12406 25832
rect 13081 25823 13139 25829
rect 13081 25820 13093 25823
rect 12400 25792 13093 25820
rect 12400 25780 12406 25792
rect 13081 25789 13093 25792
rect 13127 25820 13139 25823
rect 13127 25792 13308 25820
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 4540 25724 4936 25752
rect 2280 25712 2286 25724
rect 4908 25696 4936 25724
rect 9582 25712 9588 25764
rect 9640 25712 9646 25764
rect 9674 25712 9680 25764
rect 9732 25712 9738 25764
rect 13280 25696 13308 25792
rect 13722 25780 13728 25832
rect 13780 25780 13786 25832
rect 13998 25780 14004 25832
rect 14056 25780 14062 25832
rect 14090 25780 14096 25832
rect 14148 25829 14154 25832
rect 14148 25823 14176 25829
rect 14164 25789 14176 25823
rect 16040 25820 16068 25851
rect 14148 25783 14176 25789
rect 15304 25792 16068 25820
rect 14148 25780 14154 25783
rect 15304 25761 15332 25792
rect 19628 25761 19656 25860
rect 19981 25857 19993 25860
rect 20027 25888 20039 25891
rect 20349 25891 20407 25897
rect 20349 25888 20361 25891
rect 20027 25860 20361 25888
rect 20027 25857 20039 25860
rect 19981 25851 20039 25857
rect 20349 25857 20361 25860
rect 20395 25857 20407 25891
rect 20349 25851 20407 25857
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25888 20591 25891
rect 20622 25888 20628 25900
rect 20579 25860 20628 25888
rect 20579 25857 20591 25860
rect 20533 25851 20591 25857
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 21358 25848 21364 25900
rect 21416 25848 21422 25900
rect 21542 25848 21548 25900
rect 21600 25848 21606 25900
rect 23032 25897 23060 25928
rect 24118 25916 24124 25968
rect 24176 25916 24182 25968
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 22112 25860 22569 25888
rect 22112 25832 22140 25860
rect 22557 25857 22569 25860
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25857 23075 25891
rect 23017 25851 23075 25857
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 23624 25860 23673 25888
rect 23624 25848 23630 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 23753 25891 23811 25897
rect 23753 25857 23765 25891
rect 23799 25857 23811 25891
rect 23753 25851 23811 25857
rect 20257 25823 20315 25829
rect 20257 25789 20269 25823
rect 20303 25820 20315 25823
rect 20441 25823 20499 25829
rect 20441 25820 20453 25823
rect 20303 25792 20453 25820
rect 20303 25789 20315 25792
rect 20257 25783 20315 25789
rect 20441 25789 20453 25792
rect 20487 25789 20499 25823
rect 20441 25783 20499 25789
rect 22094 25780 22100 25832
rect 22152 25780 22158 25832
rect 23382 25780 23388 25832
rect 23440 25820 23446 25832
rect 23768 25820 23796 25851
rect 23440 25792 23796 25820
rect 23440 25780 23446 25792
rect 15289 25755 15347 25761
rect 15289 25721 15301 25755
rect 15335 25721 15347 25755
rect 15289 25715 15347 25721
rect 19613 25755 19671 25761
rect 19613 25721 19625 25755
rect 19659 25721 19671 25755
rect 19613 25715 19671 25721
rect 20165 25755 20223 25761
rect 20165 25721 20177 25755
rect 20211 25752 20223 25755
rect 23934 25752 23940 25764
rect 20211 25724 23940 25752
rect 20211 25721 20223 25724
rect 20165 25715 20223 25721
rect 23934 25712 23940 25724
rect 23992 25712 23998 25764
rect 1946 25644 1952 25696
rect 2004 25684 2010 25696
rect 2501 25687 2559 25693
rect 2501 25684 2513 25687
rect 2004 25656 2513 25684
rect 2004 25644 2010 25656
rect 2501 25653 2513 25656
rect 2547 25653 2559 25687
rect 2501 25647 2559 25653
rect 2590 25644 2596 25696
rect 2648 25684 2654 25696
rect 3050 25684 3056 25696
rect 2648 25656 3056 25684
rect 2648 25644 2654 25656
rect 3050 25644 3056 25656
rect 3108 25644 3114 25696
rect 3326 25644 3332 25696
rect 3384 25684 3390 25696
rect 4246 25684 4252 25696
rect 3384 25656 4252 25684
rect 3384 25644 3390 25656
rect 4246 25644 4252 25656
rect 4304 25644 4310 25696
rect 4430 25644 4436 25696
rect 4488 25644 4494 25696
rect 4890 25644 4896 25696
rect 4948 25644 4954 25696
rect 5810 25644 5816 25696
rect 5868 25644 5874 25696
rect 6086 25644 6092 25696
rect 6144 25684 6150 25696
rect 7098 25684 7104 25696
rect 6144 25656 7104 25684
rect 6144 25644 6150 25656
rect 7098 25644 7104 25656
rect 7156 25644 7162 25696
rect 8389 25687 8447 25693
rect 8389 25653 8401 25687
rect 8435 25684 8447 25687
rect 12342 25684 12348 25696
rect 8435 25656 12348 25684
rect 8435 25653 8447 25656
rect 8389 25647 8447 25653
rect 12342 25644 12348 25656
rect 12400 25644 12406 25696
rect 12526 25644 12532 25696
rect 12584 25644 12590 25696
rect 13262 25644 13268 25696
rect 13320 25644 13326 25696
rect 20070 25644 20076 25696
rect 20128 25644 20134 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 23106 25644 23112 25696
rect 23164 25644 23170 25696
rect 24394 25644 24400 25696
rect 24452 25644 24458 25696
rect 1104 25594 24840 25616
rect 1104 25542 3917 25594
rect 3969 25542 3981 25594
rect 4033 25542 4045 25594
rect 4097 25542 4109 25594
rect 4161 25542 4173 25594
rect 4225 25542 9851 25594
rect 9903 25542 9915 25594
rect 9967 25542 9979 25594
rect 10031 25542 10043 25594
rect 10095 25542 10107 25594
rect 10159 25542 15785 25594
rect 15837 25542 15849 25594
rect 15901 25542 15913 25594
rect 15965 25542 15977 25594
rect 16029 25542 16041 25594
rect 16093 25542 21719 25594
rect 21771 25542 21783 25594
rect 21835 25542 21847 25594
rect 21899 25542 21911 25594
rect 21963 25542 21975 25594
rect 22027 25542 24840 25594
rect 1104 25520 24840 25542
rect 1210 25440 1216 25492
rect 1268 25480 1274 25492
rect 2222 25480 2228 25492
rect 1268 25452 2228 25480
rect 1268 25440 1274 25452
rect 2222 25440 2228 25452
rect 2280 25440 2286 25492
rect 3234 25480 3240 25492
rect 2332 25452 3240 25480
rect 1581 25415 1639 25421
rect 1581 25381 1593 25415
rect 1627 25412 1639 25415
rect 2130 25412 2136 25424
rect 1627 25384 2136 25412
rect 1627 25381 1639 25384
rect 1581 25375 1639 25381
rect 2130 25372 2136 25384
rect 2188 25372 2194 25424
rect 2332 25353 2360 25452
rect 3234 25440 3240 25452
rect 3292 25440 3298 25492
rect 5442 25440 5448 25492
rect 5500 25440 5506 25492
rect 7742 25440 7748 25492
rect 7800 25480 7806 25492
rect 8297 25483 8355 25489
rect 8297 25480 8309 25483
rect 7800 25452 8309 25480
rect 7800 25440 7806 25452
rect 8297 25449 8309 25452
rect 8343 25449 8355 25483
rect 8297 25443 8355 25449
rect 8478 25440 8484 25492
rect 8536 25480 8542 25492
rect 8846 25480 8852 25492
rect 8536 25452 8852 25480
rect 8536 25440 8542 25452
rect 8846 25440 8852 25452
rect 8904 25480 8910 25492
rect 8904 25452 10364 25480
rect 8904 25440 8910 25452
rect 3329 25415 3387 25421
rect 3329 25381 3341 25415
rect 3375 25412 3387 25415
rect 3375 25384 3832 25412
rect 3375 25381 3387 25384
rect 3329 25375 3387 25381
rect 2317 25347 2375 25353
rect 2317 25313 2329 25347
rect 2363 25313 2375 25347
rect 3804 25330 3832 25384
rect 5460 25344 5488 25440
rect 2317 25307 2375 25313
rect 5092 25316 5488 25344
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 1670 25236 1676 25288
rect 1728 25236 1734 25288
rect 2130 25236 2136 25288
rect 2188 25236 2194 25288
rect 2591 25279 2649 25285
rect 2591 25245 2603 25279
rect 2637 25276 2649 25279
rect 2682 25276 2688 25288
rect 2637 25248 2688 25276
rect 2637 25245 2649 25248
rect 2591 25239 2649 25245
rect 2682 25236 2688 25248
rect 2740 25276 2746 25288
rect 4062 25276 4068 25288
rect 2740 25248 4068 25276
rect 2740 25236 2746 25248
rect 4062 25236 4068 25248
rect 4120 25236 4126 25288
rect 4341 25279 4399 25285
rect 4341 25245 4353 25279
rect 4387 25276 4399 25279
rect 4430 25276 4436 25288
rect 4387 25248 4436 25276
rect 4387 25245 4399 25248
rect 4341 25239 4399 25245
rect 4430 25236 4436 25248
rect 4488 25236 4494 25288
rect 4522 25236 4528 25288
rect 4580 25276 4586 25288
rect 5092 25276 5120 25316
rect 6546 25304 6552 25356
rect 6604 25344 6610 25356
rect 7282 25344 7288 25356
rect 6604 25316 7288 25344
rect 6604 25304 6610 25316
rect 7282 25304 7288 25316
rect 7340 25304 7346 25356
rect 8846 25304 8852 25356
rect 8904 25344 8910 25356
rect 9398 25344 9404 25356
rect 8904 25316 9404 25344
rect 8904 25304 8910 25316
rect 9398 25304 9404 25316
rect 9456 25344 9462 25356
rect 9493 25347 9551 25353
rect 9493 25344 9505 25347
rect 9456 25316 9505 25344
rect 9456 25304 9462 25316
rect 9493 25313 9505 25316
rect 9539 25313 9551 25347
rect 10336 25344 10364 25452
rect 10410 25440 10416 25492
rect 10468 25480 10474 25492
rect 10505 25483 10563 25489
rect 10505 25480 10517 25483
rect 10468 25452 10517 25480
rect 10468 25440 10474 25452
rect 10505 25449 10517 25452
rect 10551 25449 10563 25483
rect 18230 25480 18236 25492
rect 10505 25443 10563 25449
rect 17420 25452 18236 25480
rect 12713 25415 12771 25421
rect 12713 25381 12725 25415
rect 12759 25412 12771 25415
rect 17420 25412 17448 25452
rect 18230 25440 18236 25452
rect 18288 25440 18294 25492
rect 19337 25483 19395 25489
rect 19337 25449 19349 25483
rect 19383 25480 19395 25483
rect 20070 25480 20076 25492
rect 19383 25452 20076 25480
rect 19383 25449 19395 25452
rect 19337 25443 19395 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20622 25480 20628 25492
rect 20180 25452 20628 25480
rect 12759 25384 17448 25412
rect 12759 25381 12771 25384
rect 12713 25375 12771 25381
rect 19518 25372 19524 25424
rect 19576 25372 19582 25424
rect 19613 25415 19671 25421
rect 19613 25381 19625 25415
rect 19659 25412 19671 25415
rect 20180 25412 20208 25452
rect 20622 25440 20628 25452
rect 20680 25440 20686 25492
rect 21358 25440 21364 25492
rect 21416 25440 21422 25492
rect 23106 25440 23112 25492
rect 23164 25480 23170 25492
rect 23477 25483 23535 25489
rect 23477 25480 23489 25483
rect 23164 25452 23489 25480
rect 23164 25440 23170 25452
rect 23477 25449 23489 25452
rect 23523 25449 23535 25483
rect 23477 25443 23535 25449
rect 23566 25440 23572 25492
rect 23624 25440 23630 25492
rect 23658 25440 23664 25492
rect 23716 25440 23722 25492
rect 19659 25384 20208 25412
rect 23201 25415 23259 25421
rect 19659 25381 19671 25384
rect 19613 25375 19671 25381
rect 23201 25381 23213 25415
rect 23247 25412 23259 25415
rect 23584 25412 23612 25440
rect 23247 25384 23612 25412
rect 23247 25381 23259 25384
rect 23201 25375 23259 25381
rect 12526 25344 12532 25356
rect 10336 25316 11008 25344
rect 12466 25316 12532 25344
rect 9493 25307 9551 25313
rect 4580 25248 5120 25276
rect 4580 25236 4586 25248
rect 4249 25211 4307 25217
rect 2746 25180 4200 25208
rect 1854 25100 1860 25152
rect 1912 25100 1918 25152
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 2746 25140 2774 25180
rect 4172 25152 4200 25180
rect 4249 25177 4261 25211
rect 4295 25208 4307 25211
rect 4614 25208 4620 25220
rect 4295 25180 4620 25208
rect 4295 25177 4307 25180
rect 4249 25171 4307 25177
rect 4614 25168 4620 25180
rect 4672 25168 4678 25220
rect 5092 25217 5120 25248
rect 5442 25236 5448 25288
rect 5500 25236 5506 25288
rect 5703 25249 5761 25255
rect 4709 25211 4767 25217
rect 4709 25177 4721 25211
rect 4755 25177 4767 25211
rect 4709 25171 4767 25177
rect 5077 25211 5135 25217
rect 5077 25177 5089 25211
rect 5123 25177 5135 25211
rect 5703 25215 5715 25249
rect 5749 25246 5761 25249
rect 5749 25215 5764 25246
rect 6914 25236 6920 25288
rect 6972 25276 6978 25288
rect 7558 25276 7564 25288
rect 6972 25248 7564 25276
rect 6972 25236 6978 25248
rect 7558 25236 7564 25248
rect 7616 25236 7622 25288
rect 9767 25279 9825 25285
rect 9767 25245 9779 25279
rect 9813 25276 9825 25279
rect 10870 25276 10876 25288
rect 9813 25248 10876 25276
rect 9813 25245 9825 25248
rect 9767 25239 9825 25245
rect 10870 25236 10876 25248
rect 10928 25236 10934 25288
rect 5703 25209 5764 25215
rect 5736 25208 5764 25209
rect 5736 25180 8156 25208
rect 5077 25171 5135 25177
rect 1995 25112 2774 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 3510 25100 3516 25152
rect 3568 25140 3574 25152
rect 3786 25140 3792 25152
rect 3568 25112 3792 25140
rect 3568 25100 3574 25112
rect 3786 25100 3792 25112
rect 3844 25140 3850 25152
rect 3970 25140 3976 25152
rect 3844 25112 3976 25140
rect 3844 25100 3850 25112
rect 3970 25100 3976 25112
rect 4028 25100 4034 25152
rect 4154 25100 4160 25152
rect 4212 25140 4218 25152
rect 4724 25140 4752 25171
rect 8128 25152 8156 25180
rect 8662 25168 8668 25220
rect 8720 25208 8726 25220
rect 9030 25208 9036 25220
rect 8720 25180 9036 25208
rect 8720 25168 8726 25180
rect 9030 25168 9036 25180
rect 9088 25168 9094 25220
rect 9582 25168 9588 25220
rect 9640 25208 9646 25220
rect 10134 25208 10140 25220
rect 9640 25180 10140 25208
rect 9640 25168 9646 25180
rect 10134 25168 10140 25180
rect 10192 25168 10198 25220
rect 10980 25208 11008 25316
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 15378 25304 15384 25356
rect 15436 25304 15442 25356
rect 16669 25347 16727 25353
rect 16669 25313 16681 25347
rect 16715 25344 16727 25347
rect 16758 25344 16764 25356
rect 16715 25316 16764 25344
rect 16715 25313 16727 25316
rect 16669 25307 16727 25313
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 17310 25304 17316 25356
rect 17368 25304 17374 25356
rect 17402 25304 17408 25356
rect 17460 25344 17466 25356
rect 17706 25347 17764 25353
rect 17706 25344 17718 25347
rect 17460 25316 17718 25344
rect 17460 25304 17466 25316
rect 17706 25313 17718 25316
rect 17752 25313 17764 25347
rect 17706 25307 17764 25313
rect 17865 25347 17923 25353
rect 17865 25313 17877 25347
rect 17911 25344 17923 25347
rect 18506 25344 18512 25356
rect 17911 25316 18512 25344
rect 17911 25313 17923 25316
rect 17865 25307 17923 25313
rect 18506 25304 18512 25316
rect 18564 25304 18570 25356
rect 11808 25248 12296 25276
rect 11425 25211 11483 25217
rect 11425 25208 11437 25211
rect 10980 25180 11437 25208
rect 11425 25177 11437 25180
rect 11471 25177 11483 25211
rect 11425 25171 11483 25177
rect 11698 25168 11704 25220
rect 11756 25168 11762 25220
rect 11808 25217 11836 25248
rect 11793 25211 11851 25217
rect 11793 25177 11805 25211
rect 11839 25177 11851 25211
rect 11793 25171 11851 25177
rect 12161 25211 12219 25217
rect 12161 25177 12173 25211
rect 12207 25177 12219 25211
rect 12268 25208 12296 25248
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 15396 25276 15424 25304
rect 16853 25279 16911 25285
rect 16853 25276 16865 25279
rect 12400 25248 15332 25276
rect 15396 25248 16865 25276
rect 12400 25236 12406 25248
rect 12434 25208 12440 25220
rect 12268 25180 12440 25208
rect 12161 25171 12219 25177
rect 4212 25112 4752 25140
rect 5261 25143 5319 25149
rect 4212 25100 4218 25112
rect 5261 25109 5273 25143
rect 5307 25140 5319 25143
rect 6086 25140 6092 25152
rect 5307 25112 6092 25140
rect 5307 25109 5319 25112
rect 5261 25103 5319 25109
rect 6086 25100 6092 25112
rect 6144 25100 6150 25152
rect 6362 25100 6368 25152
rect 6420 25140 6426 25152
rect 6457 25143 6515 25149
rect 6457 25140 6469 25143
rect 6420 25112 6469 25140
rect 6420 25100 6426 25112
rect 6457 25109 6469 25112
rect 6503 25109 6515 25143
rect 6457 25103 6515 25109
rect 8110 25100 8116 25152
rect 8168 25140 8174 25152
rect 11514 25140 11520 25152
rect 8168 25112 11520 25140
rect 8168 25100 8174 25112
rect 11514 25100 11520 25112
rect 11572 25100 11578 25152
rect 11716 25140 11744 25168
rect 12066 25140 12072 25152
rect 11716 25112 12072 25140
rect 12066 25100 12072 25112
rect 12124 25100 12130 25152
rect 12176 25140 12204 25171
rect 12434 25168 12440 25180
rect 12492 25168 12498 25220
rect 12529 25211 12587 25217
rect 12529 25177 12541 25211
rect 12575 25208 12587 25211
rect 12618 25208 12624 25220
rect 12575 25180 12624 25208
rect 12575 25177 12587 25180
rect 12529 25171 12587 25177
rect 12250 25140 12256 25152
rect 12176 25112 12256 25140
rect 12250 25100 12256 25112
rect 12308 25100 12314 25152
rect 12342 25100 12348 25152
rect 12400 25140 12406 25152
rect 12544 25140 12572 25171
rect 12618 25168 12624 25180
rect 12676 25168 12682 25220
rect 12400 25112 12572 25140
rect 15304 25140 15332 25248
rect 16684 25220 16712 25248
rect 16853 25245 16865 25248
rect 16899 25245 16911 25279
rect 16853 25239 16911 25245
rect 17586 25236 17592 25288
rect 17644 25236 17650 25288
rect 19242 25236 19248 25288
rect 19300 25236 19306 25288
rect 19536 25276 19564 25372
rect 19702 25304 19708 25356
rect 19760 25344 19766 25356
rect 19978 25344 19984 25356
rect 19760 25316 19984 25344
rect 19760 25304 19766 25316
rect 19978 25304 19984 25316
rect 20036 25344 20042 25356
rect 20349 25347 20407 25353
rect 20349 25344 20361 25347
rect 20036 25316 20361 25344
rect 20036 25304 20042 25316
rect 20349 25313 20361 25316
rect 20395 25313 20407 25347
rect 20349 25307 20407 25313
rect 21174 25304 21180 25356
rect 21232 25344 21238 25356
rect 21821 25347 21879 25353
rect 21821 25344 21833 25347
rect 21232 25316 21833 25344
rect 21232 25304 21238 25316
rect 21821 25313 21833 25316
rect 21867 25313 21879 25347
rect 21821 25307 21879 25313
rect 23474 25304 23480 25356
rect 23532 25304 23538 25356
rect 23676 25353 23704 25440
rect 23661 25347 23719 25353
rect 23661 25313 23673 25347
rect 23707 25313 23719 25347
rect 23661 25307 23719 25313
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19536 25248 19809 25276
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 20622 25276 20628 25288
rect 20583 25248 20628 25276
rect 19797 25239 19855 25245
rect 20622 25236 20628 25248
rect 20680 25236 20686 25288
rect 22554 25236 22560 25288
rect 22612 25236 22618 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25276 23443 25279
rect 23492 25276 23520 25304
rect 23431 25248 23520 25276
rect 23431 25245 23443 25248
rect 23385 25239 23443 25245
rect 16666 25168 16672 25220
rect 16724 25168 16730 25220
rect 22094 25217 22100 25220
rect 18340 25180 21220 25208
rect 18340 25140 18368 25180
rect 21192 25152 21220 25180
rect 22088 25171 22100 25217
rect 22152 25208 22158 25220
rect 22572 25208 22600 25236
rect 23845 25211 23903 25217
rect 23845 25208 23857 25211
rect 22152 25180 22188 25208
rect 22572 25180 23857 25208
rect 22094 25168 22100 25171
rect 22152 25168 22158 25180
rect 23845 25177 23857 25180
rect 23891 25177 23903 25211
rect 23845 25171 23903 25177
rect 24213 25211 24271 25217
rect 24213 25177 24225 25211
rect 24259 25208 24271 25211
rect 25130 25208 25136 25220
rect 24259 25180 25136 25208
rect 24259 25177 24271 25180
rect 24213 25171 24271 25177
rect 25130 25168 25136 25180
rect 25188 25168 25194 25220
rect 15304 25112 18368 25140
rect 18509 25143 18567 25149
rect 12400 25100 12406 25112
rect 18509 25109 18521 25143
rect 18555 25140 18567 25143
rect 19242 25140 19248 25152
rect 18555 25112 19248 25140
rect 18555 25109 18567 25112
rect 18509 25103 18567 25109
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 21174 25100 21180 25152
rect 21232 25100 21238 25152
rect 23661 25143 23719 25149
rect 23661 25109 23673 25143
rect 23707 25140 23719 25143
rect 23750 25140 23756 25152
rect 23707 25112 23756 25140
rect 23707 25109 23719 25112
rect 23661 25103 23719 25109
rect 23750 25100 23756 25112
rect 23808 25100 23814 25152
rect 1104 25050 25000 25072
rect 1104 24998 6884 25050
rect 6936 24998 6948 25050
rect 7000 24998 7012 25050
rect 7064 24998 7076 25050
rect 7128 24998 7140 25050
rect 7192 24998 12818 25050
rect 12870 24998 12882 25050
rect 12934 24998 12946 25050
rect 12998 24998 13010 25050
rect 13062 24998 13074 25050
rect 13126 24998 18752 25050
rect 18804 24998 18816 25050
rect 18868 24998 18880 25050
rect 18932 24998 18944 25050
rect 18996 24998 19008 25050
rect 19060 24998 24686 25050
rect 24738 24998 24750 25050
rect 24802 24998 24814 25050
rect 24866 24998 24878 25050
rect 24930 24998 24942 25050
rect 24994 24998 25000 25050
rect 1104 24976 25000 24998
rect 1857 24939 1915 24945
rect 1857 24905 1869 24939
rect 1903 24905 1915 24939
rect 1857 24899 1915 24905
rect 1302 24828 1308 24880
rect 1360 24868 1366 24880
rect 1872 24868 1900 24899
rect 2038 24896 2044 24948
rect 2096 24936 2102 24948
rect 2133 24939 2191 24945
rect 2133 24936 2145 24939
rect 2096 24908 2145 24936
rect 2096 24896 2102 24908
rect 2133 24905 2145 24908
rect 2179 24905 2191 24939
rect 2133 24899 2191 24905
rect 2869 24939 2927 24945
rect 2869 24905 2881 24939
rect 2915 24936 2927 24939
rect 2958 24936 2964 24948
rect 2915 24908 2964 24936
rect 2915 24905 2927 24908
rect 2869 24899 2927 24905
rect 2958 24896 2964 24908
rect 3016 24896 3022 24948
rect 3050 24896 3056 24948
rect 3108 24936 3114 24948
rect 3987 24939 4045 24945
rect 3108 24908 3924 24936
rect 3108 24896 3114 24908
rect 1360 24840 1808 24868
rect 1872 24840 3464 24868
rect 1360 24828 1366 24840
rect 750 24760 756 24812
rect 808 24800 814 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 808 24772 1409 24800
rect 808 24760 814 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 1486 24760 1492 24812
rect 1544 24800 1550 24812
rect 1673 24803 1731 24809
rect 1673 24800 1685 24803
rect 1544 24772 1685 24800
rect 1544 24760 1550 24772
rect 1673 24769 1685 24772
rect 1719 24769 1731 24803
rect 1780 24800 1808 24840
rect 1949 24803 2007 24809
rect 1949 24800 1961 24803
rect 1780 24772 1961 24800
rect 1673 24763 1731 24769
rect 1949 24769 1961 24772
rect 1995 24769 2007 24803
rect 1949 24763 2007 24769
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24769 2283 24803
rect 2225 24763 2283 24769
rect 1118 24692 1124 24744
rect 1176 24732 1182 24744
rect 2240 24732 2268 24763
rect 2774 24760 2780 24812
rect 2832 24800 2838 24812
rect 3145 24803 3203 24809
rect 3145 24800 3157 24803
rect 2832 24772 3157 24800
rect 2832 24760 2838 24772
rect 3145 24769 3157 24772
rect 3191 24769 3203 24803
rect 3145 24763 3203 24769
rect 3234 24760 3240 24812
rect 3292 24760 3298 24812
rect 3436 24800 3464 24840
rect 3510 24828 3516 24880
rect 3568 24868 3574 24880
rect 3605 24871 3663 24877
rect 3605 24868 3617 24871
rect 3568 24840 3617 24868
rect 3568 24828 3574 24840
rect 3605 24837 3617 24840
rect 3651 24837 3663 24871
rect 3896 24868 3924 24908
rect 3987 24905 3999 24939
rect 4033 24936 4045 24939
rect 4154 24936 4160 24948
rect 4033 24908 4160 24936
rect 4033 24905 4045 24908
rect 3987 24899 4045 24905
rect 4154 24896 4160 24908
rect 4212 24896 4218 24948
rect 8202 24936 8208 24948
rect 4540 24908 8208 24936
rect 4540 24868 4568 24908
rect 8202 24896 8208 24908
rect 8260 24896 8266 24948
rect 8294 24896 8300 24948
rect 8352 24936 8358 24948
rect 12250 24936 12256 24948
rect 8352 24908 12256 24936
rect 8352 24896 8358 24908
rect 12250 24896 12256 24908
rect 12308 24896 12314 24948
rect 15010 24896 15016 24948
rect 15068 24936 15074 24948
rect 15068 24908 17172 24936
rect 15068 24896 15074 24908
rect 8846 24868 8852 24880
rect 3896 24840 4568 24868
rect 8496 24840 8852 24868
rect 3605 24831 3663 24837
rect 3786 24800 3792 24812
rect 3436 24772 3792 24800
rect 3786 24760 3792 24772
rect 3844 24760 3850 24812
rect 3970 24760 3976 24812
rect 4028 24800 4034 24812
rect 4341 24803 4399 24809
rect 4341 24800 4353 24803
rect 4028 24772 4353 24800
rect 4028 24760 4034 24772
rect 4341 24769 4353 24772
rect 4387 24769 4399 24803
rect 4341 24763 4399 24769
rect 4522 24760 4528 24812
rect 4580 24760 4586 24812
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 6454 24760 6460 24812
rect 6512 24800 6518 24812
rect 8018 24800 8024 24812
rect 6512 24772 8024 24800
rect 6512 24760 6518 24772
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 8496 24809 8524 24840
rect 8846 24828 8852 24840
rect 8904 24828 8910 24880
rect 9214 24828 9220 24880
rect 9272 24868 9278 24880
rect 12158 24868 12164 24880
rect 9272 24840 12164 24868
rect 9272 24828 9278 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 12710 24868 12716 24880
rect 12450 24840 12716 24868
rect 12450 24839 12478 24840
rect 12419 24833 12478 24839
rect 8481 24803 8539 24809
rect 8481 24769 8493 24803
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 8755 24803 8813 24809
rect 8755 24800 8767 24803
rect 8720 24772 8767 24800
rect 8720 24760 8726 24772
rect 8755 24769 8767 24772
rect 8801 24800 8813 24803
rect 11330 24800 11336 24812
rect 8801 24772 11336 24800
rect 8801 24769 8813 24772
rect 8755 24763 8813 24769
rect 11330 24760 11336 24772
rect 11388 24760 11394 24812
rect 11514 24760 11520 24812
rect 11572 24800 11578 24812
rect 12419 24800 12431 24833
rect 11572 24799 12431 24800
rect 12465 24799 12478 24833
rect 12710 24828 12716 24840
rect 12768 24828 12774 24880
rect 16758 24868 16764 24880
rect 16500 24840 16764 24868
rect 11572 24772 12478 24799
rect 11572 24760 11578 24772
rect 1176 24704 2268 24732
rect 1176 24692 1182 24704
rect 3510 24692 3516 24744
rect 3568 24692 3574 24744
rect 4062 24692 4068 24744
rect 4120 24732 4126 24744
rect 4430 24732 4436 24744
rect 4120 24704 4436 24732
rect 4120 24692 4126 24704
rect 4430 24692 4436 24704
rect 4488 24692 4494 24744
rect 5378 24735 5436 24741
rect 5378 24732 5390 24735
rect 4540 24704 5390 24732
rect 1581 24667 1639 24673
rect 1581 24633 1593 24667
rect 1627 24664 1639 24667
rect 2590 24664 2596 24676
rect 1627 24636 2596 24664
rect 1627 24633 1639 24636
rect 1581 24627 1639 24633
rect 2590 24624 2596 24636
rect 2648 24624 2654 24676
rect 4154 24624 4160 24676
rect 4212 24624 4218 24676
rect 4246 24624 4252 24676
rect 4304 24664 4310 24676
rect 4540 24664 4568 24704
rect 5378 24701 5390 24704
rect 5424 24701 5436 24735
rect 5378 24695 5436 24701
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 6362 24732 6368 24744
rect 5583 24704 6368 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 6362 24692 6368 24704
rect 6420 24692 6426 24744
rect 11790 24692 11796 24744
rect 11848 24732 11854 24744
rect 12066 24732 12072 24744
rect 11848 24704 12072 24732
rect 11848 24692 11854 24704
rect 12066 24692 12072 24704
rect 12124 24732 12130 24744
rect 12161 24735 12219 24741
rect 12161 24732 12173 24735
rect 12124 24704 12173 24732
rect 12124 24692 12130 24704
rect 12161 24701 12173 24704
rect 12207 24701 12219 24735
rect 16500 24732 16528 24840
rect 16758 24828 16764 24840
rect 16816 24868 16822 24880
rect 17144 24868 17172 24908
rect 17310 24896 17316 24948
rect 17368 24936 17374 24948
rect 17681 24939 17739 24945
rect 17681 24936 17693 24939
rect 17368 24908 17693 24936
rect 17368 24896 17374 24908
rect 17681 24905 17693 24908
rect 17727 24905 17739 24939
rect 17681 24899 17739 24905
rect 21358 24896 21364 24948
rect 21416 24896 21422 24948
rect 21542 24896 21548 24948
rect 21600 24936 21606 24948
rect 21821 24939 21879 24945
rect 21821 24936 21833 24939
rect 21600 24908 21833 24936
rect 21600 24896 21606 24908
rect 21821 24905 21833 24908
rect 21867 24905 21879 24939
rect 21821 24899 21879 24905
rect 23474 24896 23480 24948
rect 23532 24896 23538 24948
rect 18598 24868 18604 24880
rect 16816 24840 17080 24868
rect 17144 24840 18604 24868
rect 16816 24828 16822 24840
rect 16574 24760 16580 24812
rect 16632 24800 16638 24812
rect 16911 24803 16969 24809
rect 16911 24800 16923 24803
rect 16632 24772 16923 24800
rect 16632 24760 16638 24772
rect 16911 24769 16923 24772
rect 16957 24769 16969 24803
rect 17052 24800 17080 24840
rect 18248 24812 18276 24840
rect 18598 24828 18604 24840
rect 18656 24828 18662 24880
rect 19242 24828 19248 24880
rect 19300 24868 19306 24880
rect 19300 24840 20116 24868
rect 19300 24828 19306 24840
rect 17862 24800 17868 24812
rect 17052 24772 17868 24800
rect 16911 24763 16969 24769
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 18230 24760 18236 24812
rect 18288 24800 18294 24812
rect 18323 24803 18381 24809
rect 18323 24800 18335 24803
rect 18288 24772 18335 24800
rect 18288 24760 18294 24772
rect 18323 24769 18335 24772
rect 18369 24769 18381 24803
rect 18323 24763 18381 24769
rect 18690 24760 18696 24812
rect 18748 24800 18754 24812
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 18748 24772 19901 24800
rect 18748 24760 18754 24772
rect 19889 24769 19901 24772
rect 19935 24800 19947 24803
rect 19978 24800 19984 24812
rect 19935 24772 19984 24800
rect 19935 24769 19947 24772
rect 19889 24763 19947 24769
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20088 24800 20116 24840
rect 21376 24809 21404 24896
rect 21634 24828 21640 24880
rect 21692 24868 21698 24880
rect 21692 24840 22131 24868
rect 21692 24828 21698 24840
rect 20145 24803 20203 24809
rect 20145 24800 20157 24803
rect 20088 24772 20157 24800
rect 20145 24769 20157 24772
rect 20191 24769 20203 24803
rect 20145 24763 20203 24769
rect 21361 24803 21419 24809
rect 21361 24769 21373 24803
rect 21407 24769 21419 24803
rect 21361 24763 21419 24769
rect 22005 24803 22063 24809
rect 22005 24769 22017 24803
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 16669 24735 16727 24741
rect 16669 24732 16681 24735
rect 16500 24704 16681 24732
rect 12161 24695 12219 24701
rect 16669 24701 16681 24704
rect 16715 24701 16727 24735
rect 17880 24732 17908 24760
rect 18049 24735 18107 24741
rect 18049 24732 18061 24735
rect 17880 24704 18061 24732
rect 16669 24695 16727 24701
rect 18049 24701 18061 24704
rect 18095 24701 18107 24735
rect 18049 24695 18107 24701
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 21637 24735 21695 24741
rect 21637 24732 21649 24735
rect 21508 24704 21649 24732
rect 21508 24692 21514 24704
rect 21637 24701 21649 24704
rect 21683 24701 21695 24735
rect 21637 24695 21695 24701
rect 4304 24636 4568 24664
rect 4985 24667 5043 24673
rect 4304 24624 4310 24636
rect 4985 24633 4997 24667
rect 5031 24633 5043 24667
rect 8294 24664 8300 24676
rect 4985 24627 5043 24633
rect 5920 24636 8300 24664
rect 2406 24556 2412 24608
rect 2464 24556 2470 24608
rect 5000 24596 5028 24627
rect 5920 24608 5948 24636
rect 8294 24624 8300 24636
rect 8352 24624 8358 24676
rect 9493 24667 9551 24673
rect 9493 24633 9505 24667
rect 9539 24664 9551 24667
rect 9674 24664 9680 24676
rect 9539 24636 9680 24664
rect 9539 24633 9551 24636
rect 9493 24627 9551 24633
rect 9674 24624 9680 24636
rect 9732 24624 9738 24676
rect 10134 24624 10140 24676
rect 10192 24664 10198 24676
rect 10962 24664 10968 24676
rect 10192 24636 10968 24664
rect 10192 24624 10198 24636
rect 10962 24624 10968 24636
rect 11020 24664 11026 24676
rect 11698 24664 11704 24676
rect 11020 24636 11704 24664
rect 11020 24624 11026 24636
rect 11698 24624 11704 24636
rect 11756 24624 11762 24676
rect 21269 24667 21327 24673
rect 13096 24636 13308 24664
rect 5718 24596 5724 24608
rect 5000 24568 5724 24596
rect 5718 24556 5724 24568
rect 5776 24556 5782 24608
rect 5902 24556 5908 24608
rect 5960 24556 5966 24608
rect 6178 24556 6184 24608
rect 6236 24556 6242 24608
rect 8754 24556 8760 24608
rect 8812 24596 8818 24608
rect 13096 24596 13124 24636
rect 8812 24568 13124 24596
rect 8812 24556 8818 24568
rect 13170 24556 13176 24608
rect 13228 24556 13234 24608
rect 13280 24596 13308 24636
rect 21269 24633 21281 24667
rect 21315 24664 21327 24667
rect 22020 24664 22048 24763
rect 22103 24744 22131 24840
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 22707 24803 22765 24809
rect 22707 24800 22719 24803
rect 22428 24772 22719 24800
rect 22428 24760 22434 24772
rect 22707 24769 22719 24772
rect 22753 24769 22765 24803
rect 22707 24763 22765 24769
rect 24121 24803 24179 24809
rect 24121 24769 24133 24803
rect 24167 24800 24179 24803
rect 24302 24800 24308 24812
rect 24167 24772 24308 24800
rect 24167 24769 24179 24772
rect 24121 24763 24179 24769
rect 24302 24760 24308 24772
rect 24360 24760 24366 24812
rect 22094 24692 22100 24744
rect 22152 24732 22158 24744
rect 22465 24735 22523 24741
rect 22465 24732 22477 24735
rect 22152 24704 22477 24732
rect 22152 24692 22158 24704
rect 22465 24701 22477 24704
rect 22511 24701 22523 24735
rect 22465 24695 22523 24701
rect 21315 24636 22048 24664
rect 21315 24633 21327 24636
rect 21269 24627 21327 24633
rect 17770 24596 17776 24608
rect 13280 24568 17776 24596
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 18506 24556 18512 24608
rect 18564 24596 18570 24608
rect 19061 24599 19119 24605
rect 19061 24596 19073 24599
rect 18564 24568 19073 24596
rect 18564 24556 18570 24568
rect 19061 24565 19073 24568
rect 19107 24565 19119 24599
rect 19061 24559 19119 24565
rect 19886 24556 19892 24608
rect 19944 24596 19950 24608
rect 20622 24596 20628 24608
rect 19944 24568 20628 24596
rect 19944 24556 19950 24568
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 21450 24556 21456 24608
rect 21508 24556 21514 24608
rect 21542 24556 21548 24608
rect 21600 24556 21606 24608
rect 24394 24556 24400 24608
rect 24452 24556 24458 24608
rect 1104 24506 24840 24528
rect 1104 24454 3917 24506
rect 3969 24454 3981 24506
rect 4033 24454 4045 24506
rect 4097 24454 4109 24506
rect 4161 24454 4173 24506
rect 4225 24454 9851 24506
rect 9903 24454 9915 24506
rect 9967 24454 9979 24506
rect 10031 24454 10043 24506
rect 10095 24454 10107 24506
rect 10159 24454 15785 24506
rect 15837 24454 15849 24506
rect 15901 24454 15913 24506
rect 15965 24454 15977 24506
rect 16029 24454 16041 24506
rect 16093 24454 21719 24506
rect 21771 24454 21783 24506
rect 21835 24454 21847 24506
rect 21899 24454 21911 24506
rect 21963 24454 21975 24506
rect 22027 24454 24840 24506
rect 1104 24432 24840 24454
rect 2774 24352 2780 24404
rect 2832 24392 2838 24404
rect 5902 24392 5908 24404
rect 2832 24364 5908 24392
rect 2832 24352 2838 24364
rect 5902 24352 5908 24364
rect 5960 24352 5966 24404
rect 6178 24352 6184 24404
rect 6236 24392 6242 24404
rect 6236 24364 6958 24392
rect 6236 24352 6242 24364
rect 2700 24296 5304 24324
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 382 24148 388 24200
rect 440 24148 446 24200
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 1903 24182 2544 24188
rect 2700 24182 2728 24296
rect 2958 24216 2964 24268
rect 3016 24256 3022 24268
rect 4246 24256 4252 24268
rect 3016 24228 4252 24256
rect 3016 24216 3022 24228
rect 4246 24216 4252 24228
rect 4304 24216 4310 24268
rect 4798 24216 4804 24268
rect 4856 24256 4862 24268
rect 5074 24256 5080 24268
rect 4856 24228 5080 24256
rect 4856 24216 4862 24228
rect 5074 24216 5080 24228
rect 5132 24256 5138 24268
rect 5169 24259 5227 24265
rect 5169 24256 5181 24259
rect 5132 24228 5181 24256
rect 5132 24216 5138 24228
rect 5169 24225 5181 24228
rect 5215 24225 5227 24259
rect 5276 24256 5304 24296
rect 5810 24284 5816 24336
rect 5868 24284 5874 24336
rect 5902 24256 5908 24268
rect 5276 24228 5908 24256
rect 5169 24219 5227 24225
rect 5902 24216 5908 24228
rect 5960 24256 5966 24268
rect 6089 24259 6147 24265
rect 6089 24256 6101 24259
rect 5960 24228 6101 24256
rect 5960 24216 5966 24228
rect 6089 24225 6101 24228
rect 6135 24225 6147 24259
rect 6089 24219 6147 24225
rect 6362 24216 6368 24268
rect 6420 24216 6426 24268
rect 5353 24191 5411 24197
rect 5353 24188 5365 24191
rect 1903 24160 2728 24182
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 2516 24154 2728 24160
rect 5184 24160 5365 24188
rect 400 24052 428 24148
rect 5184 24132 5212 24160
rect 5353 24157 5365 24160
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 6178 24148 6184 24200
rect 6236 24197 6242 24200
rect 6236 24191 6264 24197
rect 6252 24157 6264 24191
rect 6930 24188 6958 24364
rect 8570 24352 8576 24404
rect 8628 24392 8634 24404
rect 9674 24392 9680 24404
rect 8628 24364 9680 24392
rect 8628 24352 8634 24364
rect 9674 24352 9680 24364
rect 9732 24392 9738 24404
rect 13078 24392 13084 24404
rect 9732 24364 10640 24392
rect 9732 24352 9738 24364
rect 9953 24327 10011 24333
rect 9953 24293 9965 24327
rect 9999 24324 10011 24327
rect 10042 24324 10048 24336
rect 9999 24296 10048 24324
rect 9999 24293 10011 24296
rect 9953 24287 10011 24293
rect 10042 24284 10048 24296
rect 10100 24284 10106 24336
rect 10612 24265 10640 24364
rect 11440 24364 13084 24392
rect 7009 24259 7067 24265
rect 7009 24225 7021 24259
rect 7055 24256 7067 24259
rect 10597 24259 10655 24265
rect 7055 24228 7972 24256
rect 7055 24225 7067 24228
rect 7009 24219 7067 24225
rect 7944 24197 7972 24228
rect 10597 24225 10609 24259
rect 10643 24225 10655 24259
rect 10597 24219 10655 24225
rect 7285 24191 7343 24197
rect 7285 24188 7297 24191
rect 6930 24160 7297 24188
rect 6236 24151 6264 24157
rect 7285 24157 7297 24160
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7469 24191 7527 24197
rect 7469 24157 7481 24191
rect 7515 24157 7527 24191
rect 7469 24151 7527 24157
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24157 7987 24191
rect 7929 24151 7987 24157
rect 6236 24148 6242 24151
rect 1578 24080 1584 24132
rect 1636 24080 1642 24132
rect 1946 24080 1952 24132
rect 2004 24080 2010 24132
rect 2314 24080 2320 24132
rect 2372 24080 2378 24132
rect 2424 24092 2912 24120
rect 2424 24052 2452 24092
rect 400 24024 2452 24052
rect 2682 24012 2688 24064
rect 2740 24012 2746 24064
rect 2884 24061 2912 24092
rect 4614 24080 4620 24132
rect 4672 24080 4678 24132
rect 5166 24080 5172 24132
rect 5224 24080 5230 24132
rect 7484 24120 7512 24151
rect 8938 24148 8944 24200
rect 8996 24148 9002 24200
rect 9215 24191 9273 24197
rect 9215 24157 9227 24191
rect 9261 24188 9273 24191
rect 9582 24188 9588 24200
rect 9261 24160 9588 24188
rect 9261 24157 9273 24160
rect 9215 24151 9273 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10778 24148 10784 24200
rect 10836 24188 10842 24200
rect 10871 24191 10929 24197
rect 10871 24188 10883 24191
rect 10836 24160 10883 24188
rect 10836 24148 10842 24160
rect 10871 24157 10883 24160
rect 10917 24188 10929 24191
rect 11440 24188 11468 24364
rect 13078 24352 13084 24364
rect 13136 24392 13142 24404
rect 15010 24392 15016 24404
rect 13136 24364 15016 24392
rect 13136 24352 13142 24364
rect 15010 24352 15016 24364
rect 15068 24352 15074 24404
rect 17957 24395 18015 24401
rect 17957 24392 17969 24395
rect 17052 24364 17969 24392
rect 13906 24284 13912 24336
rect 13964 24324 13970 24336
rect 17052 24324 17080 24364
rect 17957 24361 17969 24364
rect 18003 24361 18015 24395
rect 17957 24355 18015 24361
rect 19242 24352 19248 24404
rect 19300 24352 19306 24404
rect 19426 24352 19432 24404
rect 19484 24392 19490 24404
rect 20438 24392 20444 24404
rect 19484 24364 20444 24392
rect 19484 24352 19490 24364
rect 20438 24352 20444 24364
rect 20496 24352 20502 24404
rect 20993 24395 21051 24401
rect 20993 24361 21005 24395
rect 21039 24392 21051 24395
rect 21450 24392 21456 24404
rect 21039 24364 21456 24392
rect 21039 24361 21051 24364
rect 20993 24355 21051 24361
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 23382 24352 23388 24404
rect 23440 24352 23446 24404
rect 23842 24352 23848 24404
rect 23900 24352 23906 24404
rect 13964 24296 15792 24324
rect 13964 24284 13970 24296
rect 12066 24216 12072 24268
rect 12124 24256 12130 24268
rect 12621 24259 12679 24265
rect 12621 24256 12633 24259
rect 12124 24228 12633 24256
rect 12124 24216 12130 24228
rect 12360 24200 12388 24228
rect 12621 24225 12633 24228
rect 12667 24225 12679 24259
rect 12621 24219 12679 24225
rect 14826 24216 14832 24268
rect 14884 24256 14890 24268
rect 15013 24259 15071 24265
rect 15013 24256 15025 24259
rect 14884 24228 15025 24256
rect 14884 24216 14890 24228
rect 15013 24225 15025 24228
rect 15059 24225 15071 24259
rect 15013 24219 15071 24225
rect 15654 24216 15660 24268
rect 15712 24216 15718 24268
rect 15764 24256 15792 24296
rect 16963 24296 17080 24324
rect 16050 24259 16108 24265
rect 16050 24256 16062 24259
rect 15764 24228 16062 24256
rect 16050 24225 16062 24228
rect 16096 24225 16108 24259
rect 16050 24219 16108 24225
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 16963 24256 16991 24296
rect 17678 24284 17684 24336
rect 17736 24324 17742 24336
rect 17862 24324 17868 24336
rect 17736 24296 17868 24324
rect 17736 24284 17742 24296
rect 17862 24284 17868 24296
rect 17920 24324 17926 24336
rect 18690 24324 18696 24336
rect 17920 24296 18696 24324
rect 17920 24284 17926 24296
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 19260 24324 19288 24352
rect 19260 24296 20576 24324
rect 16255 24228 16991 24256
rect 19628 24228 19840 24256
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 19628 24200 19656 24228
rect 10917 24160 11468 24188
rect 10917 24157 10929 24160
rect 10871 24151 10929 24157
rect 12342 24148 12348 24200
rect 12400 24148 12406 24200
rect 15197 24191 15255 24197
rect 12879 24161 12937 24167
rect 12879 24158 12891 24161
rect 7116 24092 7512 24120
rect 2869 24055 2927 24061
rect 2869 24021 2881 24055
rect 2915 24021 2927 24055
rect 4632 24052 4660 24080
rect 6178 24052 6184 24064
rect 4632 24024 6184 24052
rect 2869 24015 2927 24021
rect 6178 24012 6184 24024
rect 6236 24012 6242 24064
rect 7116 24061 7144 24092
rect 7650 24080 7656 24132
rect 7708 24120 7714 24132
rect 11330 24120 11336 24132
rect 7708 24092 11336 24120
rect 7708 24080 7714 24092
rect 11330 24080 11336 24092
rect 11388 24080 11394 24132
rect 12820 24130 12891 24158
rect 12820 24120 12848 24130
rect 12879 24127 12891 24130
rect 12925 24158 12937 24161
rect 12925 24127 12940 24158
rect 15197 24157 15209 24191
rect 15243 24157 15255 24191
rect 15197 24151 15255 24157
rect 12879 24121 12940 24127
rect 11532 24092 12848 24120
rect 12912 24120 12940 24121
rect 12912 24092 14412 24120
rect 7101 24055 7159 24061
rect 7101 24021 7113 24055
rect 7147 24021 7159 24055
rect 7101 24015 7159 24021
rect 7558 24012 7564 24064
rect 7616 24012 7622 24064
rect 7745 24055 7803 24061
rect 7745 24021 7757 24055
rect 7791 24052 7803 24055
rect 8110 24052 8116 24064
rect 7791 24024 8116 24052
rect 7791 24021 7803 24024
rect 7745 24015 7803 24021
rect 8110 24012 8116 24024
rect 8168 24012 8174 24064
rect 8570 24012 8576 24064
rect 8628 24052 8634 24064
rect 9490 24052 9496 24064
rect 8628 24024 9496 24052
rect 8628 24012 8634 24024
rect 9490 24012 9496 24024
rect 9548 24052 9554 24064
rect 11532 24052 11560 24092
rect 14384 24064 14412 24092
rect 9548 24024 11560 24052
rect 11609 24055 11667 24061
rect 9548 24012 9554 24024
rect 11609 24021 11621 24055
rect 11655 24052 11667 24055
rect 12158 24052 12164 24064
rect 11655 24024 12164 24052
rect 11655 24021 11667 24024
rect 11609 24015 11667 24021
rect 12158 24012 12164 24024
rect 12216 24012 12222 24064
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 13814 24052 13820 24064
rect 13679 24024 13820 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 14366 24012 14372 24064
rect 14424 24012 14430 24064
rect 15212 24052 15240 24151
rect 15930 24148 15936 24200
rect 15988 24148 15994 24200
rect 16945 24191 17003 24197
rect 16945 24188 16957 24191
rect 16776 24160 16957 24188
rect 16776 24132 16804 24160
rect 16945 24157 16957 24160
rect 16991 24157 17003 24191
rect 16945 24151 17003 24157
rect 17219 24191 17277 24197
rect 17219 24157 17231 24191
rect 17265 24188 17277 24191
rect 17310 24188 17316 24200
rect 17265 24160 17316 24188
rect 17265 24157 17277 24160
rect 17219 24151 17277 24157
rect 17310 24148 17316 24160
rect 17368 24188 17374 24200
rect 19426 24188 19432 24200
rect 17368 24160 19432 24188
rect 17368 24148 17374 24160
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 19610 24148 19616 24200
rect 19668 24148 19674 24200
rect 19702 24148 19708 24200
rect 19760 24148 19766 24200
rect 19812 24197 19840 24228
rect 20548 24197 20576 24296
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20533 24191 20591 24197
rect 20533 24157 20545 24191
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 20901 24191 20959 24197
rect 20901 24157 20913 24191
rect 20947 24157 20959 24191
rect 20901 24151 20959 24157
rect 23569 24191 23627 24197
rect 23569 24157 23581 24191
rect 23615 24157 23627 24191
rect 23569 24151 23627 24157
rect 16758 24080 16764 24132
rect 16816 24080 16822 24132
rect 19996 24120 20024 24151
rect 20916 24120 20944 24151
rect 19536 24092 20024 24120
rect 20364 24092 20944 24120
rect 23584 24120 23612 24151
rect 23658 24148 23664 24200
rect 23716 24148 23722 24200
rect 23934 24148 23940 24200
rect 23992 24148 23998 24200
rect 25866 24120 25872 24132
rect 23584 24092 25872 24120
rect 15470 24052 15476 24064
rect 15212 24024 15476 24052
rect 15470 24012 15476 24024
rect 15528 24012 15534 24064
rect 16853 24055 16911 24061
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 17494 24052 17500 24064
rect 16899 24024 17500 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 17494 24012 17500 24024
rect 17552 24012 17558 24064
rect 19536 24061 19564 24092
rect 19521 24055 19579 24061
rect 19521 24021 19533 24055
rect 19567 24021 19579 24055
rect 19521 24015 19579 24021
rect 19886 24012 19892 24064
rect 19944 24012 19950 24064
rect 20364 24061 20392 24092
rect 25866 24080 25872 24092
rect 25924 24080 25930 24132
rect 20349 24055 20407 24061
rect 20349 24021 20361 24055
rect 20395 24021 20407 24055
rect 20349 24015 20407 24021
rect 20622 24012 20628 24064
rect 20680 24052 20686 24064
rect 23382 24052 23388 24064
rect 20680 24024 23388 24052
rect 20680 24012 20686 24024
rect 23382 24012 23388 24024
rect 23440 24012 23446 24064
rect 24121 24055 24179 24061
rect 24121 24021 24133 24055
rect 24167 24052 24179 24055
rect 25130 24052 25136 24064
rect 24167 24024 25136 24052
rect 24167 24021 24179 24024
rect 24121 24015 24179 24021
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 1104 23962 25000 23984
rect 1104 23910 6884 23962
rect 6936 23910 6948 23962
rect 7000 23910 7012 23962
rect 7064 23910 7076 23962
rect 7128 23910 7140 23962
rect 7192 23910 12818 23962
rect 12870 23910 12882 23962
rect 12934 23910 12946 23962
rect 12998 23910 13010 23962
rect 13062 23910 13074 23962
rect 13126 23910 18752 23962
rect 18804 23910 18816 23962
rect 18868 23910 18880 23962
rect 18932 23910 18944 23962
rect 18996 23910 19008 23962
rect 19060 23910 24686 23962
rect 24738 23910 24750 23962
rect 24802 23910 24814 23962
rect 24866 23910 24878 23962
rect 24930 23910 24942 23962
rect 24994 23910 25000 23962
rect 1104 23888 25000 23910
rect 2406 23808 2412 23860
rect 2464 23848 2470 23860
rect 2464 23820 2774 23848
rect 2464 23808 2470 23820
rect 2746 23780 2774 23820
rect 3510 23808 3516 23860
rect 3568 23808 3574 23860
rect 4062 23808 4068 23860
rect 4120 23808 4126 23860
rect 7650 23848 7656 23860
rect 5092 23820 7656 23848
rect 5092 23780 5120 23820
rect 7650 23808 7656 23820
rect 7708 23808 7714 23860
rect 8036 23820 10088 23848
rect 8036 23780 8064 23820
rect 2746 23752 5120 23780
rect 7024 23752 8064 23780
rect 2038 23672 2044 23724
rect 2096 23712 2102 23724
rect 2222 23712 2228 23724
rect 2096 23684 2228 23712
rect 2096 23672 2102 23684
rect 2222 23672 2228 23684
rect 2280 23712 2286 23724
rect 2501 23715 2559 23721
rect 2501 23712 2513 23715
rect 2280 23684 2513 23712
rect 2280 23672 2286 23684
rect 2501 23681 2513 23684
rect 2547 23681 2559 23715
rect 2501 23675 2559 23681
rect 2775 23715 2833 23721
rect 2775 23681 2787 23715
rect 2821 23712 2833 23715
rect 3326 23712 3332 23724
rect 2821 23684 3332 23712
rect 2821 23681 2833 23684
rect 2775 23675 2833 23681
rect 3326 23672 3332 23684
rect 3384 23672 3390 23724
rect 3786 23672 3792 23724
rect 3844 23712 3850 23724
rect 3881 23715 3939 23721
rect 3881 23712 3893 23715
rect 3844 23684 3893 23712
rect 3844 23672 3850 23684
rect 3881 23681 3893 23684
rect 3927 23681 3939 23715
rect 3881 23675 3939 23681
rect 3970 23672 3976 23724
rect 4028 23712 4034 23724
rect 7024 23712 7052 23752
rect 8110 23740 8116 23792
rect 8168 23780 8174 23792
rect 8168 23752 8524 23780
rect 8168 23740 8174 23752
rect 4028 23684 7052 23712
rect 7191 23715 7249 23721
rect 4028 23672 4034 23684
rect 7191 23681 7203 23715
rect 7237 23712 7249 23715
rect 7237 23684 8156 23712
rect 7237 23681 7249 23684
rect 7191 23675 7249 23681
rect 1394 23604 1400 23656
rect 1452 23604 1458 23656
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23613 1731 23647
rect 1673 23607 1731 23613
rect 842 23536 848 23588
rect 900 23576 906 23588
rect 1026 23576 1032 23588
rect 900 23548 1032 23576
rect 900 23536 906 23548
rect 1026 23536 1032 23548
rect 1084 23536 1090 23588
rect 1688 23508 1716 23607
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 5350 23644 5356 23656
rect 3476 23616 5356 23644
rect 3476 23604 3482 23616
rect 5350 23604 5356 23616
rect 5408 23604 5414 23656
rect 5442 23604 5448 23656
rect 5500 23644 5506 23656
rect 6917 23647 6975 23653
rect 6917 23644 6929 23647
rect 5500 23616 6929 23644
rect 5500 23604 5506 23616
rect 6917 23613 6929 23616
rect 6963 23613 6975 23647
rect 8128 23644 8156 23684
rect 8202 23672 8208 23724
rect 8260 23712 8266 23724
rect 8496 23721 8524 23752
rect 8754 23740 8760 23792
rect 8812 23780 8818 23792
rect 9600 23789 9628 23820
rect 8849 23783 8907 23789
rect 8849 23780 8861 23783
rect 8812 23752 8861 23780
rect 8812 23740 8818 23752
rect 8849 23749 8861 23752
rect 8895 23749 8907 23783
rect 8849 23743 8907 23749
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9585 23783 9643 23789
rect 9171 23752 9534 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 8297 23715 8355 23721
rect 8297 23712 8309 23715
rect 8260 23684 8309 23712
rect 8260 23672 8266 23684
rect 8297 23681 8309 23684
rect 8343 23681 8355 23715
rect 8297 23675 8355 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23681 8539 23715
rect 8481 23675 8539 23681
rect 9214 23672 9220 23724
rect 9272 23672 9278 23724
rect 9506 23712 9534 23752
rect 9585 23749 9597 23783
rect 9631 23780 9643 23783
rect 9631 23752 9665 23780
rect 9631 23749 9643 23752
rect 9585 23743 9643 23749
rect 9950 23740 9956 23792
rect 10008 23740 10014 23792
rect 10060 23780 10088 23820
rect 10134 23808 10140 23860
rect 10192 23808 10198 23860
rect 11974 23808 11980 23860
rect 12032 23808 12038 23860
rect 12434 23808 12440 23860
rect 12492 23848 12498 23860
rect 13446 23848 13452 23860
rect 12492 23820 13452 23848
rect 12492 23808 12498 23820
rect 13446 23808 13452 23820
rect 13504 23848 13510 23860
rect 13504 23820 14964 23848
rect 13504 23808 13510 23820
rect 11790 23780 11796 23792
rect 10060 23752 11796 23780
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 9766 23712 9772 23724
rect 9506 23684 9772 23712
rect 9766 23672 9772 23684
rect 9824 23712 9830 23724
rect 11698 23712 11704 23724
rect 9824 23684 11704 23712
rect 9824 23672 9830 23684
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 11885 23715 11943 23721
rect 11885 23681 11897 23715
rect 11931 23712 11943 23715
rect 11992 23712 12020 23808
rect 14826 23740 14832 23792
rect 14884 23740 14890 23792
rect 11931 23684 12020 23712
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 8570 23644 8576 23656
rect 8128 23616 8576 23644
rect 6917 23607 6975 23613
rect 2222 23536 2228 23588
rect 2280 23576 2286 23588
rect 2498 23576 2504 23588
rect 2280 23548 2504 23576
rect 2280 23536 2286 23548
rect 2498 23536 2504 23548
rect 2556 23536 2562 23588
rect 3694 23536 3700 23588
rect 3752 23576 3758 23588
rect 6454 23576 6460 23588
rect 3752 23548 6460 23576
rect 3752 23536 3758 23548
rect 6454 23536 6460 23548
rect 6512 23536 6518 23588
rect 6730 23508 6736 23520
rect 1688 23480 6736 23508
rect 6730 23468 6736 23480
rect 6788 23468 6794 23520
rect 6932 23508 6960 23607
rect 8570 23604 8576 23616
rect 8628 23604 8634 23656
rect 10042 23644 10048 23656
rect 9890 23616 10048 23644
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 11146 23604 11152 23656
rect 11204 23644 11210 23656
rect 11900 23644 11928 23675
rect 12250 23672 12256 23724
rect 12308 23672 12314 23724
rect 12618 23672 12624 23724
rect 12676 23672 12682 23724
rect 13630 23672 13636 23724
rect 13688 23721 13694 23724
rect 13688 23715 13716 23721
rect 13704 23681 13716 23715
rect 13688 23675 13716 23681
rect 13688 23672 13694 23675
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 14658 23712 14780 23716
rect 14844 23712 14872 23740
rect 14936 23721 14964 23820
rect 15654 23808 15660 23860
rect 15712 23808 15718 23860
rect 15930 23808 15936 23860
rect 15988 23808 15994 23860
rect 19245 23851 19303 23857
rect 19245 23817 19257 23851
rect 19291 23848 19303 23851
rect 19702 23848 19708 23860
rect 19291 23820 19708 23848
rect 19291 23817 19303 23820
rect 19245 23811 19303 23817
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 22370 23848 22376 23860
rect 22066 23820 22376 23848
rect 14658 23688 14872 23712
rect 11204 23616 11928 23644
rect 12268 23644 12296 23672
rect 12526 23644 12532 23656
rect 12268 23616 12532 23644
rect 11204 23604 11210 23616
rect 12526 23604 12532 23616
rect 12584 23644 12590 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12584 23616 12817 23644
rect 12584 23604 12590 23616
rect 12805 23613 12817 23616
rect 12851 23613 12863 23647
rect 12805 23607 12863 23613
rect 13170 23604 13176 23656
rect 13228 23644 13234 23656
rect 13265 23647 13323 23653
rect 13265 23644 13277 23647
rect 13228 23616 13277 23644
rect 13228 23604 13234 23616
rect 13265 23613 13277 23616
rect 13311 23613 13323 23647
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 13265 23607 13323 23613
rect 13397 23616 13553 23644
rect 7650 23508 7656 23520
rect 6932 23480 7656 23508
rect 7650 23468 7656 23480
rect 7708 23468 7714 23520
rect 7834 23468 7840 23520
rect 7892 23508 7898 23520
rect 7929 23511 7987 23517
rect 7929 23508 7941 23511
rect 7892 23480 7941 23508
rect 7892 23468 7898 23480
rect 7929 23477 7941 23480
rect 7975 23508 7987 23511
rect 8202 23508 8208 23520
rect 7975 23480 8208 23508
rect 7975 23477 7987 23480
rect 7929 23471 7987 23477
rect 8202 23468 8208 23480
rect 8260 23468 8266 23520
rect 8386 23468 8392 23520
rect 8444 23468 8450 23520
rect 12066 23468 12072 23520
rect 12124 23468 12130 23520
rect 13262 23468 13268 23520
rect 13320 23508 13326 23520
rect 13397 23508 13425 23616
rect 13541 23613 13553 23616
rect 13587 23644 13599 23647
rect 13998 23644 14004 23656
rect 13587 23616 14004 23644
rect 13587 23613 13599 23616
rect 13541 23607 13599 23613
rect 13998 23604 14004 23616
rect 14056 23604 14062 23656
rect 14658 23653 14686 23688
rect 14752 23684 14872 23688
rect 14919 23715 14977 23721
rect 14919 23681 14931 23715
rect 14965 23681 14977 23715
rect 15948 23712 15976 23808
rect 16482 23740 16488 23792
rect 16540 23780 16546 23792
rect 22066 23780 22094 23820
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 22833 23851 22891 23857
rect 22833 23817 22845 23851
rect 22879 23817 22891 23851
rect 22833 23811 22891 23817
rect 16540 23752 22094 23780
rect 22848 23780 22876 23811
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 23348 23820 24164 23848
rect 23348 23808 23354 23820
rect 24136 23789 24164 23820
rect 24121 23783 24179 23789
rect 22848 23752 23520 23780
rect 16540 23740 16546 23752
rect 16209 23715 16267 23721
rect 16209 23712 16221 23715
rect 15948 23684 16221 23712
rect 14919 23675 14977 23681
rect 16209 23681 16221 23684
rect 16255 23681 16267 23715
rect 16209 23675 16267 23681
rect 17862 23672 17868 23724
rect 17920 23672 17926 23724
rect 18121 23715 18179 23721
rect 18121 23712 18133 23715
rect 17972 23684 18133 23712
rect 14645 23647 14703 23653
rect 14645 23613 14657 23647
rect 14691 23613 14703 23647
rect 17972 23644 18000 23684
rect 18121 23681 18133 23684
rect 18167 23712 18179 23715
rect 18506 23712 18512 23724
rect 18167 23684 18512 23712
rect 18167 23681 18179 23684
rect 18121 23675 18179 23681
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 19337 23715 19395 23721
rect 19337 23681 19349 23715
rect 19383 23712 19395 23715
rect 19518 23712 19524 23724
rect 19383 23684 19524 23712
rect 19383 23681 19395 23684
rect 19337 23675 19395 23681
rect 19518 23672 19524 23684
rect 19576 23672 19582 23724
rect 19611 23715 19669 23721
rect 19611 23681 19623 23715
rect 19657 23712 19669 23715
rect 20530 23712 20536 23724
rect 19657 23684 20536 23712
rect 19657 23681 19669 23684
rect 19611 23675 19669 23681
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 21634 23672 21640 23724
rect 21692 23712 21698 23724
rect 22738 23712 22744 23724
rect 21692 23684 22744 23712
rect 21692 23672 21698 23684
rect 22738 23672 22744 23684
rect 22796 23712 22802 23724
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 22796 23684 23029 23712
rect 22796 23672 22802 23684
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 23492 23721 23520 23752
rect 24121 23749 24133 23783
rect 24167 23749 24179 23783
rect 24121 23743 24179 23749
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23385 23675 23443 23681
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23681 23535 23715
rect 23477 23675 23535 23681
rect 14645 23607 14703 23613
rect 17880 23616 18000 23644
rect 23400 23644 23428 23675
rect 23934 23672 23940 23724
rect 23992 23672 23998 23724
rect 23400 23616 23796 23644
rect 13320 23480 13425 23508
rect 13320 23468 13326 23480
rect 13998 23468 14004 23520
rect 14056 23508 14062 23520
rect 14274 23508 14280 23520
rect 14056 23480 14280 23508
rect 14056 23468 14062 23480
rect 14274 23468 14280 23480
rect 14332 23468 14338 23520
rect 14461 23511 14519 23517
rect 14461 23477 14473 23511
rect 14507 23508 14519 23511
rect 17880 23508 17908 23616
rect 23768 23585 23796 23616
rect 23753 23579 23811 23585
rect 23753 23545 23765 23579
rect 23799 23545 23811 23579
rect 23753 23539 23811 23545
rect 14507 23480 17908 23508
rect 14507 23477 14519 23480
rect 14461 23471 14519 23477
rect 19610 23468 19616 23520
rect 19668 23508 19674 23520
rect 20349 23511 20407 23517
rect 20349 23508 20361 23511
rect 19668 23480 20361 23508
rect 19668 23468 19674 23480
rect 20349 23477 20361 23480
rect 20395 23477 20407 23511
rect 20349 23471 20407 23477
rect 23290 23468 23296 23520
rect 23348 23468 23354 23520
rect 23566 23468 23572 23520
rect 23624 23468 23630 23520
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 1104 23418 24840 23440
rect 1104 23366 3917 23418
rect 3969 23366 3981 23418
rect 4033 23366 4045 23418
rect 4097 23366 4109 23418
rect 4161 23366 4173 23418
rect 4225 23366 9851 23418
rect 9903 23366 9915 23418
rect 9967 23366 9979 23418
rect 10031 23366 10043 23418
rect 10095 23366 10107 23418
rect 10159 23366 15785 23418
rect 15837 23366 15849 23418
rect 15901 23366 15913 23418
rect 15965 23366 15977 23418
rect 16029 23366 16041 23418
rect 16093 23366 21719 23418
rect 21771 23366 21783 23418
rect 21835 23366 21847 23418
rect 21899 23366 21911 23418
rect 21963 23366 21975 23418
rect 22027 23366 24840 23418
rect 1104 23344 24840 23366
rect 2038 23264 2044 23316
rect 2096 23264 2102 23316
rect 2222 23264 2228 23316
rect 2280 23264 2286 23316
rect 2590 23264 2596 23316
rect 2648 23304 2654 23316
rect 2648 23276 3188 23304
rect 2648 23264 2654 23276
rect 2056 23168 2084 23264
rect 3160 23236 3188 23276
rect 3234 23264 3240 23316
rect 3292 23304 3298 23316
rect 3329 23307 3387 23313
rect 3329 23304 3341 23307
rect 3292 23276 3341 23304
rect 3292 23264 3298 23276
rect 3329 23273 3341 23276
rect 3375 23273 3387 23307
rect 4801 23307 4859 23313
rect 4801 23304 4813 23307
rect 3329 23267 3387 23273
rect 3804 23276 4813 23304
rect 3804 23236 3832 23276
rect 4801 23273 4813 23276
rect 4847 23273 4859 23307
rect 4801 23267 4859 23273
rect 9214 23264 9220 23316
rect 9272 23304 9278 23316
rect 9953 23307 10011 23313
rect 9953 23304 9965 23307
rect 9272 23276 9965 23304
rect 9272 23264 9278 23276
rect 9953 23273 9965 23276
rect 9999 23273 10011 23307
rect 9953 23267 10011 23273
rect 12342 23264 12348 23316
rect 12400 23304 12406 23316
rect 14826 23304 14832 23316
rect 12400 23276 14832 23304
rect 12400 23264 12406 23276
rect 3160 23208 3832 23236
rect 2317 23171 2375 23177
rect 2317 23168 2329 23171
rect 2056 23140 2329 23168
rect 2317 23137 2329 23140
rect 2363 23137 2375 23171
rect 3789 23171 3847 23177
rect 3789 23168 3801 23171
rect 2317 23131 2375 23137
rect 3252 23140 3801 23168
rect 1026 23060 1032 23112
rect 1084 23100 1090 23112
rect 2041 23103 2099 23109
rect 2041 23100 2053 23103
rect 1084 23072 2053 23100
rect 1084 23060 1090 23072
rect 2041 23069 2053 23072
rect 2087 23069 2099 23103
rect 2591 23103 2649 23109
rect 2591 23100 2603 23103
rect 2041 23063 2099 23069
rect 2516 23072 2603 23100
rect 2516 23044 2544 23072
rect 2591 23069 2603 23072
rect 2637 23069 2649 23103
rect 2591 23063 2649 23069
rect 842 22992 848 23044
rect 900 22992 906 23044
rect 2498 22992 2504 23044
rect 2556 22992 2562 23044
rect 860 22964 888 22992
rect 3252 22964 3280 23140
rect 3789 23137 3801 23140
rect 3835 23137 3847 23171
rect 3789 23131 3847 23137
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 11054 23128 11060 23180
rect 11112 23128 11118 23180
rect 14108 23177 14136 23276
rect 14826 23264 14832 23276
rect 14884 23304 14890 23316
rect 15010 23304 15016 23316
rect 14884 23276 15016 23304
rect 14884 23264 14890 23276
rect 15010 23264 15016 23276
rect 15068 23304 15074 23316
rect 16758 23304 16764 23316
rect 15068 23276 16764 23304
rect 15068 23264 15074 23276
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 19886 23264 19892 23316
rect 19944 23264 19950 23316
rect 23753 23307 23811 23313
rect 23753 23273 23765 23307
rect 23799 23304 23811 23307
rect 23934 23304 23940 23316
rect 23799 23276 23940 23304
rect 23799 23273 23811 23276
rect 23753 23267 23811 23273
rect 23934 23264 23940 23276
rect 23992 23264 23998 23316
rect 18417 23239 18475 23245
rect 18417 23205 18429 23239
rect 18463 23205 18475 23239
rect 18417 23199 18475 23205
rect 14093 23171 14151 23177
rect 14093 23137 14105 23171
rect 14139 23137 14151 23171
rect 18432 23168 18460 23199
rect 19904 23177 19932 23264
rect 19337 23171 19395 23177
rect 18432 23140 19288 23168
rect 14093 23131 14151 23137
rect 3326 23060 3332 23112
rect 3384 23100 3390 23112
rect 3384 23090 3740 23100
rect 3896 23090 4108 23100
rect 3384 23073 4108 23090
rect 3384 23072 4059 23073
rect 3384 23060 3390 23072
rect 3712 23062 3924 23072
rect 3326 22964 3332 22976
rect 860 22936 3332 22964
rect 3326 22924 3332 22936
rect 3384 22924 3390 22976
rect 3896 22964 3924 23062
rect 4047 23039 4059 23072
rect 4093 23042 4108 23073
rect 4154 23060 4160 23112
rect 4212 23100 4218 23112
rect 5994 23100 6000 23112
rect 4212 23072 6000 23100
rect 4212 23060 4218 23072
rect 5994 23060 6000 23072
rect 6052 23060 6058 23112
rect 6178 23060 6184 23112
rect 6236 23100 6242 23112
rect 6546 23100 6552 23112
rect 6236 23072 6552 23100
rect 6236 23060 6242 23072
rect 6546 23060 6552 23072
rect 6604 23060 6610 23112
rect 7558 23060 7564 23112
rect 7616 23100 7622 23112
rect 8021 23103 8079 23109
rect 8021 23100 8033 23103
rect 7616 23072 8033 23100
rect 7616 23060 7622 23072
rect 8021 23069 8033 23072
rect 8067 23069 8079 23103
rect 8021 23063 8079 23069
rect 8386 23060 8392 23112
rect 8444 23100 8450 23112
rect 8481 23103 8539 23109
rect 8481 23100 8493 23103
rect 8444 23072 8493 23100
rect 8444 23060 8450 23072
rect 8481 23069 8493 23072
rect 8527 23069 8539 23103
rect 8481 23063 8539 23069
rect 8938 23060 8944 23112
rect 8996 23060 9002 23112
rect 9215 23103 9273 23109
rect 9215 23069 9227 23103
rect 9261 23100 9273 23103
rect 9261 23072 10548 23100
rect 9261 23069 9273 23072
rect 9215 23063 9273 23069
rect 4093 23039 4105 23042
rect 4047 23033 4105 23039
rect 6730 23032 6736 23044
rect 4816 23004 6736 23032
rect 4246 22964 4252 22976
rect 3896 22936 4252 22964
rect 4246 22924 4252 22936
rect 4304 22964 4310 22976
rect 4816 22964 4844 23004
rect 6730 22992 6736 23004
rect 6788 22992 6794 23044
rect 8757 23035 8815 23041
rect 8757 23001 8769 23035
rect 8803 23032 8815 23035
rect 10042 23032 10048 23044
rect 8803 23004 10048 23032
rect 8803 23001 8815 23004
rect 8757 22995 8815 23001
rect 10042 22992 10048 23004
rect 10100 22992 10106 23044
rect 4304 22936 4844 22964
rect 4304 22924 4310 22936
rect 4890 22924 4896 22976
rect 4948 22964 4954 22976
rect 9398 22964 9404 22976
rect 4948 22936 9404 22964
rect 4948 22924 4954 22936
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 10520 22964 10548 23072
rect 10870 23060 10876 23112
rect 10928 23060 10934 23112
rect 10965 23103 11023 23109
rect 10965 23069 10977 23103
rect 11011 23100 11023 23103
rect 12158 23100 12164 23112
rect 11011 23072 12164 23100
rect 11011 23069 11023 23072
rect 10965 23063 11023 23069
rect 12158 23060 12164 23072
rect 12216 23060 12222 23112
rect 14274 23060 14280 23112
rect 14332 23100 14338 23112
rect 14367 23103 14425 23109
rect 14367 23100 14379 23103
rect 14332 23072 14379 23100
rect 14332 23060 14338 23072
rect 14367 23069 14379 23072
rect 14413 23100 14425 23103
rect 15102 23100 15108 23112
rect 14413 23072 15108 23100
rect 14413 23069 14425 23072
rect 14367 23063 14425 23069
rect 15102 23060 15108 23072
rect 15160 23060 15166 23112
rect 16758 23060 16764 23112
rect 16816 23100 16822 23112
rect 17402 23100 17408 23112
rect 16816 23072 17408 23100
rect 16816 23060 16822 23072
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 18506 23060 18512 23112
rect 18564 23100 18570 23112
rect 19260 23109 19288 23140
rect 19337 23137 19349 23171
rect 19383 23168 19395 23171
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 19383 23140 19717 23168
rect 19383 23137 19395 23140
rect 19337 23131 19395 23137
rect 19705 23137 19717 23140
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 19889 23171 19947 23177
rect 19889 23137 19901 23171
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 18601 23103 18659 23109
rect 18601 23100 18613 23103
rect 18564 23072 18613 23100
rect 18564 23060 18570 23072
rect 18601 23069 18613 23072
rect 18647 23069 18659 23103
rect 18601 23063 18659 23069
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19610 23060 19616 23112
rect 19668 23060 19674 23112
rect 19978 23060 19984 23112
rect 20036 23100 20042 23112
rect 20622 23100 20628 23112
rect 20036 23072 20628 23100
rect 20036 23060 20042 23072
rect 20622 23060 20628 23072
rect 20680 23100 20686 23112
rect 20680 23072 21016 23100
rect 20680 23060 20686 23072
rect 10597 23035 10655 23041
rect 10597 23001 10609 23035
rect 10643 23032 10655 23035
rect 11146 23032 11152 23044
rect 10643 23004 11152 23032
rect 10643 23001 10655 23004
rect 10597 22995 10655 23001
rect 11146 22992 11152 23004
rect 11204 22992 11210 23044
rect 11330 22992 11336 23044
rect 11388 22992 11394 23044
rect 11422 22992 11428 23044
rect 11480 22992 11486 23044
rect 11790 22992 11796 23044
rect 11848 23032 11854 23044
rect 19426 23032 19432 23044
rect 11848 23004 19432 23032
rect 11848 22992 11854 23004
rect 19426 22992 19432 23004
rect 19484 22992 19490 23044
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 20870 23035 20928 23041
rect 20870 23032 20882 23035
rect 20772 23004 20882 23032
rect 20772 22992 20778 23004
rect 20870 23001 20882 23004
rect 20916 23001 20928 23035
rect 20988 23032 21016 23072
rect 21726 23060 21732 23112
rect 21784 23100 21790 23112
rect 22097 23103 22155 23109
rect 22097 23100 22109 23103
rect 21784 23072 22109 23100
rect 21784 23060 21790 23072
rect 22097 23069 22109 23072
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 22370 23060 22376 23112
rect 22428 23060 22434 23112
rect 23750 23060 23756 23112
rect 23808 23100 23814 23112
rect 23937 23103 23995 23109
rect 23937 23100 23949 23103
rect 23808 23072 23949 23100
rect 23808 23060 23814 23072
rect 23937 23069 23949 23072
rect 23983 23069 23995 23103
rect 23937 23063 23995 23069
rect 22388 23032 22416 23060
rect 20988 23004 22416 23032
rect 22629 23035 22687 23041
rect 20870 22995 20928 23001
rect 22629 23001 22641 23035
rect 22675 23032 22687 23035
rect 22738 23032 22744 23044
rect 22675 23004 22744 23032
rect 22675 23001 22687 23004
rect 22629 22995 22687 23001
rect 22738 22992 22744 23004
rect 22796 22992 22802 23044
rect 11440 22964 11468 22992
rect 10520 22936 11468 22964
rect 11514 22924 11520 22976
rect 11572 22964 11578 22976
rect 11701 22967 11759 22973
rect 11701 22964 11713 22967
rect 11572 22936 11713 22964
rect 11572 22924 11578 22936
rect 11701 22933 11713 22936
rect 11747 22933 11759 22967
rect 11701 22927 11759 22933
rect 11882 22924 11888 22976
rect 11940 22964 11946 22976
rect 14550 22964 14556 22976
rect 11940 22936 14556 22964
rect 11940 22924 11946 22936
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 15102 22924 15108 22976
rect 15160 22924 15166 22976
rect 17126 22924 17132 22976
rect 17184 22964 17190 22976
rect 17402 22964 17408 22976
rect 17184 22936 17408 22964
rect 17184 22924 17190 22936
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 19889 22967 19947 22973
rect 19889 22933 19901 22967
rect 19935 22964 19947 22967
rect 21358 22964 21364 22976
rect 19935 22936 21364 22964
rect 19935 22933 19947 22936
rect 19889 22927 19947 22933
rect 21358 22924 21364 22936
rect 21416 22924 21422 22976
rect 22005 22967 22063 22973
rect 22005 22933 22017 22967
rect 22051 22964 22063 22967
rect 22094 22964 22100 22976
rect 22051 22936 22100 22964
rect 22051 22933 22063 22936
rect 22005 22927 22063 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22186 22924 22192 22976
rect 22244 22924 22250 22976
rect 24121 22967 24179 22973
rect 24121 22933 24133 22967
rect 24167 22964 24179 22967
rect 25130 22964 25136 22976
rect 24167 22936 25136 22964
rect 24167 22933 24179 22936
rect 24121 22927 24179 22933
rect 25130 22924 25136 22936
rect 25188 22924 25194 22976
rect 1104 22874 25000 22896
rect 1104 22822 6884 22874
rect 6936 22822 6948 22874
rect 7000 22822 7012 22874
rect 7064 22822 7076 22874
rect 7128 22822 7140 22874
rect 7192 22822 12818 22874
rect 12870 22822 12882 22874
rect 12934 22822 12946 22874
rect 12998 22822 13010 22874
rect 13062 22822 13074 22874
rect 13126 22822 18752 22874
rect 18804 22822 18816 22874
rect 18868 22822 18880 22874
rect 18932 22822 18944 22874
rect 18996 22822 19008 22874
rect 19060 22822 24686 22874
rect 24738 22822 24750 22874
rect 24802 22822 24814 22874
rect 24866 22822 24878 22874
rect 24930 22822 24942 22874
rect 24994 22822 25000 22874
rect 1104 22800 25000 22822
rect 2682 22720 2688 22772
rect 2740 22760 2746 22772
rect 3329 22763 3387 22769
rect 2740 22732 3280 22760
rect 2740 22720 2746 22732
rect 1302 22652 1308 22704
rect 1360 22692 1366 22704
rect 3252 22692 3280 22732
rect 3329 22729 3341 22763
rect 3375 22760 3387 22763
rect 3510 22760 3516 22772
rect 3375 22732 3516 22760
rect 3375 22729 3387 22732
rect 3329 22723 3387 22729
rect 3510 22720 3516 22732
rect 3568 22760 3574 22772
rect 6086 22760 6092 22772
rect 3568 22732 6092 22760
rect 3568 22720 3574 22732
rect 6086 22720 6092 22732
rect 6144 22720 6150 22772
rect 8110 22720 8116 22772
rect 8168 22760 8174 22772
rect 10778 22760 10784 22772
rect 8168 22732 10784 22760
rect 8168 22720 8174 22732
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 11054 22720 11060 22772
rect 11112 22720 11118 22772
rect 11422 22720 11428 22772
rect 11480 22760 11486 22772
rect 12250 22760 12256 22772
rect 11480 22732 12256 22760
rect 11480 22720 11486 22732
rect 12250 22720 12256 22732
rect 12308 22720 12314 22772
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 14458 22760 14464 22772
rect 13872 22732 14464 22760
rect 13872 22720 13878 22732
rect 14458 22720 14464 22732
rect 14516 22720 14522 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 15378 22760 15384 22772
rect 14792 22732 15384 22760
rect 14792 22720 14798 22732
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 19426 22720 19432 22772
rect 19484 22760 19490 22772
rect 19886 22760 19892 22772
rect 19484 22732 19892 22760
rect 19484 22720 19490 22732
rect 19886 22720 19892 22732
rect 19944 22720 19950 22772
rect 20714 22720 20720 22772
rect 20772 22720 20778 22772
rect 21085 22763 21143 22769
rect 21085 22729 21097 22763
rect 21131 22760 21143 22763
rect 21726 22760 21732 22772
rect 21131 22732 21732 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 21726 22720 21732 22732
rect 21784 22720 21790 22772
rect 22278 22720 22284 22772
rect 22336 22720 22342 22772
rect 23198 22720 23204 22772
rect 23256 22760 23262 22772
rect 24213 22763 24271 22769
rect 24213 22760 24225 22763
rect 23256 22732 24225 22760
rect 23256 22720 23262 22732
rect 24213 22729 24225 22732
rect 24259 22729 24271 22763
rect 24213 22723 24271 22729
rect 5442 22692 5448 22704
rect 1360 22664 3188 22692
rect 3252 22664 5448 22692
rect 1360 22652 1366 22664
rect 842 22584 848 22636
rect 900 22624 906 22636
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 900 22596 1409 22624
rect 900 22584 906 22596
rect 1320 22488 1348 22596
rect 1397 22593 1409 22596
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 1671 22627 1729 22633
rect 1671 22593 1683 22627
rect 1717 22624 1729 22627
rect 2866 22624 2872 22636
rect 1717 22596 2872 22624
rect 1717 22593 1729 22596
rect 1671 22587 1729 22593
rect 2866 22584 2872 22596
rect 2924 22624 2930 22636
rect 3160 22633 3188 22664
rect 5442 22652 5448 22664
rect 5500 22652 5506 22704
rect 7834 22692 7840 22704
rect 6564 22664 7840 22692
rect 2961 22627 3019 22633
rect 2961 22624 2973 22627
rect 2924 22596 2973 22624
rect 2924 22584 2930 22596
rect 2961 22593 2973 22596
rect 3007 22593 3019 22627
rect 2961 22587 3019 22593
rect 3145 22627 3203 22633
rect 3145 22593 3157 22627
rect 3191 22593 3203 22627
rect 3145 22587 3203 22593
rect 4431 22627 4489 22633
rect 4431 22593 4443 22627
rect 4477 22624 4489 22627
rect 6564 22624 6592 22664
rect 7834 22652 7840 22664
rect 7892 22652 7898 22704
rect 10426 22664 13032 22692
rect 10303 22657 10361 22663
rect 4477 22596 6592 22624
rect 6639 22627 6697 22633
rect 4477 22593 4489 22596
rect 4431 22587 4489 22593
rect 6639 22593 6651 22627
rect 6685 22624 6697 22627
rect 6730 22624 6736 22636
rect 6685 22596 6736 22624
rect 6685 22593 6697 22596
rect 6639 22587 6697 22593
rect 6730 22584 6736 22596
rect 6788 22584 6794 22636
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 10045 22627 10103 22633
rect 10045 22624 10057 22627
rect 9732 22596 10057 22624
rect 9732 22584 9738 22596
rect 10045 22593 10057 22596
rect 10091 22593 10103 22627
rect 10303 22623 10315 22657
rect 10349 22654 10361 22657
rect 10426 22654 10454 22664
rect 10349 22636 10454 22654
rect 10376 22626 10454 22636
rect 10303 22617 10324 22623
rect 10045 22587 10103 22593
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22525 4215 22559
rect 4157 22519 4215 22525
rect 1394 22488 1400 22500
rect 1320 22460 1400 22488
rect 1394 22448 1400 22460
rect 1452 22448 1458 22500
rect 2590 22448 2596 22500
rect 2648 22488 2654 22500
rect 4062 22488 4068 22500
rect 2648 22460 4068 22488
rect 2648 22448 2654 22460
rect 4062 22448 4068 22460
rect 4120 22448 4126 22500
rect 2406 22380 2412 22432
rect 2464 22380 2470 22432
rect 4172 22420 4200 22519
rect 6178 22516 6184 22568
rect 6236 22556 6242 22568
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 6236 22528 6377 22556
rect 6236 22516 6242 22528
rect 6365 22525 6377 22528
rect 6411 22525 6423 22559
rect 6365 22519 6423 22525
rect 4890 22420 4896 22432
rect 4172 22392 4896 22420
rect 4890 22380 4896 22392
rect 4948 22380 4954 22432
rect 5166 22380 5172 22432
rect 5224 22380 5230 22432
rect 6730 22380 6736 22432
rect 6788 22420 6794 22432
rect 7377 22423 7435 22429
rect 7377 22420 7389 22423
rect 6788 22392 7389 22420
rect 6788 22380 6794 22392
rect 7377 22389 7389 22392
rect 7423 22389 7435 22423
rect 10060 22420 10088 22587
rect 10318 22584 10324 22617
rect 10376 22584 10382 22626
rect 12618 22584 12624 22636
rect 12676 22624 12682 22636
rect 12894 22624 12900 22636
rect 12676 22596 12900 22624
rect 12676 22584 12682 22596
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 13004 22624 13032 22664
rect 13170 22652 13176 22704
rect 13228 22692 13234 22704
rect 13446 22692 13452 22704
rect 13228 22664 13452 22692
rect 13228 22652 13234 22664
rect 13446 22652 13452 22664
rect 13504 22652 13510 22704
rect 16666 22652 16672 22704
rect 16724 22652 16730 22704
rect 16574 22624 16580 22636
rect 13004 22596 16580 22624
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 16684 22624 16712 22652
rect 17770 22633 17776 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16684 22596 16865 22624
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 17727 22627 17776 22633
rect 17727 22593 17739 22627
rect 17773 22593 17776 22627
rect 17727 22587 17776 22593
rect 17770 22584 17776 22587
rect 17828 22584 17834 22636
rect 20732 22624 20760 22720
rect 22296 22692 22324 22720
rect 22738 22692 22744 22704
rect 22296 22664 22744 22692
rect 22738 22652 22744 22664
rect 22796 22692 22802 22704
rect 22796 22664 23244 22692
rect 22796 22652 22802 22664
rect 22095 22637 22153 22643
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 20732 22596 21281 22624
rect 21269 22593 21281 22596
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21453 22627 21511 22633
rect 21453 22593 21465 22627
rect 21499 22593 21511 22627
rect 21453 22587 21511 22593
rect 16669 22559 16727 22565
rect 16669 22525 16681 22559
rect 16715 22556 16727 22559
rect 16758 22556 16764 22568
rect 16715 22528 16764 22556
rect 16715 22525 16727 22528
rect 16669 22519 16727 22525
rect 16758 22516 16764 22528
rect 16816 22516 16822 22568
rect 17589 22559 17647 22565
rect 17589 22556 17601 22559
rect 17420 22528 17601 22556
rect 17310 22448 17316 22500
rect 17368 22448 17374 22500
rect 10962 22420 10968 22432
rect 10060 22392 10968 22420
rect 7377 22383 7435 22389
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 12342 22380 12348 22432
rect 12400 22420 12406 22432
rect 12618 22420 12624 22432
rect 12400 22392 12624 22420
rect 12400 22380 12406 22392
rect 12618 22380 12624 22392
rect 12676 22380 12682 22432
rect 14826 22380 14832 22432
rect 14884 22380 14890 22432
rect 15654 22380 15660 22432
rect 15712 22420 15718 22432
rect 16942 22420 16948 22432
rect 15712 22392 16948 22420
rect 15712 22380 15718 22392
rect 16942 22380 16948 22392
rect 17000 22420 17006 22432
rect 17420 22420 17448 22528
rect 17589 22525 17601 22528
rect 17635 22525 17647 22559
rect 17589 22519 17647 22525
rect 17862 22516 17868 22568
rect 17920 22516 17926 22568
rect 21468 22556 21496 22587
rect 21634 22584 21640 22636
rect 21692 22584 21698 22636
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22624 21879 22627
rect 22002 22624 22008 22636
rect 21867 22596 22008 22624
rect 21867 22593 21879 22596
rect 21821 22587 21879 22593
rect 21726 22556 21732 22568
rect 21468 22528 21732 22556
rect 21726 22516 21732 22528
rect 21784 22516 21790 22568
rect 19978 22448 19984 22500
rect 20036 22488 20042 22500
rect 21836 22488 21864 22587
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 22095 22603 22107 22637
rect 22141 22624 22153 22637
rect 22646 22624 22652 22636
rect 22141 22603 22652 22624
rect 22095 22597 22652 22603
rect 22110 22596 22652 22597
rect 22646 22584 22652 22596
rect 22704 22584 22710 22636
rect 23216 22633 23244 22664
rect 23201 22627 23259 22633
rect 23201 22593 23213 22627
rect 23247 22593 23259 22627
rect 23201 22587 23259 22593
rect 23474 22584 23480 22636
rect 23532 22584 23538 22636
rect 20036 22460 21864 22488
rect 20036 22448 20042 22460
rect 17000 22392 17448 22420
rect 17000 22380 17006 22392
rect 18506 22380 18512 22432
rect 18564 22380 18570 22432
rect 19242 22380 19248 22432
rect 19300 22420 19306 22432
rect 20622 22420 20628 22432
rect 19300 22392 20628 22420
rect 19300 22380 19306 22392
rect 20622 22380 20628 22392
rect 20680 22380 20686 22432
rect 21545 22423 21603 22429
rect 21545 22389 21557 22423
rect 21591 22420 21603 22423
rect 22278 22420 22284 22432
rect 21591 22392 22284 22420
rect 21591 22389 21603 22392
rect 21545 22383 21603 22389
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 22830 22380 22836 22432
rect 22888 22380 22894 22432
rect 1104 22330 24840 22352
rect 1104 22278 3917 22330
rect 3969 22278 3981 22330
rect 4033 22278 4045 22330
rect 4097 22278 4109 22330
rect 4161 22278 4173 22330
rect 4225 22278 9851 22330
rect 9903 22278 9915 22330
rect 9967 22278 9979 22330
rect 10031 22278 10043 22330
rect 10095 22278 10107 22330
rect 10159 22278 15785 22330
rect 15837 22278 15849 22330
rect 15901 22278 15913 22330
rect 15965 22278 15977 22330
rect 16029 22278 16041 22330
rect 16093 22278 21719 22330
rect 21771 22278 21783 22330
rect 21835 22278 21847 22330
rect 21899 22278 21911 22330
rect 21963 22278 21975 22330
rect 22027 22278 24840 22330
rect 1104 22256 24840 22278
rect 3050 22176 3056 22228
rect 3108 22176 3114 22228
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 3786 22216 3792 22228
rect 3660 22188 3792 22216
rect 3660 22176 3666 22188
rect 3786 22176 3792 22188
rect 3844 22216 3850 22228
rect 3973 22219 4031 22225
rect 3973 22216 3985 22219
rect 3844 22188 3985 22216
rect 3844 22176 3850 22188
rect 3973 22185 3985 22188
rect 4019 22185 4031 22219
rect 3973 22179 4031 22185
rect 11057 22219 11115 22225
rect 11057 22185 11069 22219
rect 11103 22216 11115 22219
rect 11103 22188 11468 22216
rect 11103 22185 11115 22188
rect 11057 22179 11115 22185
rect 5994 22108 6000 22160
rect 6052 22108 6058 22160
rect 6546 22108 6552 22160
rect 6604 22108 6610 22160
rect 8478 22108 8484 22160
rect 8536 22148 8542 22160
rect 9490 22148 9496 22160
rect 8536 22120 9496 22148
rect 8536 22108 8542 22120
rect 9490 22108 9496 22120
rect 9548 22108 9554 22160
rect 2314 22040 2320 22092
rect 2372 22040 2378 22092
rect 5166 22040 5172 22092
rect 5224 22040 5230 22092
rect 6178 22040 6184 22092
rect 6236 22080 6242 22092
rect 6641 22083 6699 22089
rect 6641 22080 6653 22083
rect 6236 22052 6653 22080
rect 6236 22040 6242 22052
rect 6564 22024 6592 22052
rect 6641 22049 6653 22052
rect 6687 22049 6699 22083
rect 6641 22043 6699 22049
rect 9398 22040 9404 22092
rect 9456 22080 9462 22092
rect 9858 22080 9864 22092
rect 9456 22052 9864 22080
rect 9456 22040 9462 22052
rect 9858 22040 9864 22052
rect 9916 22080 9922 22092
rect 10045 22083 10103 22089
rect 10045 22080 10057 22083
rect 9916 22052 10057 22080
rect 9916 22040 9922 22052
rect 10045 22049 10057 22052
rect 10091 22049 10103 22083
rect 11440 22066 11468 22188
rect 12894 22176 12900 22228
rect 12952 22176 12958 22228
rect 13630 22176 13636 22228
rect 13688 22216 13694 22228
rect 13688 22188 17264 22216
rect 13688 22176 13694 22188
rect 10045 22043 10103 22049
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 14826 22040 14832 22092
rect 14884 22080 14890 22092
rect 15013 22083 15071 22089
rect 15013 22080 15025 22083
rect 14884 22052 15025 22080
rect 14884 22040 14890 22052
rect 15013 22049 15025 22052
rect 15059 22049 15071 22083
rect 15013 22043 15071 22049
rect 15286 22040 15292 22092
rect 15344 22040 15350 22092
rect 17236 22024 17264 22188
rect 17310 22176 17316 22228
rect 17368 22176 17374 22228
rect 18506 22176 18512 22228
rect 18564 22176 18570 22228
rect 22097 22219 22155 22225
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22186 22216 22192 22228
rect 22143 22188 22192 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 22830 22216 22836 22228
rect 22296 22188 22836 22216
rect 1026 21972 1032 22024
rect 1084 22012 1090 22024
rect 1210 22012 1216 22024
rect 1084 21984 1216 22012
rect 1084 21972 1090 21984
rect 1210 21972 1216 21984
rect 1268 21972 1274 22024
rect 2133 22015 2191 22021
rect 2133 21981 2145 22015
rect 2179 22012 2191 22015
rect 2406 22012 2412 22024
rect 2179 21984 2412 22012
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 2501 22015 2559 22021
rect 2501 21981 2513 22015
rect 2547 22012 2559 22015
rect 3142 22012 3148 22024
rect 2547 21984 3148 22012
rect 2547 21981 2559 21984
rect 2501 21975 2559 21981
rect 3142 21972 3148 21984
rect 3200 21972 3206 22024
rect 3234 21972 3240 22024
rect 3292 21972 3298 22024
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 5000 22002 5210 22012
rect 5000 21984 5212 22002
rect 1762 21904 1768 21956
rect 1820 21904 1826 21956
rect 2038 21904 2044 21956
rect 2096 21904 2102 21956
rect 3804 21944 3832 21975
rect 2746 21916 3832 21944
rect 1210 21836 1216 21888
rect 1268 21876 1274 21888
rect 2746 21876 2774 21916
rect 3970 21904 3976 21956
rect 4028 21944 4034 21956
rect 5000 21953 5028 21984
rect 5182 21974 5212 21984
rect 4709 21947 4767 21953
rect 4709 21944 4721 21947
rect 4028 21916 4721 21944
rect 4028 21904 4034 21916
rect 4709 21913 4721 21916
rect 4755 21913 4767 21947
rect 4709 21907 4767 21913
rect 4985 21947 5043 21953
rect 4985 21913 4997 21947
rect 5031 21913 5043 21947
rect 4985 21907 5043 21913
rect 5074 21904 5080 21956
rect 5132 21904 5138 21956
rect 5184 21944 5212 21974
rect 5442 21972 5448 22024
rect 5500 21972 5506 22024
rect 5810 21972 5816 22024
rect 5868 22021 5874 22024
rect 5868 22015 5885 22021
rect 5873 21981 5885 22015
rect 5868 21975 5885 21981
rect 5868 21972 5874 21975
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6822 21972 6828 22024
rect 6880 22012 6886 22024
rect 6915 22015 6973 22021
rect 6915 22012 6927 22015
rect 6880 21984 6927 22012
rect 6880 21972 6886 21984
rect 6915 21981 6927 21984
rect 6961 22012 6973 22015
rect 8202 22012 8208 22024
rect 6961 21984 8208 22012
rect 6961 21981 6973 21984
rect 6915 21975 6973 21981
rect 8202 21972 8208 21984
rect 8260 21972 8266 22024
rect 8570 21972 8576 22024
rect 8628 22012 8634 22024
rect 9030 22012 9036 22024
rect 8628 21984 9036 22012
rect 8628 21972 8634 21984
rect 9030 21972 9036 21984
rect 9088 22012 9094 22024
rect 10287 22015 10345 22021
rect 10287 22012 10299 22015
rect 9088 22002 10042 22012
rect 10152 22002 10299 22012
rect 9088 21984 10299 22002
rect 9088 21972 9094 21984
rect 10014 21974 10180 21984
rect 10287 21981 10299 21984
rect 10333 21981 10345 22015
rect 13354 22012 13360 22024
rect 10287 21975 10345 21981
rect 10428 21984 13360 22012
rect 5184 21916 5580 21944
rect 1268 21848 2774 21876
rect 1268 21836 1274 21848
rect 2866 21836 2872 21888
rect 2924 21836 2930 21888
rect 3142 21836 3148 21888
rect 3200 21876 3206 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 3200 21848 3433 21876
rect 3200 21836 3206 21848
rect 3421 21845 3433 21848
rect 3467 21876 3479 21879
rect 4614 21876 4620 21888
rect 3467 21848 4620 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 5552 21876 5580 21916
rect 5626 21904 5632 21956
rect 5684 21944 5690 21956
rect 10428 21944 10456 21984
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 5684 21916 10456 21944
rect 11164 21916 11744 21944
rect 5684 21904 5690 21916
rect 5902 21876 5908 21888
rect 5552 21848 5908 21876
rect 5902 21836 5908 21848
rect 5960 21876 5966 21888
rect 6178 21876 6184 21888
rect 5960 21848 6184 21876
rect 5960 21836 5966 21848
rect 6178 21836 6184 21848
rect 6236 21836 6242 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 7432 21848 7665 21876
rect 7432 21836 7438 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 7653 21839 7711 21845
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 8662 21876 8668 21888
rect 8444 21848 8668 21876
rect 8444 21836 8450 21848
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 11164 21876 11192 21916
rect 9824 21848 11192 21876
rect 9824 21836 9830 21848
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 11609 21879 11667 21885
rect 11609 21876 11621 21879
rect 11296 21848 11621 21876
rect 11296 21836 11302 21848
rect 11609 21845 11621 21848
rect 11655 21845 11667 21879
rect 11716 21876 11744 21916
rect 11790 21904 11796 21956
rect 11848 21944 11854 21956
rect 11885 21947 11943 21953
rect 11885 21944 11897 21947
rect 11848 21916 11897 21944
rect 11848 21904 11854 21916
rect 11885 21913 11897 21916
rect 11931 21913 11943 21947
rect 11885 21907 11943 21913
rect 11974 21904 11980 21956
rect 12032 21904 12038 21956
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12124 21916 12357 21944
rect 12124 21904 12130 21916
rect 12345 21913 12357 21916
rect 12391 21944 12403 21947
rect 14108 21944 14136 21975
rect 12391 21916 14136 21944
rect 12391 21913 12403 21916
rect 12345 21907 12403 21913
rect 12713 21879 12771 21885
rect 12713 21876 12725 21879
rect 11716 21848 12725 21876
rect 11609 21839 11667 21845
rect 12713 21845 12725 21848
rect 12759 21876 12771 21879
rect 14292 21876 14320 21975
rect 15102 21972 15108 22024
rect 15160 22021 15166 22024
rect 15160 22015 15188 22021
rect 15176 21981 15188 22015
rect 15160 21975 15188 21981
rect 15160 21972 15166 21975
rect 16114 21972 16120 22024
rect 16172 22012 16178 22024
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 16172 21984 16313 22012
rect 16172 21972 16178 21984
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 16301 21975 16359 21981
rect 16482 21972 16488 22024
rect 16540 22012 16546 22024
rect 16575 22015 16633 22021
rect 16575 22012 16587 22015
rect 16540 21984 16587 22012
rect 16540 21972 16546 21984
rect 16575 21981 16587 21984
rect 16621 21981 16633 22015
rect 16575 21975 16633 21981
rect 17218 21972 17224 22024
rect 17276 21972 17282 22024
rect 18417 22015 18475 22021
rect 18417 21981 18429 22015
rect 18463 22012 18475 22015
rect 18524 22012 18552 22176
rect 21634 22108 21640 22160
rect 21692 22148 21698 22160
rect 22296 22148 22324 22188
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 23201 22219 23259 22225
rect 23201 22185 23213 22219
rect 23247 22216 23259 22219
rect 23566 22216 23572 22228
rect 23247 22188 23572 22216
rect 23247 22185 23259 22188
rect 23201 22179 23259 22185
rect 23566 22176 23572 22188
rect 23624 22176 23630 22228
rect 21692 22120 22324 22148
rect 22373 22151 22431 22157
rect 21692 22108 21698 22120
rect 19242 22040 19248 22092
rect 19300 22040 19306 22092
rect 20346 22040 20352 22092
rect 20404 22080 20410 22092
rect 20404 22052 21128 22080
rect 20404 22040 20410 22052
rect 18463 21984 18552 22012
rect 19512 22015 19570 22021
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 19512 21981 19524 22015
rect 19558 22012 19570 22015
rect 20254 22012 20260 22024
rect 19558 21984 20260 22012
rect 19558 21981 19570 21984
rect 19512 21975 19570 21981
rect 16132 21944 16160 21972
rect 15764 21916 16160 21944
rect 17236 21944 17264 21972
rect 19628 21956 19656 21984
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20806 21972 20812 22024
rect 20864 21972 20870 22024
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 17236 21916 19334 21944
rect 12759 21848 14320 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 15378 21836 15384 21888
rect 15436 21876 15442 21888
rect 15764 21876 15792 21916
rect 15436 21848 15792 21876
rect 15933 21879 15991 21885
rect 15436 21836 15442 21848
rect 15933 21845 15945 21879
rect 15979 21876 15991 21879
rect 17678 21876 17684 21888
rect 15979 21848 17684 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 17678 21836 17684 21848
rect 17736 21836 17742 21888
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 18598 21876 18604 21888
rect 18279 21848 18604 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 19306 21876 19334 21916
rect 19610 21904 19616 21956
rect 19668 21904 19674 21956
rect 20438 21944 20444 21956
rect 19720 21916 20444 21944
rect 19720 21876 19748 21916
rect 20438 21904 20444 21916
rect 20496 21904 20502 21956
rect 20714 21904 20720 21956
rect 20772 21944 20778 21956
rect 21008 21944 21036 21975
rect 20772 21916 21036 21944
rect 21100 21944 21128 22052
rect 22020 22021 22048 22120
rect 22373 22117 22385 22151
rect 22419 22148 22431 22151
rect 22462 22148 22468 22160
rect 22419 22120 22468 22148
rect 22419 22117 22431 22120
rect 22373 22111 22431 22117
rect 22462 22108 22468 22120
rect 22520 22108 22526 22160
rect 25682 22108 25688 22160
rect 25740 22108 25746 22160
rect 22278 22040 22284 22092
rect 22336 22040 22342 22092
rect 23290 22040 23296 22092
rect 23348 22080 23354 22092
rect 23385 22083 23443 22089
rect 23385 22080 23397 22083
rect 23348 22052 23397 22080
rect 23348 22040 23354 22052
rect 23385 22049 23397 22052
rect 23431 22049 23443 22083
rect 25700 22080 25728 22108
rect 23385 22043 23443 22049
rect 23584 22052 25728 22080
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 22152 21984 22569 22012
rect 22152 21972 22158 21984
rect 22557 21981 22569 21984
rect 22603 21981 22615 22015
rect 22557 21975 22615 21981
rect 23106 21972 23112 22024
rect 23164 21972 23170 22024
rect 23584 22021 23612 22052
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 24213 22015 24271 22021
rect 24213 21981 24225 22015
rect 24259 22012 24271 22015
rect 25682 22012 25688 22024
rect 24259 21984 25688 22012
rect 24259 21981 24271 21984
rect 24213 21975 24271 21981
rect 25682 21972 25688 21984
rect 25740 21972 25746 22024
rect 23474 21944 23480 21956
rect 21100 21916 23480 21944
rect 20772 21904 20778 21916
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23937 21947 23995 21953
rect 23937 21913 23949 21947
rect 23983 21944 23995 21947
rect 25130 21944 25136 21956
rect 23983 21916 25136 21944
rect 23983 21913 23995 21916
rect 23937 21907 23995 21913
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 19306 21848 19748 21876
rect 20625 21879 20683 21885
rect 20625 21845 20637 21879
rect 20671 21876 20683 21879
rect 20898 21876 20904 21888
rect 20671 21848 20904 21876
rect 20671 21845 20683 21848
rect 20625 21839 20683 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 20990 21836 20996 21888
rect 21048 21836 21054 21888
rect 21358 21836 21364 21888
rect 21416 21876 21422 21888
rect 21634 21876 21640 21888
rect 21416 21848 21640 21876
rect 21416 21836 21422 21848
rect 21634 21836 21640 21848
rect 21692 21836 21698 21888
rect 22278 21836 22284 21888
rect 22336 21836 22342 21888
rect 23382 21836 23388 21888
rect 23440 21836 23446 21888
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 24029 21879 24087 21885
rect 24029 21876 24041 21879
rect 23808 21848 24041 21876
rect 23808 21836 23814 21848
rect 24029 21845 24041 21848
rect 24075 21845 24087 21879
rect 24029 21839 24087 21845
rect 1104 21786 25000 21808
rect 1104 21734 6884 21786
rect 6936 21734 6948 21786
rect 7000 21734 7012 21786
rect 7064 21734 7076 21786
rect 7128 21734 7140 21786
rect 7192 21734 12818 21786
rect 12870 21734 12882 21786
rect 12934 21734 12946 21786
rect 12998 21734 13010 21786
rect 13062 21734 13074 21786
rect 13126 21734 18752 21786
rect 18804 21734 18816 21786
rect 18868 21734 18880 21786
rect 18932 21734 18944 21786
rect 18996 21734 19008 21786
rect 19060 21734 24686 21786
rect 24738 21734 24750 21786
rect 24802 21734 24814 21786
rect 24866 21734 24878 21786
rect 24930 21734 24942 21786
rect 24994 21734 25000 21786
rect 1104 21712 25000 21734
rect 842 21632 848 21684
rect 900 21672 906 21684
rect 1762 21672 1768 21684
rect 900 21644 1768 21672
rect 900 21632 906 21644
rect 1762 21632 1768 21644
rect 1820 21632 1826 21684
rect 2314 21632 2320 21684
rect 2372 21672 2378 21684
rect 2409 21675 2467 21681
rect 2409 21672 2421 21675
rect 2372 21644 2421 21672
rect 2372 21632 2378 21644
rect 2409 21641 2421 21644
rect 2455 21641 2467 21675
rect 2409 21635 2467 21641
rect 2498 21632 2504 21684
rect 2556 21672 2562 21684
rect 2961 21675 3019 21681
rect 2961 21672 2973 21675
rect 2556 21644 2973 21672
rect 2556 21632 2562 21644
rect 2961 21641 2973 21644
rect 3007 21641 3019 21675
rect 2961 21635 3019 21641
rect 3237 21675 3295 21681
rect 3237 21641 3249 21675
rect 3283 21672 3295 21675
rect 4154 21672 4160 21684
rect 3283 21644 4160 21672
rect 3283 21641 3295 21644
rect 3237 21635 3295 21641
rect 1302 21564 1308 21616
rect 1360 21604 1366 21616
rect 2976 21604 3004 21635
rect 4154 21632 4160 21644
rect 4212 21632 4218 21684
rect 5074 21672 5080 21684
rect 5000 21644 5080 21672
rect 3970 21604 3976 21616
rect 1360 21576 2820 21604
rect 2976 21576 3976 21604
rect 1360 21564 1366 21576
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1671 21539 1729 21545
rect 1671 21505 1683 21539
rect 1717 21536 1729 21539
rect 2590 21536 2596 21548
rect 1717 21508 2596 21536
rect 1717 21505 1729 21508
rect 1671 21499 1729 21505
rect 2590 21496 2596 21508
rect 2648 21496 2654 21548
rect 2792 21545 2820 21576
rect 3970 21564 3976 21576
rect 4028 21604 4034 21616
rect 5000 21604 5028 21644
rect 5074 21632 5080 21644
rect 5132 21632 5138 21684
rect 5166 21632 5172 21684
rect 5224 21672 5230 21684
rect 5721 21675 5779 21681
rect 5721 21672 5733 21675
rect 5224 21644 5733 21672
rect 5224 21632 5230 21644
rect 5721 21641 5733 21644
rect 5767 21641 5779 21675
rect 5721 21635 5779 21641
rect 6178 21632 6184 21684
rect 6236 21672 6242 21684
rect 6236 21644 6592 21672
rect 6236 21632 6242 21644
rect 6564 21613 6592 21644
rect 7098 21632 7104 21684
rect 7156 21672 7162 21684
rect 7156 21644 7786 21672
rect 7156 21632 7162 21644
rect 4028 21576 5028 21604
rect 6549 21607 6607 21613
rect 4028 21564 4034 21576
rect 6549 21573 6561 21607
rect 6595 21573 6607 21607
rect 6549 21567 6607 21573
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 6825 21607 6883 21613
rect 6825 21604 6837 21607
rect 6696 21576 6837 21604
rect 6696 21564 6702 21576
rect 6825 21573 6837 21576
rect 6871 21573 6883 21607
rect 6825 21567 6883 21573
rect 6917 21607 6975 21613
rect 6917 21573 6929 21607
rect 6963 21604 6975 21607
rect 7374 21604 7380 21616
rect 6963 21576 7380 21604
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 7650 21564 7656 21616
rect 7708 21564 7714 21616
rect 7758 21604 7786 21644
rect 8478 21632 8484 21684
rect 8536 21632 8542 21684
rect 9585 21675 9643 21681
rect 9585 21641 9597 21675
rect 9631 21672 9643 21675
rect 9674 21672 9680 21684
rect 9631 21644 9680 21672
rect 9631 21641 9643 21644
rect 9585 21635 9643 21641
rect 9674 21632 9680 21644
rect 9732 21632 9738 21684
rect 9769 21675 9827 21681
rect 9769 21641 9781 21675
rect 9815 21672 9827 21675
rect 11054 21672 11060 21684
rect 9815 21644 11060 21672
rect 9815 21641 9827 21644
rect 9769 21635 9827 21641
rect 11054 21632 11060 21644
rect 11112 21632 11118 21684
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 12805 21675 12863 21681
rect 12805 21672 12817 21675
rect 12032 21644 12817 21672
rect 12032 21632 12038 21644
rect 12805 21641 12817 21644
rect 12851 21641 12863 21675
rect 12805 21635 12863 21641
rect 14277 21675 14335 21681
rect 14277 21641 14289 21675
rect 14323 21672 14335 21675
rect 14734 21672 14740 21684
rect 14323 21644 14740 21672
rect 14323 21641 14335 21644
rect 14277 21635 14335 21641
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 20346 21672 20352 21684
rect 14844 21644 20352 21672
rect 14844 21604 14872 21644
rect 20346 21632 20352 21644
rect 20404 21632 20410 21684
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 20864 21644 20913 21672
rect 20864 21632 20870 21644
rect 20901 21641 20913 21644
rect 20947 21641 20959 21675
rect 20901 21635 20959 21641
rect 7758 21576 8984 21604
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 2777 21499 2835 21505
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21505 3111 21539
rect 3053 21499 3111 21505
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21536 4767 21539
rect 4890 21536 4896 21548
rect 4755 21508 4896 21536
rect 4755 21505 4767 21508
rect 4709 21499 4767 21505
rect 3068 21400 3096 21499
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 5000 21545 5166 21546
rect 4983 21539 5166 21545
rect 4983 21505 4995 21539
rect 5029 21536 5166 21539
rect 5902 21536 5908 21548
rect 5029 21518 5908 21536
rect 5029 21505 5041 21518
rect 5138 21508 5908 21518
rect 4983 21499 5041 21505
rect 5902 21496 5908 21508
rect 5960 21496 5966 21548
rect 6086 21496 6092 21548
rect 6144 21536 6150 21548
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 6144 21508 7297 21536
rect 6144 21496 6150 21508
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 8662 21496 8668 21548
rect 8720 21536 8726 21548
rect 8757 21539 8815 21545
rect 8757 21536 8769 21539
rect 8720 21508 8769 21536
rect 8720 21496 8726 21508
rect 8757 21505 8769 21508
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 8846 21496 8852 21548
rect 8904 21496 8910 21548
rect 8956 21536 8984 21576
rect 12544 21576 14872 21604
rect 9214 21536 9220 21548
rect 8956 21508 9220 21536
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 9398 21496 9404 21548
rect 9456 21536 9462 21548
rect 12035 21539 12093 21545
rect 12035 21536 12047 21539
rect 9456 21508 12047 21536
rect 9456 21496 9462 21508
rect 12035 21505 12047 21508
rect 12081 21536 12093 21539
rect 12544 21536 12572 21576
rect 15194 21564 15200 21616
rect 15252 21604 15258 21616
rect 15252 21576 15976 21604
rect 15252 21564 15258 21576
rect 12081 21508 12572 21536
rect 12081 21505 12093 21508
rect 12035 21499 12093 21505
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 13265 21539 13323 21545
rect 13265 21536 13277 21539
rect 12676 21508 13277 21536
rect 12676 21496 12682 21508
rect 13265 21505 13277 21508
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 13539 21539 13597 21545
rect 13539 21505 13551 21539
rect 13585 21536 13597 21539
rect 13630 21536 13636 21548
rect 13585 21508 13636 21536
rect 13585 21505 13597 21508
rect 13539 21499 13597 21505
rect 13630 21496 13636 21508
rect 13688 21496 13694 21548
rect 14274 21496 14280 21548
rect 14332 21536 14338 21548
rect 15010 21536 15016 21548
rect 14332 21508 15016 21536
rect 14332 21496 14338 21508
rect 15010 21496 15016 21508
rect 15068 21536 15074 21548
rect 15105 21539 15163 21545
rect 15105 21536 15117 21539
rect 15068 21508 15117 21536
rect 15068 21496 15074 21508
rect 15105 21505 15117 21508
rect 15151 21505 15163 21539
rect 15378 21536 15384 21548
rect 15339 21508 15384 21536
rect 15105 21499 15163 21505
rect 15378 21496 15384 21508
rect 15436 21496 15442 21548
rect 15470 21496 15476 21548
rect 15528 21536 15534 21548
rect 15838 21536 15844 21548
rect 15528 21508 15844 21536
rect 15528 21496 15534 21508
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 15948 21536 15976 21576
rect 16114 21564 16120 21616
rect 16172 21604 16178 21616
rect 16758 21604 16764 21616
rect 16172 21576 16764 21604
rect 16172 21564 16178 21576
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 18598 21564 18604 21616
rect 18656 21604 18662 21616
rect 18656 21576 18920 21604
rect 18656 21564 18662 21576
rect 17770 21545 17776 21548
rect 17727 21539 17776 21545
rect 15948 21508 16970 21536
rect 8484 21480 8536 21486
rect 6730 21428 6736 21480
rect 6788 21428 6794 21480
rect 9582 21428 9588 21480
rect 9640 21468 9646 21480
rect 11330 21468 11336 21480
rect 9640 21440 11336 21468
rect 9640 21428 9646 21440
rect 11330 21428 11336 21440
rect 11388 21428 11394 21480
rect 11790 21428 11796 21480
rect 11848 21428 11854 21480
rect 16715 21471 16773 21477
rect 16715 21437 16727 21471
rect 16761 21437 16773 21471
rect 16715 21431 16773 21437
rect 8484 21422 8536 21428
rect 2056 21372 3096 21400
rect 1302 21292 1308 21344
rect 1360 21332 1366 21344
rect 2056 21332 2084 21372
rect 4522 21360 4528 21412
rect 4580 21360 4586 21412
rect 1360 21304 2084 21332
rect 1360 21292 1366 21304
rect 3694 21292 3700 21344
rect 3752 21332 3758 21344
rect 4338 21332 4344 21344
rect 3752 21304 4344 21332
rect 3752 21292 3758 21304
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 4540 21332 4568 21360
rect 5810 21332 5816 21344
rect 4540 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 7837 21335 7895 21341
rect 7837 21301 7849 21335
rect 7883 21332 7895 21335
rect 8386 21332 8392 21344
rect 7883 21304 8392 21332
rect 7883 21301 7895 21304
rect 7837 21295 7895 21301
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 11422 21292 11428 21344
rect 11480 21332 11486 21344
rect 13538 21332 13544 21344
rect 11480 21304 13544 21332
rect 11480 21292 11486 21304
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 15010 21292 15016 21344
rect 15068 21292 15074 21344
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 16730 21332 16758 21431
rect 16850 21428 16856 21480
rect 16908 21428 16914 21480
rect 16942 21400 16970 21508
rect 17727 21505 17739 21539
rect 17773 21505 17776 21539
rect 17727 21499 17776 21505
rect 17770 21496 17776 21499
rect 17828 21496 17834 21548
rect 18892 21545 18920 21576
rect 19610 21564 19616 21616
rect 19668 21604 19674 21616
rect 19668 21576 19840 21604
rect 19668 21564 19674 21576
rect 19812 21545 19840 21576
rect 19978 21564 19984 21616
rect 20036 21564 20042 21616
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21536 18567 21539
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18555 21508 18797 21536
rect 18555 21505 18567 21508
rect 18509 21499 18567 21505
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21505 18935 21539
rect 18877 21499 18935 21505
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 19996 21536 20024 21564
rect 19935 21508 20024 21536
rect 20131 21539 20189 21545
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20131 21505 20143 21539
rect 20177 21536 20189 21539
rect 20254 21536 20260 21548
rect 20177 21508 20260 21536
rect 20177 21505 20189 21508
rect 20131 21499 20189 21505
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 17589 21471 17647 21477
rect 17589 21468 17601 21471
rect 17420 21440 17601 21468
rect 17420 21400 17448 21440
rect 17589 21437 17601 21440
rect 17635 21437 17647 21471
rect 17589 21431 17647 21437
rect 17862 21428 17868 21480
rect 17920 21428 17926 21480
rect 16942 21372 17448 21400
rect 18601 21403 18659 21409
rect 18601 21369 18613 21403
rect 18647 21400 18659 21403
rect 19058 21400 19064 21412
rect 18647 21372 19064 21400
rect 18647 21369 18659 21372
rect 18601 21363 18659 21369
rect 19058 21360 19064 21372
rect 19116 21360 19122 21412
rect 19794 21360 19800 21412
rect 19852 21400 19858 21412
rect 19904 21400 19932 21499
rect 20254 21496 20260 21508
rect 20312 21496 20318 21548
rect 20916 21536 20944 21635
rect 20990 21632 20996 21684
rect 21048 21632 21054 21684
rect 21266 21632 21272 21684
rect 21324 21672 21330 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 21324 21644 22017 21672
rect 21324 21632 21330 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 22278 21632 22284 21684
rect 22336 21632 22342 21684
rect 24397 21675 24455 21681
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24486 21672 24492 21684
rect 24443 21644 24492 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 21008 21604 21036 21632
rect 22296 21604 22324 21632
rect 24121 21607 24179 21613
rect 24121 21604 24133 21607
rect 21008 21576 21404 21604
rect 22296 21576 24133 21604
rect 21269 21539 21327 21545
rect 21269 21536 21281 21539
rect 20916 21508 21281 21536
rect 21269 21505 21281 21508
rect 21315 21505 21327 21539
rect 21269 21499 21327 21505
rect 21376 21468 21404 21576
rect 24121 21573 24133 21576
rect 24167 21573 24179 21607
rect 24121 21567 24179 21573
rect 21450 21496 21456 21548
rect 21508 21536 21514 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21508 21508 21833 21536
rect 21508 21496 21514 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 21376 21440 21557 21468
rect 21545 21437 21557 21440
rect 21591 21437 21603 21471
rect 23400 21468 23428 21499
rect 23566 21496 23572 21548
rect 23624 21496 23630 21548
rect 23661 21539 23719 21545
rect 23661 21505 23673 21539
rect 23707 21536 23719 21539
rect 24210 21536 24216 21548
rect 23707 21508 24216 21536
rect 23707 21505 23719 21508
rect 23661 21499 23719 21505
rect 24210 21496 24216 21508
rect 24268 21496 24274 21548
rect 23750 21468 23756 21480
rect 23400 21440 23756 21468
rect 21545 21431 21603 21437
rect 23750 21428 23756 21440
rect 23808 21428 23814 21480
rect 19852 21372 19932 21400
rect 21453 21403 21511 21409
rect 19852 21360 19858 21372
rect 21453 21369 21465 21403
rect 21499 21400 21511 21403
rect 23658 21400 23664 21412
rect 21499 21372 23664 21400
rect 21499 21369 21511 21372
rect 21453 21363 21511 21369
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 17126 21332 17132 21344
rect 16730 21304 17132 21332
rect 17126 21292 17132 21304
rect 17184 21292 17190 21344
rect 17218 21292 17224 21344
rect 17276 21332 17282 21344
rect 17770 21332 17776 21344
rect 17276 21304 17776 21332
rect 17276 21292 17282 21304
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 18969 21335 19027 21341
rect 18969 21332 18981 21335
rect 18840 21304 18981 21332
rect 18840 21292 18846 21304
rect 18969 21301 18981 21304
rect 19015 21301 19027 21335
rect 18969 21295 19027 21301
rect 19610 21292 19616 21344
rect 19668 21292 19674 21344
rect 21358 21292 21364 21344
rect 21416 21292 21422 21344
rect 23474 21292 23480 21344
rect 23532 21292 23538 21344
rect 23842 21292 23848 21344
rect 23900 21292 23906 21344
rect 1104 21242 24840 21264
rect 1104 21190 3917 21242
rect 3969 21190 3981 21242
rect 4033 21190 4045 21242
rect 4097 21190 4109 21242
rect 4161 21190 4173 21242
rect 4225 21190 9851 21242
rect 9903 21190 9915 21242
rect 9967 21190 9979 21242
rect 10031 21190 10043 21242
rect 10095 21190 10107 21242
rect 10159 21190 15785 21242
rect 15837 21190 15849 21242
rect 15901 21190 15913 21242
rect 15965 21190 15977 21242
rect 16029 21190 16041 21242
rect 16093 21190 21719 21242
rect 21771 21190 21783 21242
rect 21835 21190 21847 21242
rect 21899 21190 21911 21242
rect 21963 21190 21975 21242
rect 22027 21190 24840 21242
rect 1104 21168 24840 21190
rect 2501 21131 2559 21137
rect 2501 21097 2513 21131
rect 2547 21128 2559 21131
rect 7098 21128 7104 21140
rect 2547 21100 7104 21128
rect 2547 21097 2559 21100
rect 2501 21091 2559 21097
rect 7098 21088 7104 21100
rect 7156 21088 7162 21140
rect 7484 21100 8432 21128
rect 2777 21063 2835 21069
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 2958 21060 2964 21072
rect 2823 21032 2964 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 2958 21020 2964 21032
rect 3016 21020 3022 21072
rect 1210 20952 1216 21004
rect 1268 20992 1274 21004
rect 7484 21001 7512 21100
rect 8404 21060 8432 21100
rect 8478 21088 8484 21140
rect 8536 21088 8542 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 8904 21100 9965 21128
rect 8904 21088 8910 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 9953 21091 10011 21097
rect 10980 21100 17816 21128
rect 8404 21032 8616 21060
rect 7469 20995 7527 21001
rect 7469 20992 7481 20995
rect 1268 20964 2360 20992
rect 1268 20952 1274 20964
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 1762 20924 1768 20936
rect 1719 20896 1768 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 2332 20933 2360 20964
rect 4724 20964 7481 20992
rect 2317 20927 2375 20933
rect 2317 20893 2329 20927
rect 2363 20893 2375 20927
rect 2317 20887 2375 20893
rect 2593 20927 2651 20933
rect 2593 20893 2605 20927
rect 2639 20893 2651 20927
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 2593 20887 2651 20893
rect 2746 20896 3801 20924
rect 1302 20816 1308 20868
rect 1360 20856 1366 20868
rect 2608 20856 2636 20887
rect 1360 20828 2636 20856
rect 1360 20816 1366 20828
rect 2130 20748 2136 20800
rect 2188 20788 2194 20800
rect 2746 20788 2774 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 3970 20884 3976 20936
rect 4028 20924 4034 20936
rect 4063 20927 4121 20933
rect 4063 20924 4075 20927
rect 4028 20896 4075 20924
rect 4028 20884 4034 20896
rect 4063 20893 4075 20896
rect 4109 20893 4121 20927
rect 4063 20887 4121 20893
rect 3326 20816 3332 20868
rect 3384 20856 3390 20868
rect 4724 20856 4752 20964
rect 7469 20961 7481 20964
rect 7515 20961 7527 20995
rect 7469 20955 7527 20961
rect 8202 20952 8208 21004
rect 8260 20992 8266 21004
rect 8478 20992 8484 21004
rect 8260 20964 8484 20992
rect 8260 20952 8266 20964
rect 8478 20952 8484 20964
rect 8536 20952 8542 21004
rect 8588 20992 8616 21032
rect 8938 20992 8944 21004
rect 8588 20964 8944 20992
rect 8938 20952 8944 20964
rect 8996 20952 9002 21004
rect 9766 20952 9772 21004
rect 9824 20992 9830 21004
rect 10134 20992 10140 21004
rect 9824 20964 10140 20992
rect 9824 20952 9830 20964
rect 10134 20952 10140 20964
rect 10192 20992 10198 21004
rect 10321 20995 10379 21001
rect 10321 20992 10333 20995
rect 10192 20964 10333 20992
rect 10192 20952 10198 20964
rect 10321 20961 10333 20964
rect 10367 20961 10379 20995
rect 10321 20955 10379 20961
rect 5074 20884 5080 20936
rect 5132 20924 5138 20936
rect 5626 20924 5632 20936
rect 5132 20896 5632 20924
rect 5132 20884 5138 20896
rect 5626 20884 5632 20896
rect 5684 20884 5690 20936
rect 5902 20884 5908 20936
rect 5960 20884 5966 20936
rect 7727 20917 7785 20923
rect 3384 20828 4752 20856
rect 5920 20856 5948 20884
rect 7727 20883 7739 20917
rect 7773 20914 7785 20917
rect 7834 20914 7840 20936
rect 7773 20886 7840 20914
rect 7773 20883 7785 20886
rect 7834 20884 7840 20886
rect 7892 20884 7898 20936
rect 9122 20924 9128 20936
rect 8034 20896 9128 20924
rect 7727 20877 7785 20883
rect 5920 20828 7696 20856
rect 3384 20816 3390 20828
rect 2188 20760 2774 20788
rect 2188 20748 2194 20760
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 4801 20791 4859 20797
rect 4801 20788 4813 20791
rect 4120 20760 4813 20788
rect 4120 20748 4126 20760
rect 4801 20757 4813 20760
rect 4847 20757 4859 20791
rect 4801 20751 4859 20757
rect 6086 20748 6092 20800
rect 6144 20788 6150 20800
rect 6362 20788 6368 20800
rect 6144 20760 6368 20788
rect 6144 20748 6150 20760
rect 6362 20748 6368 20760
rect 6420 20748 6426 20800
rect 7668 20788 7696 20828
rect 8034 20788 8062 20896
rect 9122 20884 9128 20896
rect 9180 20933 9186 20936
rect 9180 20927 9241 20933
rect 9180 20893 9195 20927
rect 9229 20893 9241 20927
rect 9180 20887 9241 20893
rect 9180 20884 9186 20887
rect 9858 20884 9864 20936
rect 9916 20924 9922 20936
rect 10563 20927 10621 20933
rect 10563 20924 10575 20927
rect 9916 20896 10575 20924
rect 9916 20884 9922 20896
rect 10563 20893 10575 20896
rect 10609 20893 10621 20927
rect 10563 20887 10621 20893
rect 8938 20816 8944 20868
rect 8996 20856 9002 20868
rect 10980 20856 11008 21100
rect 15010 21020 15016 21072
rect 15068 21060 15074 21072
rect 17788 21060 17816 21100
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 17957 21131 18015 21137
rect 17957 21128 17969 21131
rect 17920 21100 17969 21128
rect 17920 21088 17926 21100
rect 17957 21097 17969 21100
rect 18003 21097 18015 21131
rect 19334 21128 19340 21140
rect 17957 21091 18015 21097
rect 18892 21100 19340 21128
rect 18892 21060 18920 21100
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 19610 21088 19616 21140
rect 19668 21088 19674 21140
rect 20441 21131 20499 21137
rect 20441 21097 20453 21131
rect 20487 21128 20499 21131
rect 21358 21128 21364 21140
rect 20487 21100 21364 21128
rect 20487 21097 20499 21100
rect 20441 21091 20499 21097
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 15068 21032 15516 21060
rect 17788 21032 18920 21060
rect 18969 21063 19027 21069
rect 15068 21020 15074 21032
rect 11790 20952 11796 21004
rect 11848 20992 11854 21004
rect 11974 20992 11980 21004
rect 11848 20964 11980 20992
rect 11848 20952 11854 20964
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 13412 20964 14749 20992
rect 13412 20952 13418 20964
rect 14737 20961 14749 20964
rect 14783 20961 14795 20995
rect 14737 20955 14795 20961
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 15488 20992 15516 21032
rect 18969 21029 18981 21063
rect 19015 21060 19027 21063
rect 19015 21032 19564 21060
rect 19015 21029 19027 21032
rect 18969 21023 19027 21029
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15488 20964 15669 20992
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 15746 20952 15752 21004
rect 15804 21001 15810 21004
rect 15804 20995 15832 21001
rect 15820 20961 15832 20995
rect 15804 20955 15832 20961
rect 15933 20995 15991 21001
rect 15933 20961 15945 20995
rect 15979 20992 15991 20995
rect 16114 20992 16120 21004
rect 15979 20964 16120 20992
rect 15979 20961 15991 20964
rect 15933 20955 15991 20961
rect 15804 20952 15810 20955
rect 16114 20952 16120 20964
rect 16172 20952 16178 21004
rect 16758 20952 16764 21004
rect 16816 20992 16822 21004
rect 16942 20992 16948 21004
rect 16816 20964 16948 20992
rect 16816 20952 16822 20964
rect 16942 20952 16948 20964
rect 17000 20952 17006 21004
rect 18782 20992 18788 21004
rect 18708 20964 18788 20992
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 12158 20924 12164 20936
rect 11204 20896 12164 20924
rect 11204 20884 11210 20896
rect 12158 20884 12164 20896
rect 12216 20933 12222 20936
rect 12216 20927 12277 20933
rect 12216 20893 12231 20927
rect 12265 20893 12277 20927
rect 12216 20887 12277 20893
rect 12216 20884 12222 20887
rect 14826 20884 14832 20936
rect 14884 20924 14890 20936
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 14884 20896 14933 20924
rect 14884 20884 14890 20896
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 16666 20884 16672 20936
rect 16724 20924 16730 20936
rect 17187 20927 17245 20933
rect 17187 20924 17199 20927
rect 16724 20896 17199 20924
rect 16724 20884 16730 20896
rect 17187 20893 17199 20896
rect 17233 20893 17245 20927
rect 17187 20887 17245 20893
rect 18604 20927 18662 20933
rect 18604 20893 18616 20927
rect 18650 20924 18662 20927
rect 18708 20924 18736 20964
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20992 18935 20995
rect 18923 20964 19012 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 18650 20896 18736 20924
rect 18984 20924 19012 20964
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 19116 20964 19472 20992
rect 19116 20952 19122 20964
rect 19150 20924 19156 20936
rect 18984 20896 19156 20924
rect 18650 20893 18662 20896
rect 18604 20887 18662 20893
rect 19150 20884 19156 20896
rect 19208 20924 19214 20936
rect 19444 20933 19472 20964
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 8996 20828 11008 20856
rect 8996 20816 9002 20828
rect 11054 20816 11060 20868
rect 11112 20856 11118 20868
rect 11514 20856 11520 20868
rect 11112 20828 11520 20856
rect 11112 20816 11118 20828
rect 11514 20816 11520 20828
rect 11572 20816 11578 20868
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 13630 20856 13636 20868
rect 12676 20828 13636 20856
rect 12676 20816 12682 20828
rect 13630 20816 13636 20828
rect 13688 20816 13694 20868
rect 19061 20859 19119 20865
rect 19061 20825 19073 20859
rect 19107 20856 19119 20859
rect 19337 20859 19395 20865
rect 19337 20856 19349 20859
rect 19107 20828 19349 20856
rect 19107 20825 19119 20828
rect 19061 20819 19119 20825
rect 19337 20825 19349 20828
rect 19383 20825 19395 20859
rect 19536 20856 19564 21032
rect 19628 20924 19656 21088
rect 20714 21020 20720 21072
rect 20772 21020 20778 21072
rect 20898 21020 20904 21072
rect 20956 21020 20962 21072
rect 20916 20933 20944 21020
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 22388 20964 22569 20992
rect 22388 20936 22416 20964
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 20349 20927 20407 20933
rect 20349 20924 20361 20927
rect 19628 20896 20361 20924
rect 20349 20893 20361 20896
rect 20395 20893 20407 20927
rect 20349 20887 20407 20893
rect 20901 20927 20959 20933
rect 20901 20893 20913 20927
rect 20947 20893 20959 20927
rect 20901 20887 20959 20893
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 22462 20884 22468 20936
rect 22520 20924 22526 20936
rect 24029 20927 24087 20933
rect 24029 20924 24041 20927
rect 22520 20896 24041 20924
rect 22520 20884 22526 20896
rect 24029 20893 24041 20896
rect 24075 20893 24087 20927
rect 24029 20887 24087 20893
rect 20162 20856 20168 20868
rect 19536 20828 20168 20856
rect 19337 20819 19395 20825
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 21174 20816 21180 20868
rect 21232 20856 21238 20868
rect 22646 20856 22652 20868
rect 21232 20828 22652 20856
rect 21232 20816 21238 20828
rect 22646 20816 22652 20828
rect 22704 20856 22710 20868
rect 22802 20859 22860 20865
rect 22802 20856 22814 20859
rect 22704 20828 22814 20856
rect 22704 20816 22710 20828
rect 22802 20825 22814 20828
rect 22848 20825 22860 20859
rect 22802 20819 22860 20825
rect 8202 20788 8208 20800
rect 7668 20760 8208 20788
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 9122 20748 9128 20800
rect 9180 20788 9186 20800
rect 9674 20788 9680 20800
rect 9180 20760 9680 20788
rect 9180 20748 9186 20760
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 10134 20748 10140 20800
rect 10192 20788 10198 20800
rect 10686 20788 10692 20800
rect 10192 20760 10692 20788
rect 10192 20748 10198 20760
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11333 20791 11391 20797
rect 11333 20788 11345 20791
rect 11020 20760 11345 20788
rect 11020 20748 11026 20760
rect 11333 20757 11345 20760
rect 11379 20757 11391 20791
rect 11333 20751 11391 20757
rect 12710 20748 12716 20800
rect 12768 20788 12774 20800
rect 12989 20791 13047 20797
rect 12989 20788 13001 20791
rect 12768 20760 13001 20788
rect 12768 20748 12774 20760
rect 12989 20757 13001 20760
rect 13035 20757 13047 20791
rect 12989 20751 13047 20757
rect 13446 20748 13452 20800
rect 13504 20788 13510 20800
rect 13814 20788 13820 20800
rect 13504 20760 13820 20788
rect 13504 20748 13510 20760
rect 13814 20748 13820 20760
rect 13872 20748 13878 20800
rect 14090 20748 14096 20800
rect 14148 20788 14154 20800
rect 15102 20788 15108 20800
rect 14148 20760 15108 20788
rect 14148 20748 14154 20760
rect 15102 20748 15108 20760
rect 15160 20748 15166 20800
rect 16577 20791 16635 20797
rect 16577 20757 16589 20791
rect 16623 20788 16635 20791
rect 20806 20788 20812 20800
rect 16623 20760 20812 20788
rect 16623 20757 16635 20760
rect 16577 20751 16635 20757
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 23290 20748 23296 20800
rect 23348 20788 23354 20800
rect 23937 20791 23995 20797
rect 23937 20788 23949 20791
rect 23348 20760 23949 20788
rect 23348 20748 23354 20760
rect 23937 20757 23949 20760
rect 23983 20757 23995 20791
rect 23937 20751 23995 20757
rect 24121 20791 24179 20797
rect 24121 20757 24133 20791
rect 24167 20788 24179 20791
rect 24210 20788 24216 20800
rect 24167 20760 24216 20788
rect 24167 20757 24179 20760
rect 24121 20751 24179 20757
rect 24210 20748 24216 20760
rect 24268 20748 24274 20800
rect 1104 20698 25000 20720
rect 1104 20646 6884 20698
rect 6936 20646 6948 20698
rect 7000 20646 7012 20698
rect 7064 20646 7076 20698
rect 7128 20646 7140 20698
rect 7192 20646 12818 20698
rect 12870 20646 12882 20698
rect 12934 20646 12946 20698
rect 12998 20646 13010 20698
rect 13062 20646 13074 20698
rect 13126 20646 18752 20698
rect 18804 20646 18816 20698
rect 18868 20646 18880 20698
rect 18932 20646 18944 20698
rect 18996 20646 19008 20698
rect 19060 20646 24686 20698
rect 24738 20646 24750 20698
rect 24802 20646 24814 20698
rect 24866 20646 24878 20698
rect 24930 20646 24942 20698
rect 24994 20646 25000 20698
rect 1104 20624 25000 20646
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 7834 20584 7840 20596
rect 4028 20556 7840 20584
rect 4028 20544 4034 20556
rect 7834 20544 7840 20556
rect 7892 20544 7898 20596
rect 11238 20584 11244 20596
rect 10704 20556 11244 20584
rect 4890 20516 4896 20528
rect 4816 20488 4896 20516
rect 1671 20451 1729 20457
rect 1671 20417 1683 20451
rect 1717 20448 1729 20451
rect 2038 20448 2044 20460
rect 1717 20420 2044 20448
rect 1717 20417 1729 20420
rect 1671 20411 1729 20417
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 2590 20408 2596 20460
rect 2648 20448 2654 20460
rect 3053 20451 3111 20457
rect 3053 20448 3065 20451
rect 2648 20420 3065 20448
rect 2648 20408 2654 20420
rect 3053 20417 3065 20420
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 3786 20408 3792 20460
rect 3844 20408 3850 20460
rect 3878 20408 3884 20460
rect 3936 20457 3942 20460
rect 3936 20451 3964 20457
rect 3952 20417 3964 20451
rect 3936 20411 3964 20417
rect 3936 20408 3942 20411
rect 4062 20408 4068 20460
rect 4120 20408 4126 20460
rect 4816 20457 4844 20488
rect 4890 20476 4896 20488
rect 4948 20516 4954 20528
rect 6638 20516 6644 20528
rect 4948 20488 6644 20516
rect 4948 20476 4954 20488
rect 6638 20476 6644 20488
rect 6696 20476 6702 20528
rect 9950 20476 9956 20528
rect 10008 20476 10014 20528
rect 10226 20476 10232 20528
rect 10284 20516 10290 20528
rect 10502 20516 10508 20528
rect 10284 20488 10508 20516
rect 10284 20476 10290 20488
rect 10502 20476 10508 20488
rect 10560 20476 10566 20528
rect 10704 20525 10732 20556
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 12526 20584 12532 20596
rect 11624 20556 12532 20584
rect 10689 20519 10747 20525
rect 10689 20485 10701 20519
rect 10735 20485 10747 20519
rect 10689 20479 10747 20485
rect 11057 20519 11115 20525
rect 11057 20485 11069 20519
rect 11103 20516 11115 20519
rect 11146 20516 11152 20528
rect 11103 20488 11152 20516
rect 11103 20485 11115 20488
rect 11057 20479 11115 20485
rect 11146 20476 11152 20488
rect 11204 20516 11210 20528
rect 11624 20516 11652 20556
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 15378 20544 15384 20596
rect 15436 20544 15442 20596
rect 16666 20544 16672 20596
rect 16724 20584 16730 20596
rect 17126 20584 17132 20596
rect 16724 20556 17132 20584
rect 16724 20544 16730 20556
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 18785 20587 18843 20593
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 19150 20584 19156 20596
rect 18831 20556 19156 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 19150 20544 19156 20556
rect 19208 20544 19214 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19610 20584 19616 20596
rect 19484 20556 19616 20584
rect 19484 20544 19490 20556
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 20438 20544 20444 20596
rect 20496 20544 20502 20596
rect 22462 20544 22468 20596
rect 22520 20544 22526 20596
rect 23750 20544 23756 20596
rect 23808 20544 23814 20596
rect 11204 20488 11652 20516
rect 11204 20476 11210 20488
rect 11790 20476 11796 20528
rect 11848 20516 11854 20528
rect 12434 20516 12440 20528
rect 11848 20488 12440 20516
rect 11848 20476 11854 20488
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 5075 20451 5133 20457
rect 5075 20417 5087 20451
rect 5121 20448 5133 20451
rect 8570 20448 8576 20460
rect 5121 20420 8576 20448
rect 5121 20417 5133 20420
rect 5075 20411 5133 20417
rect 8570 20408 8576 20420
rect 8628 20408 8634 20460
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 10594 20448 10600 20460
rect 10367 20420 10600 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 12544 20457 12572 20544
rect 14185 20519 14243 20525
rect 14185 20485 14197 20519
rect 14231 20516 14243 20519
rect 15102 20516 15108 20528
rect 14231 20488 15108 20516
rect 14231 20485 14243 20488
rect 14185 20479 14243 20485
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 18230 20476 18236 20528
rect 18288 20476 18294 20528
rect 20456 20516 20484 20544
rect 20456 20488 22876 20516
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20417 12587 20451
rect 12529 20411 12587 20417
rect 13354 20408 13360 20460
rect 13412 20457 13418 20460
rect 13412 20451 13440 20457
rect 13428 20417 13440 20451
rect 13412 20411 13440 20417
rect 13412 20408 13418 20411
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 14369 20451 14427 20457
rect 14369 20448 14381 20451
rect 14332 20420 14381 20448
rect 14332 20408 14338 20420
rect 14369 20417 14381 20420
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 14643 20451 14701 20457
rect 14643 20448 14655 20451
rect 14608 20420 14655 20448
rect 14608 20408 14614 20420
rect 14643 20417 14655 20420
rect 14689 20448 14701 20451
rect 14734 20448 14740 20460
rect 14689 20420 14740 20448
rect 14689 20417 14701 20420
rect 14643 20411 14701 20417
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17000 20420 17785 20448
rect 17000 20408 17006 20420
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 18047 20451 18105 20457
rect 18047 20417 18059 20451
rect 18093 20448 18105 20451
rect 18248 20448 18276 20476
rect 18093 20420 18276 20448
rect 18093 20417 18105 20420
rect 18047 20411 18105 20417
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22373 20451 22431 20457
rect 22373 20448 22385 20451
rect 22152 20420 22385 20448
rect 22152 20408 22158 20420
rect 22373 20417 22385 20420
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 22646 20408 22652 20460
rect 22704 20408 22710 20460
rect 22738 20408 22744 20460
rect 22796 20408 22802 20460
rect 22848 20448 22876 20488
rect 22922 20448 22928 20460
rect 22848 20420 22928 20448
rect 22922 20408 22928 20420
rect 22980 20457 22986 20460
rect 22980 20451 23041 20457
rect 22980 20417 22995 20451
rect 23029 20417 23041 20451
rect 23768 20448 23796 20544
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23768 20420 24133 20448
rect 22980 20411 23041 20417
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 22980 20408 22986 20411
rect 24210 20408 24216 20460
rect 24268 20408 24274 20460
rect 1394 20340 1400 20392
rect 1452 20340 1458 20392
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 3142 20380 3148 20392
rect 2915 20352 3148 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 3804 20380 3832 20408
rect 10968 20392 11020 20398
rect 3804 20352 4844 20380
rect 3510 20272 3516 20324
rect 3568 20272 3574 20324
rect 2406 20204 2412 20256
rect 2464 20204 2470 20256
rect 4706 20204 4712 20256
rect 4764 20204 4770 20256
rect 4816 20244 4844 20352
rect 11330 20340 11336 20392
rect 11388 20380 11394 20392
rect 12250 20380 12256 20392
rect 11388 20352 12256 20380
rect 11388 20340 11394 20352
rect 12250 20340 12256 20352
rect 12308 20340 12314 20392
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20349 12403 20383
rect 12345 20343 12403 20349
rect 10968 20334 11020 20340
rect 9398 20312 9404 20324
rect 5736 20284 9404 20312
rect 5736 20244 5764 20284
rect 9398 20272 9404 20284
rect 9456 20272 9462 20324
rect 11238 20272 11244 20324
rect 11296 20272 11302 20324
rect 4816 20216 5764 20244
rect 5810 20204 5816 20256
rect 5868 20204 5874 20256
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 7282 20244 7288 20256
rect 5960 20216 7288 20244
rect 5960 20204 5966 20216
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 12360 20244 12388 20343
rect 12710 20340 12716 20392
rect 12768 20380 12774 20392
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12768 20352 13001 20380
rect 12768 20340 12774 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 12989 20343 13047 20349
rect 13265 20383 13323 20389
rect 13265 20349 13277 20383
rect 13311 20380 13323 20383
rect 13906 20380 13912 20392
rect 13311 20352 13912 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 13906 20340 13912 20352
rect 13964 20380 13970 20392
rect 14182 20380 14188 20392
rect 13964 20352 14188 20380
rect 13964 20340 13970 20352
rect 14182 20340 14188 20352
rect 14240 20340 14246 20392
rect 22278 20340 22284 20392
rect 22336 20380 22342 20392
rect 22756 20380 22784 20408
rect 22336 20352 22784 20380
rect 22336 20340 22342 20352
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 23532 20352 24409 20380
rect 23532 20340 23538 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 22189 20315 22247 20321
rect 13924 20284 14320 20312
rect 13924 20244 13952 20284
rect 11388 20216 13952 20244
rect 14292 20244 14320 20284
rect 22189 20281 22201 20315
rect 22235 20312 22247 20315
rect 22646 20312 22652 20324
rect 22235 20284 22652 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 22646 20272 22652 20284
rect 22704 20272 22710 20324
rect 14826 20244 14832 20256
rect 14292 20216 14832 20244
rect 11388 20204 11394 20216
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 18506 20244 18512 20256
rect 16448 20216 18512 20244
rect 16448 20204 16454 20216
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 22830 20204 22836 20256
rect 22888 20244 22894 20256
rect 23842 20244 23848 20256
rect 22888 20216 23848 20244
rect 22888 20204 22894 20216
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 24302 20204 24308 20256
rect 24360 20204 24366 20256
rect 1104 20154 24840 20176
rect 1104 20102 3917 20154
rect 3969 20102 3981 20154
rect 4033 20102 4045 20154
rect 4097 20102 4109 20154
rect 4161 20102 4173 20154
rect 4225 20102 9851 20154
rect 9903 20102 9915 20154
rect 9967 20102 9979 20154
rect 10031 20102 10043 20154
rect 10095 20102 10107 20154
rect 10159 20102 15785 20154
rect 15837 20102 15849 20154
rect 15901 20102 15913 20154
rect 15965 20102 15977 20154
rect 16029 20102 16041 20154
rect 16093 20102 21719 20154
rect 21771 20102 21783 20154
rect 21835 20102 21847 20154
rect 21899 20102 21911 20154
rect 21963 20102 21975 20154
rect 22027 20102 24840 20154
rect 1104 20080 24840 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1854 20040 1860 20052
rect 1627 20012 1860 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 1854 20000 1860 20012
rect 1912 20000 1918 20052
rect 3329 20043 3387 20049
rect 3329 20009 3341 20043
rect 3375 20040 3387 20043
rect 3510 20040 3516 20052
rect 3375 20012 3516 20040
rect 3375 20009 3387 20012
rect 3329 20003 3387 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 4338 20000 4344 20052
rect 4396 20000 4402 20052
rect 9766 20000 9772 20052
rect 9824 20000 9830 20052
rect 10594 20000 10600 20052
rect 10652 20040 10658 20052
rect 11149 20043 11207 20049
rect 11149 20040 11161 20043
rect 10652 20012 11161 20040
rect 10652 20000 10658 20012
rect 11149 20009 11161 20012
rect 11195 20009 11207 20043
rect 11149 20003 11207 20009
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 13262 20040 13268 20052
rect 12032 20012 13268 20040
rect 12032 20000 12038 20012
rect 4356 19972 4384 20000
rect 2976 19944 4384 19972
rect 2130 19864 2136 19916
rect 2188 19904 2194 19916
rect 2317 19907 2375 19913
rect 2317 19904 2329 19907
rect 2188 19876 2329 19904
rect 2188 19864 2194 19876
rect 2317 19873 2329 19876
rect 2363 19873 2375 19907
rect 2317 19867 2375 19873
rect 750 19796 756 19848
rect 808 19836 814 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 808 19808 1501 19836
rect 808 19796 814 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 1489 19799 1547 19805
rect 2038 19796 2044 19848
rect 2096 19836 2102 19848
rect 2559 19839 2617 19845
rect 2559 19836 2571 19839
rect 2096 19808 2571 19836
rect 2096 19796 2102 19808
rect 2559 19805 2571 19808
rect 2605 19836 2617 19839
rect 2976 19836 3004 19944
rect 5810 19864 5816 19916
rect 5868 19864 5874 19916
rect 7650 19864 7656 19916
rect 7708 19904 7714 19916
rect 8018 19904 8024 19916
rect 7708 19876 8024 19904
rect 7708 19864 7714 19876
rect 8018 19864 8024 19876
rect 8076 19864 8082 19916
rect 9784 19904 9812 20000
rect 12544 19913 12572 20012
rect 13262 20000 13268 20012
rect 13320 20000 13326 20052
rect 13538 20000 13544 20052
rect 13596 20000 13602 20052
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 16114 20040 16120 20052
rect 14332 20012 16120 20040
rect 14332 20000 14338 20012
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16632 20012 17264 20040
rect 16632 20000 16638 20012
rect 14458 19932 14464 19984
rect 14516 19972 14522 19984
rect 15378 19972 15384 19984
rect 14516 19944 15384 19972
rect 14516 19932 14522 19944
rect 15378 19932 15384 19944
rect 15436 19932 15442 19984
rect 17236 19972 17264 20012
rect 20898 20000 20904 20052
rect 20956 20040 20962 20052
rect 20956 20012 21772 20040
rect 20956 20000 20962 20012
rect 17770 19972 17776 19984
rect 17236 19944 17776 19972
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9784 19876 10149 19904
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 16298 19864 16304 19916
rect 16356 19864 16362 19916
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16577 19907 16635 19913
rect 16577 19904 16589 19907
rect 16448 19876 16589 19904
rect 16448 19864 16454 19876
rect 16577 19873 16589 19876
rect 16623 19873 16635 19907
rect 16577 19867 16635 19873
rect 16715 19907 16773 19913
rect 16715 19873 16727 19907
rect 16761 19904 16773 19907
rect 17236 19904 17264 19944
rect 17770 19932 17776 19944
rect 17828 19932 17834 19984
rect 16761 19876 17264 19904
rect 16761 19873 16773 19876
rect 16715 19867 16773 19873
rect 17678 19864 17684 19916
rect 17736 19864 17742 19916
rect 19242 19904 19248 19916
rect 19203 19876 19248 19904
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 2605 19808 3004 19836
rect 3789 19839 3847 19845
rect 2605 19805 2617 19808
rect 2559 19799 2617 19805
rect 3789 19805 3801 19839
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 5445 19839 5503 19845
rect 5445 19836 5457 19839
rect 4939 19808 5457 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 5445 19805 5457 19808
rect 5491 19805 5503 19839
rect 5445 19799 5503 19805
rect 1302 19728 1308 19780
rect 1360 19768 1366 19780
rect 3804 19768 3832 19799
rect 5626 19796 5632 19848
rect 5684 19836 5690 19848
rect 5905 19839 5963 19845
rect 5905 19836 5917 19839
rect 5684 19808 5917 19836
rect 5684 19796 5690 19808
rect 5905 19805 5917 19808
rect 5951 19805 5963 19839
rect 5905 19799 5963 19805
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 6915 19839 6973 19845
rect 6687 19808 6776 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 6748 19780 6776 19808
rect 6915 19805 6927 19839
rect 6961 19836 6973 19839
rect 7282 19836 7288 19848
rect 6961 19808 7288 19836
rect 6961 19805 6973 19808
rect 6915 19799 6973 19805
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7374 19796 7380 19848
rect 7432 19836 7438 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 7432 19808 8217 19836
rect 7432 19796 7438 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 10411 19839 10469 19845
rect 10411 19805 10423 19839
rect 10457 19836 10469 19839
rect 10870 19836 10876 19848
rect 10457 19808 10876 19836
rect 10457 19805 10469 19808
rect 10411 19799 10469 19805
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 12802 19845 12808 19848
rect 12771 19839 12808 19845
rect 12771 19805 12783 19839
rect 12771 19799 12808 19805
rect 12802 19796 12808 19799
rect 12860 19796 12866 19848
rect 14274 19796 14280 19848
rect 14332 19836 14338 19848
rect 15657 19839 15715 19845
rect 15657 19836 15669 19839
rect 14332 19808 15669 19836
rect 14332 19796 14338 19808
rect 15657 19805 15669 19808
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19805 15899 19839
rect 15841 19799 15899 19805
rect 1360 19740 3832 19768
rect 1360 19728 1366 19740
rect 4982 19728 4988 19780
rect 5040 19768 5046 19780
rect 5169 19771 5227 19777
rect 5169 19768 5181 19771
rect 5040 19740 5181 19768
rect 5040 19728 5046 19740
rect 5169 19737 5181 19740
rect 5215 19737 5227 19771
rect 5169 19731 5227 19737
rect 5350 19728 5356 19780
rect 5408 19728 5414 19780
rect 5537 19771 5595 19777
rect 5537 19737 5549 19771
rect 5583 19768 5595 19771
rect 5810 19768 5816 19780
rect 5583 19740 5816 19768
rect 5583 19737 5595 19740
rect 5537 19731 5595 19737
rect 5810 19728 5816 19740
rect 5868 19728 5874 19780
rect 6730 19728 6736 19780
rect 6788 19728 6794 19780
rect 6822 19728 6828 19780
rect 6880 19768 6886 19780
rect 6880 19740 7786 19768
rect 6880 19728 6886 19740
rect 3973 19703 4031 19709
rect 3973 19669 3985 19703
rect 4019 19700 4031 19703
rect 5368 19700 5396 19728
rect 6273 19703 6331 19709
rect 6273 19700 6285 19703
rect 4019 19672 6285 19700
rect 4019 19669 4031 19672
rect 3973 19663 4031 19669
rect 6273 19669 6285 19672
rect 6319 19669 6331 19703
rect 6273 19663 6331 19669
rect 6454 19660 6460 19712
rect 6512 19660 6518 19712
rect 7650 19660 7656 19712
rect 7708 19660 7714 19712
rect 7758 19700 7786 19740
rect 9122 19728 9128 19780
rect 9180 19768 9186 19780
rect 15010 19768 15016 19780
rect 9180 19740 15016 19768
rect 9180 19728 9186 19740
rect 15010 19728 15016 19740
rect 15068 19768 15074 19780
rect 15856 19768 15884 19799
rect 16850 19796 16856 19848
rect 16908 19796 16914 19848
rect 17696 19836 17724 19864
rect 19061 19839 19119 19845
rect 19061 19836 19073 19839
rect 17696 19808 19073 19836
rect 19061 19805 19073 19808
rect 19107 19805 19119 19839
rect 19260 19836 19288 19864
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 19260 19808 20729 19836
rect 19061 19799 19119 19805
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 15068 19740 15884 19768
rect 19076 19768 19104 19799
rect 20806 19796 20812 19848
rect 20864 19836 20870 19848
rect 20973 19839 21031 19845
rect 20973 19836 20985 19839
rect 20864 19808 20985 19836
rect 20864 19796 20870 19808
rect 20973 19805 20985 19808
rect 21019 19836 21031 19839
rect 21266 19836 21272 19848
rect 21019 19808 21272 19836
rect 21019 19805 21031 19808
rect 20973 19799 21031 19805
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 21744 19836 21772 20012
rect 22094 20000 22100 20052
rect 22152 20000 22158 20052
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 22462 20040 22468 20052
rect 22336 20012 22468 20040
rect 22336 20000 22342 20012
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 23937 20043 23995 20049
rect 23937 20009 23949 20043
rect 23983 20040 23995 20043
rect 24026 20040 24032 20052
rect 23983 20012 24032 20040
rect 23983 20009 23995 20012
rect 23937 20003 23995 20009
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 22296 19972 22324 20000
rect 22204 19944 22324 19972
rect 22204 19913 22232 19944
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 22431 19839 22489 19845
rect 22431 19836 22443 19839
rect 21744 19808 22443 19836
rect 22431 19805 22443 19808
rect 22477 19805 22489 19839
rect 22431 19799 22489 19805
rect 23658 19796 23664 19848
rect 23716 19796 23722 19848
rect 19490 19771 19548 19777
rect 19490 19768 19502 19771
rect 19076 19740 19502 19768
rect 15068 19728 15074 19740
rect 19490 19737 19502 19740
rect 19536 19737 19548 19771
rect 19490 19731 19548 19737
rect 21082 19728 21088 19780
rect 21140 19768 21146 19780
rect 24210 19768 24216 19780
rect 21140 19740 24216 19768
rect 21140 19728 21146 19740
rect 24210 19728 24216 19740
rect 24268 19728 24274 19780
rect 11330 19700 11336 19712
rect 7758 19672 11336 19700
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 14090 19700 14096 19712
rect 12768 19672 14096 19700
rect 12768 19660 12774 19672
rect 14090 19660 14096 19672
rect 14148 19700 14154 19712
rect 16942 19700 16948 19712
rect 14148 19672 16948 19700
rect 14148 19660 14154 19672
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 18138 19700 18144 19712
rect 17543 19672 18144 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 18877 19703 18935 19709
rect 18877 19669 18889 19703
rect 18923 19700 18935 19703
rect 19150 19700 19156 19712
rect 18923 19672 19156 19700
rect 18923 19669 18935 19672
rect 18877 19663 18935 19669
rect 19150 19660 19156 19672
rect 19208 19660 19214 19712
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 23198 19660 23204 19712
rect 23256 19660 23262 19712
rect 1104 19610 25000 19632
rect 1104 19558 6884 19610
rect 6936 19558 6948 19610
rect 7000 19558 7012 19610
rect 7064 19558 7076 19610
rect 7128 19558 7140 19610
rect 7192 19558 12818 19610
rect 12870 19558 12882 19610
rect 12934 19558 12946 19610
rect 12998 19558 13010 19610
rect 13062 19558 13074 19610
rect 13126 19558 18752 19610
rect 18804 19558 18816 19610
rect 18868 19558 18880 19610
rect 18932 19558 18944 19610
rect 18996 19558 19008 19610
rect 19060 19558 24686 19610
rect 24738 19558 24750 19610
rect 24802 19558 24814 19610
rect 24866 19558 24878 19610
rect 24930 19558 24942 19610
rect 24994 19558 25000 19610
rect 1104 19536 25000 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 1946 19456 1952 19508
rect 2004 19496 2010 19508
rect 3053 19499 3111 19505
rect 3053 19496 3065 19499
rect 2004 19468 3065 19496
rect 2004 19456 2010 19468
rect 3053 19465 3065 19468
rect 3099 19465 3111 19499
rect 3053 19459 3111 19465
rect 3513 19499 3571 19505
rect 3513 19465 3525 19499
rect 3559 19496 3571 19499
rect 4614 19496 4620 19508
rect 3559 19468 4620 19496
rect 3559 19465 3571 19468
rect 3513 19459 3571 19465
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 4706 19456 4712 19508
rect 4764 19456 4770 19508
rect 5810 19456 5816 19508
rect 5868 19496 5874 19508
rect 5905 19499 5963 19505
rect 5905 19496 5917 19499
rect 5868 19468 5917 19496
rect 5868 19456 5874 19468
rect 5905 19465 5917 19468
rect 5951 19465 5963 19499
rect 5905 19459 5963 19465
rect 6362 19456 6368 19508
rect 6420 19496 6426 19508
rect 7101 19499 7159 19505
rect 7101 19496 7113 19499
rect 6420 19468 7113 19496
rect 6420 19456 6426 19468
rect 7101 19465 7113 19468
rect 7147 19496 7159 19499
rect 7742 19496 7748 19508
rect 7147 19468 7748 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 8202 19456 8208 19508
rect 8260 19456 8266 19508
rect 9122 19496 9128 19508
rect 8772 19468 9128 19496
rect 4724 19428 4752 19456
rect 3252 19400 4752 19428
rect 4816 19400 7788 19428
rect 842 19320 848 19372
rect 900 19360 906 19372
rect 1397 19363 1455 19369
rect 1397 19360 1409 19363
rect 900 19332 1409 19360
rect 900 19320 906 19332
rect 1397 19329 1409 19332
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 1854 19360 1860 19372
rect 1719 19332 1860 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 1947 19363 2005 19369
rect 1947 19329 1959 19363
rect 1993 19360 2005 19363
rect 2038 19360 2044 19372
rect 1993 19332 2044 19360
rect 1993 19329 2005 19332
rect 1947 19323 2005 19329
rect 2038 19320 2044 19332
rect 2096 19320 2102 19372
rect 3252 19369 3280 19400
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3326 19320 3332 19372
rect 3384 19320 3390 19372
rect 3786 19320 3792 19372
rect 3844 19320 3850 19372
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 4816 19360 4844 19400
rect 4672 19332 4844 19360
rect 4672 19320 4678 19332
rect 4890 19320 4896 19372
rect 4948 19320 4954 19372
rect 5167 19363 5225 19369
rect 5167 19329 5179 19363
rect 5213 19360 5225 19363
rect 7190 19360 7196 19372
rect 5213 19332 7196 19360
rect 5213 19329 5225 19332
rect 5167 19323 5225 19329
rect 7190 19320 7196 19332
rect 7248 19320 7254 19372
rect 7374 19320 7380 19372
rect 7432 19320 7438 19372
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 7760 19360 7788 19400
rect 7834 19388 7840 19440
rect 7892 19388 7898 19440
rect 8772 19428 8800 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 9214 19456 9220 19508
rect 9272 19496 9278 19508
rect 14274 19496 14280 19508
rect 9272 19468 14280 19496
rect 9272 19456 9278 19468
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 16850 19456 16856 19508
rect 16908 19496 16914 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 16908 19468 17693 19496
rect 16908 19456 16914 19468
rect 17681 19465 17693 19468
rect 17727 19465 17739 19499
rect 17681 19459 17739 19465
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 19978 19496 19984 19508
rect 19300 19468 19984 19496
rect 19300 19456 19306 19468
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19465 20223 19499
rect 20165 19459 20223 19465
rect 20809 19499 20867 19505
rect 20809 19465 20821 19499
rect 20855 19496 20867 19499
rect 21082 19496 21088 19508
rect 20855 19468 21088 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 12710 19428 12716 19440
rect 7944 19400 8800 19428
rect 8864 19400 12716 19428
rect 7944 19360 7972 19400
rect 7760 19332 7972 19360
rect 8018 19320 8024 19372
rect 8076 19360 8082 19372
rect 8864 19369 8892 19400
rect 12710 19388 12716 19400
rect 12768 19388 12774 19440
rect 13538 19388 13544 19440
rect 13596 19388 13602 19440
rect 13906 19388 13912 19440
rect 13964 19428 13970 19440
rect 19794 19428 19800 19440
rect 13964 19400 16954 19428
rect 13964 19388 13970 19400
rect 8849 19363 8907 19369
rect 8849 19360 8861 19363
rect 8076 19332 8861 19360
rect 8076 19320 8082 19332
rect 3804 19292 3832 19320
rect 3804 19264 4936 19292
rect 2682 19116 2688 19168
rect 2740 19116 2746 19168
rect 4908 19156 4936 19264
rect 7650 19252 7656 19304
rect 7708 19252 7714 19304
rect 8312 19168 8340 19332
rect 8849 19329 8861 19332
rect 8895 19329 8907 19363
rect 8849 19323 8907 19329
rect 9123 19363 9181 19369
rect 9123 19329 9135 19363
rect 9169 19360 9181 19363
rect 10594 19360 10600 19372
rect 9169 19332 10600 19360
rect 9169 19329 9181 19332
rect 9123 19323 9181 19329
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 11790 19360 11796 19372
rect 11751 19332 11796 19360
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 12728 19360 12756 19388
rect 13437 19363 13495 19369
rect 13437 19360 13449 19363
rect 12728 19332 13449 19360
rect 13437 19329 13449 19332
rect 13483 19329 13495 19363
rect 13556 19360 13584 19388
rect 13691 19363 13749 19369
rect 13691 19360 13703 19363
rect 13556 19332 13703 19360
rect 13437 19323 13495 19329
rect 13691 19329 13703 19332
rect 13737 19329 13749 19363
rect 13691 19323 13749 19329
rect 16390 19320 16396 19372
rect 16448 19320 16454 19372
rect 16926 19369 16954 19400
rect 19168 19400 19800 19428
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 16911 19363 16969 19369
rect 16911 19329 16923 19363
rect 16957 19329 16969 19363
rect 16911 19323 16969 19329
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 11514 19292 11520 19304
rect 11296 19264 11520 19292
rect 11296 19252 11302 19264
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 16408 19292 16436 19320
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 16408 19264 16497 19292
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 11054 19224 11060 19236
rect 9600 19196 11060 19224
rect 5810 19156 5816 19168
rect 4908 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 8294 19116 8300 19168
rect 8352 19116 8358 19168
rect 8389 19159 8447 19165
rect 8389 19125 8401 19159
rect 8435 19156 8447 19159
rect 9600 19156 9628 19196
rect 11054 19184 11060 19196
rect 11112 19184 11118 19236
rect 8435 19128 9628 19156
rect 8435 19125 8447 19128
rect 8389 19119 8447 19125
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9732 19128 9873 19156
rect 9732 19116 9738 19128
rect 9861 19125 9873 19128
rect 9907 19125 9919 19159
rect 9861 19119 9919 19125
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10410 19156 10416 19168
rect 10192 19128 10416 19156
rect 10192 19116 10198 19128
rect 10410 19116 10416 19128
rect 10468 19116 10474 19168
rect 12526 19116 12532 19168
rect 12584 19116 12590 19168
rect 14458 19116 14464 19168
rect 14516 19116 14522 19168
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16684 19156 16712 19323
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19168 19369 19196 19400
rect 19794 19388 19800 19400
rect 19852 19388 19858 19440
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 19116 19332 19165 19360
rect 19116 19320 19122 19332
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19426 19320 19432 19372
rect 19484 19320 19490 19372
rect 20180 19360 20208 19459
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19465 21235 19499
rect 21177 19459 21235 19465
rect 20438 19388 20444 19440
rect 20496 19428 20502 19440
rect 21192 19428 21220 19459
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22373 19499 22431 19505
rect 22373 19496 22385 19499
rect 22244 19468 22385 19496
rect 22244 19456 22250 19468
rect 22373 19465 22385 19468
rect 22419 19465 22431 19499
rect 22373 19459 22431 19465
rect 23198 19456 23204 19508
rect 23256 19456 23262 19508
rect 23290 19456 23296 19508
rect 23348 19456 23354 19508
rect 23566 19456 23572 19508
rect 23624 19456 23630 19508
rect 23842 19456 23848 19508
rect 23900 19496 23906 19508
rect 23900 19468 25636 19496
rect 23900 19456 23906 19468
rect 23216 19428 23244 19456
rect 20496 19400 21128 19428
rect 21192 19400 21864 19428
rect 20496 19388 20502 19400
rect 21100 19369 21128 19400
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 20180 19332 20545 19360
rect 20533 19329 20545 19332
rect 20579 19360 20591 19363
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 20579 19332 20913 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20901 19329 20913 19332
rect 20947 19329 20959 19363
rect 20901 19323 20959 19329
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21836 19369 21864 19400
rect 22480 19400 23244 19428
rect 22480 19369 22508 19400
rect 21361 19363 21419 19369
rect 21361 19360 21373 19363
rect 21324 19332 21373 19360
rect 21324 19320 21330 19332
rect 21361 19329 21373 19332
rect 21407 19329 21419 19363
rect 21361 19323 21419 19329
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 22143 19332 22477 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 22646 19320 22652 19372
rect 22704 19320 22710 19372
rect 22922 19320 22928 19372
rect 22980 19360 22986 19372
rect 23308 19360 23336 19456
rect 23584 19428 23612 19456
rect 23492 19400 23612 19428
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 22980 19332 23244 19360
rect 23308 19332 23397 19360
rect 22980 19320 22986 19332
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20855 19264 21005 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19292 22431 19295
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22419 19264 22569 19292
rect 22419 19261 22431 19264
rect 22373 19255 22431 19261
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 23216 19292 23244 19332
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 23290 19292 23296 19304
rect 23216 19264 23296 19292
rect 22557 19255 22615 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 23201 19227 23259 19233
rect 20088 19196 20852 19224
rect 20088 19156 20116 19196
rect 20824 19168 20852 19196
rect 23201 19193 23213 19227
rect 23247 19224 23259 19227
rect 23492 19224 23520 19400
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 23569 19363 23627 19369
rect 23569 19329 23581 19363
rect 23615 19360 23627 19363
rect 25498 19360 25504 19372
rect 23615 19332 25504 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 25498 19320 25504 19332
rect 25556 19320 25562 19372
rect 24397 19295 24455 19301
rect 24397 19261 24409 19295
rect 24443 19292 24455 19295
rect 25130 19292 25136 19304
rect 24443 19264 25136 19292
rect 24443 19261 24455 19264
rect 24397 19255 24455 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 23247 19196 23520 19224
rect 23247 19193 23259 19196
rect 23201 19187 23259 19193
rect 25498 19184 25504 19236
rect 25556 19224 25562 19236
rect 25608 19224 25636 19468
rect 25556 19196 25636 19224
rect 25556 19184 25562 19196
rect 16172 19128 20116 19156
rect 16172 19116 16178 19128
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 20625 19159 20683 19165
rect 20625 19156 20637 19159
rect 20312 19128 20637 19156
rect 20312 19116 20318 19128
rect 20625 19125 20637 19128
rect 20671 19125 20683 19159
rect 20625 19119 20683 19125
rect 20806 19116 20812 19168
rect 20864 19116 20870 19168
rect 21913 19159 21971 19165
rect 21913 19125 21925 19159
rect 21959 19156 21971 19159
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21959 19128 22201 19156
rect 21959 19125 21971 19128
rect 21913 19119 21971 19125
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 22189 19119 22247 19125
rect 23842 19116 23848 19168
rect 23900 19116 23906 19168
rect 1104 19066 24840 19088
rect 1104 19014 3917 19066
rect 3969 19014 3981 19066
rect 4033 19014 4045 19066
rect 4097 19014 4109 19066
rect 4161 19014 4173 19066
rect 4225 19014 9851 19066
rect 9903 19014 9915 19066
rect 9967 19014 9979 19066
rect 10031 19014 10043 19066
rect 10095 19014 10107 19066
rect 10159 19014 15785 19066
rect 15837 19014 15849 19066
rect 15901 19014 15913 19066
rect 15965 19014 15977 19066
rect 16029 19014 16041 19066
rect 16093 19014 21719 19066
rect 21771 19014 21783 19066
rect 21835 19014 21847 19066
rect 21899 19014 21911 19066
rect 21963 19014 21975 19066
rect 22027 19014 24840 19066
rect 1104 18992 24840 19014
rect 1394 18912 1400 18964
rect 1452 18912 1458 18964
rect 4522 18952 4528 18964
rect 3252 18924 4528 18952
rect 1412 18816 1440 18912
rect 3252 18893 3280 18924
rect 4522 18912 4528 18924
rect 4580 18912 4586 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7524 18924 8125 18952
rect 7524 18912 7530 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 12710 18952 12716 18964
rect 10560 18924 12716 18952
rect 10560 18912 10566 18924
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 16114 18912 16120 18964
rect 16172 18912 16178 18964
rect 16298 18912 16304 18964
rect 16356 18952 16362 18964
rect 17037 18955 17095 18961
rect 17037 18952 17049 18955
rect 16356 18924 17049 18952
rect 16356 18912 16362 18924
rect 17037 18921 17049 18924
rect 17083 18921 17095 18955
rect 17037 18915 17095 18921
rect 19705 18955 19763 18961
rect 19705 18921 19717 18955
rect 19751 18952 19763 18955
rect 20254 18952 20260 18964
rect 19751 18924 20260 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 20254 18912 20260 18924
rect 20312 18912 20318 18964
rect 20438 18912 20444 18964
rect 20496 18912 20502 18964
rect 21542 18912 21548 18964
rect 21600 18952 21606 18964
rect 21600 18924 22094 18952
rect 21600 18912 21606 18924
rect 3237 18887 3295 18893
rect 3237 18853 3249 18887
rect 3283 18853 3295 18887
rect 3237 18847 3295 18853
rect 4614 18844 4620 18896
rect 4672 18884 4678 18896
rect 5902 18884 5908 18896
rect 4672 18856 5908 18884
rect 4672 18844 4678 18856
rect 5902 18844 5908 18856
rect 5960 18844 5966 18896
rect 16132 18884 16160 18912
rect 16040 18856 16160 18884
rect 19981 18887 20039 18893
rect 9128 18828 9180 18834
rect 1578 18816 1584 18828
rect 1412 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 6730 18776 6736 18828
rect 6788 18816 6794 18828
rect 7101 18819 7159 18825
rect 7101 18816 7113 18819
rect 6788 18788 7113 18816
rect 6788 18776 6794 18788
rect 7101 18785 7113 18788
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 14458 18776 14464 18828
rect 14516 18776 14522 18828
rect 16040 18825 16068 18856
rect 19981 18853 19993 18887
rect 20027 18884 20039 18887
rect 20456 18884 20484 18912
rect 20027 18856 20484 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 19150 18776 19156 18828
rect 19208 18776 19214 18828
rect 22066 18816 22094 18924
rect 22833 18887 22891 18893
rect 22833 18853 22845 18887
rect 22879 18884 22891 18887
rect 23474 18884 23480 18896
rect 22879 18856 23480 18884
rect 22879 18853 22891 18856
rect 22833 18847 22891 18853
rect 23474 18844 23480 18856
rect 23532 18844 23538 18896
rect 23569 18887 23627 18893
rect 23569 18853 23581 18887
rect 23615 18884 23627 18887
rect 25130 18884 25136 18896
rect 23615 18856 25136 18884
rect 23615 18853 23627 18856
rect 23569 18847 23627 18853
rect 25130 18844 25136 18856
rect 25188 18844 25194 18896
rect 22066 18788 23888 18816
rect 9128 18770 9180 18776
rect 1855 18751 1913 18757
rect 1855 18717 1867 18751
rect 1901 18748 1913 18751
rect 2314 18748 2320 18760
rect 1901 18720 2320 18748
rect 1901 18717 1913 18720
rect 1855 18711 1913 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 3789 18751 3847 18757
rect 3789 18717 3801 18751
rect 3835 18717 3847 18751
rect 3789 18711 3847 18717
rect 1302 18640 1308 18692
rect 1360 18680 1366 18692
rect 3053 18683 3111 18689
rect 3053 18680 3065 18683
rect 1360 18652 3065 18680
rect 1360 18640 1366 18652
rect 3053 18649 3065 18652
rect 3099 18649 3111 18683
rect 3804 18680 3832 18711
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 4063 18751 4121 18757
rect 4063 18748 4075 18751
rect 4028 18720 4075 18748
rect 4028 18708 4034 18720
rect 4063 18717 4075 18720
rect 4109 18748 4121 18751
rect 4522 18748 4528 18760
rect 4109 18720 4528 18748
rect 4109 18717 4121 18720
rect 4063 18711 4121 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 4706 18708 4712 18760
rect 4764 18748 4770 18760
rect 6362 18748 6368 18760
rect 4764 18720 6368 18748
rect 4764 18708 4770 18720
rect 6362 18708 6368 18720
rect 6420 18748 6426 18760
rect 7343 18751 7401 18757
rect 7343 18748 7355 18751
rect 6420 18720 7355 18748
rect 6420 18708 6426 18720
rect 7343 18717 7355 18720
rect 7389 18717 7401 18751
rect 7343 18711 7401 18717
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9674 18748 9680 18760
rect 9539 18720 9680 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9824 18720 9873 18748
rect 9824 18708 9830 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 10243 18751 10301 18757
rect 10243 18748 10255 18751
rect 9861 18711 9919 18717
rect 9968 18720 10255 18748
rect 4540 18680 4568 18708
rect 9968 18692 9996 18720
rect 10243 18717 10255 18720
rect 10289 18748 10301 18751
rect 10410 18748 10416 18760
rect 10289 18720 10416 18748
rect 10289 18717 10301 18720
rect 10243 18711 10301 18717
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 11238 18708 11244 18760
rect 11296 18708 11302 18760
rect 11515 18751 11573 18757
rect 11515 18748 11527 18751
rect 11440 18720 11527 18748
rect 11440 18692 11468 18720
rect 11515 18717 11527 18720
rect 11561 18717 11573 18751
rect 14553 18751 14611 18757
rect 14553 18748 14565 18751
rect 11515 18711 11573 18717
rect 11624 18720 14565 18748
rect 7098 18680 7104 18692
rect 3804 18652 4108 18680
rect 4540 18652 7104 18680
rect 3053 18643 3111 18649
rect 4080 18624 4108 18652
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 7834 18640 7840 18692
rect 7892 18680 7898 18692
rect 9125 18683 9183 18689
rect 9125 18680 9137 18683
rect 7892 18652 9137 18680
rect 7892 18640 7898 18652
rect 9125 18649 9137 18652
rect 9171 18649 9183 18683
rect 9125 18643 9183 18649
rect 9950 18640 9956 18692
rect 10008 18640 10014 18692
rect 10870 18680 10876 18692
rect 10336 18652 10876 18680
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 2866 18612 2872 18624
rect 2639 18584 2872 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 4062 18572 4068 18624
rect 4120 18572 4126 18624
rect 4798 18572 4804 18624
rect 4856 18572 4862 18624
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 10336 18612 10364 18652
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 11422 18640 11428 18692
rect 11480 18640 11486 18692
rect 8720 18584 10364 18612
rect 8720 18572 8726 18584
rect 10410 18572 10416 18624
rect 10468 18572 10474 18624
rect 10888 18612 10916 18640
rect 11624 18612 11652 18720
rect 14553 18717 14565 18720
rect 14599 18748 14611 18751
rect 14918 18748 14924 18760
rect 14599 18720 14924 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 15010 18708 15016 18760
rect 15068 18708 15074 18760
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 16299 18751 16357 18757
rect 16299 18748 16311 18751
rect 16264 18720 16311 18748
rect 16264 18708 16270 18720
rect 16299 18717 16311 18720
rect 16345 18717 16357 18751
rect 16299 18711 16357 18717
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17184 18720 17601 18748
rect 17184 18708 17190 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 17831 18751 17889 18757
rect 17831 18748 17843 18751
rect 17589 18711 17647 18717
rect 17696 18720 17843 18748
rect 11992 18652 14228 18680
rect 11992 18624 12020 18652
rect 10888 18584 11652 18612
rect 11974 18572 11980 18624
rect 12032 18572 12038 18624
rect 12250 18572 12256 18624
rect 12308 18572 12314 18624
rect 14200 18612 14228 18652
rect 14274 18640 14280 18692
rect 14332 18640 14338 18692
rect 14642 18640 14648 18692
rect 14700 18640 14706 18692
rect 15746 18680 15752 18692
rect 15396 18652 15752 18680
rect 15396 18621 15424 18652
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 17696 18680 17724 18720
rect 17831 18717 17843 18720
rect 17877 18717 17889 18751
rect 19168 18748 19196 18776
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19168 18720 19625 18748
rect 17831 18711 17889 18717
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18748 20223 18751
rect 20622 18748 20628 18760
rect 20211 18720 20628 18748
rect 20211 18717 20223 18720
rect 20165 18711 20223 18717
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 22741 18751 22799 18757
rect 22741 18717 22753 18751
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 21174 18680 21180 18692
rect 16592 18652 21180 18680
rect 16592 18624 16620 18652
rect 21174 18640 21180 18652
rect 21232 18640 21238 18692
rect 22756 18680 22784 18711
rect 22922 18708 22928 18760
rect 22980 18708 22986 18760
rect 23106 18708 23112 18760
rect 23164 18748 23170 18760
rect 23201 18751 23259 18757
rect 23201 18748 23213 18751
rect 23164 18720 23213 18748
rect 23164 18708 23170 18720
rect 23201 18717 23213 18720
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23382 18708 23388 18760
rect 23440 18708 23446 18760
rect 23860 18757 23888 18788
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 23750 18680 23756 18692
rect 22756 18652 23756 18680
rect 23750 18640 23756 18652
rect 23808 18640 23814 18692
rect 15381 18615 15439 18621
rect 15381 18612 15393 18615
rect 14200 18584 15393 18612
rect 15381 18581 15393 18584
rect 15427 18581 15439 18615
rect 15381 18575 15439 18581
rect 15562 18572 15568 18624
rect 15620 18572 15626 18624
rect 16574 18572 16580 18624
rect 16632 18572 16638 18624
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18380 18584 18613 18612
rect 18380 18572 18386 18584
rect 18601 18581 18613 18584
rect 18647 18581 18659 18615
rect 18601 18575 18659 18581
rect 23014 18572 23020 18624
rect 23072 18572 23078 18624
rect 24121 18615 24179 18621
rect 24121 18581 24133 18615
rect 24167 18612 24179 18615
rect 25314 18612 25320 18624
rect 24167 18584 25320 18612
rect 24167 18581 24179 18584
rect 24121 18575 24179 18581
rect 25314 18572 25320 18584
rect 25372 18572 25378 18624
rect 1104 18522 25000 18544
rect 1104 18470 6884 18522
rect 6936 18470 6948 18522
rect 7000 18470 7012 18522
rect 7064 18470 7076 18522
rect 7128 18470 7140 18522
rect 7192 18470 12818 18522
rect 12870 18470 12882 18522
rect 12934 18470 12946 18522
rect 12998 18470 13010 18522
rect 13062 18470 13074 18522
rect 13126 18470 18752 18522
rect 18804 18470 18816 18522
rect 18868 18470 18880 18522
rect 18932 18470 18944 18522
rect 18996 18470 19008 18522
rect 19060 18470 24686 18522
rect 24738 18470 24750 18522
rect 24802 18470 24814 18522
rect 24866 18470 24878 18522
rect 24930 18470 24942 18522
rect 24994 18470 25000 18522
rect 1104 18448 25000 18470
rect 934 18368 940 18420
rect 992 18408 998 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 992 18380 5549 18408
rect 992 18368 998 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 5537 18371 5595 18377
rect 5626 18368 5632 18420
rect 5684 18408 5690 18420
rect 8294 18408 8300 18420
rect 5684 18380 8300 18408
rect 5684 18368 5690 18380
rect 1210 18300 1216 18352
rect 1268 18340 1274 18352
rect 3513 18343 3571 18349
rect 3513 18340 3525 18343
rect 1268 18312 3525 18340
rect 1268 18300 1274 18312
rect 3513 18309 3525 18312
rect 3559 18309 3571 18343
rect 3513 18303 3571 18309
rect 4062 18300 4068 18352
rect 4120 18300 4126 18352
rect 4706 18340 4712 18352
rect 4246 18312 4712 18340
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 1854 18232 1860 18284
rect 1912 18272 1918 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 1912 18244 2053 18272
rect 1912 18232 1918 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2314 18272 2320 18284
rect 2275 18244 2320 18272
rect 2041 18235 2099 18241
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 3973 18275 4031 18281
rect 3973 18241 3985 18275
rect 4019 18272 4031 18275
rect 4080 18272 4108 18300
rect 4019 18244 4108 18272
rect 4019 18241 4031 18244
rect 3973 18235 4031 18241
rect 4154 18232 4160 18284
rect 4212 18272 4218 18284
rect 4246 18281 4274 18312
rect 4706 18300 4712 18312
rect 4764 18300 4770 18352
rect 4246 18275 4305 18281
rect 4246 18272 4259 18275
rect 4212 18244 4259 18272
rect 4212 18232 4218 18244
rect 4247 18241 4259 18244
rect 4293 18241 4305 18275
rect 4247 18235 4305 18241
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 5445 18275 5503 18281
rect 4396 18244 5028 18272
rect 4396 18232 4402 18244
rect 5000 18216 5028 18244
rect 5445 18241 5457 18275
rect 5491 18272 5503 18275
rect 5626 18272 5632 18284
rect 5491 18244 5632 18272
rect 5491 18241 5503 18244
rect 5445 18235 5503 18241
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 7944 18272 7972 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 9122 18368 9128 18420
rect 9180 18408 9186 18420
rect 9217 18411 9275 18417
rect 9217 18408 9229 18411
rect 9180 18380 9229 18408
rect 9180 18368 9186 18380
rect 9217 18377 9229 18380
rect 9263 18377 9275 18411
rect 9217 18371 9275 18377
rect 11606 18368 11612 18420
rect 11664 18408 11670 18420
rect 11701 18411 11759 18417
rect 11701 18408 11713 18411
rect 11664 18380 11713 18408
rect 11664 18368 11670 18380
rect 11701 18377 11713 18380
rect 11747 18377 11759 18411
rect 11701 18371 11759 18377
rect 11808 18380 14596 18408
rect 8018 18300 8024 18352
rect 8076 18340 8082 18352
rect 8076 18312 8614 18340
rect 8076 18300 8082 18312
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 7944 18244 8217 18272
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8478 18272 8484 18284
rect 8439 18244 8484 18272
rect 8205 18235 8263 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 8586 18272 8614 18312
rect 8938 18300 8944 18352
rect 8996 18340 9002 18352
rect 11808 18340 11836 18380
rect 8996 18312 11836 18340
rect 12069 18343 12127 18349
rect 8996 18300 9002 18312
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12250 18340 12256 18352
rect 12115 18312 12256 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 12805 18343 12863 18349
rect 12805 18340 12817 18343
rect 12676 18312 12817 18340
rect 12676 18300 12682 18312
rect 12805 18309 12817 18312
rect 12851 18309 12863 18343
rect 14568 18340 14596 18380
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14700 18380 15209 18408
rect 14700 18368 14706 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15304 18380 18828 18408
rect 15304 18340 15332 18380
rect 14568 18312 15332 18340
rect 18800 18340 18828 18380
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21416 18380 24164 18408
rect 21416 18368 21422 18380
rect 22802 18343 22860 18349
rect 22802 18340 22814 18343
rect 18800 18312 22814 18340
rect 12805 18303 12863 18309
rect 22802 18309 22814 18312
rect 22848 18340 22860 18343
rect 23106 18340 23112 18352
rect 22848 18312 23112 18340
rect 22848 18309 22860 18312
rect 22802 18303 22860 18309
rect 23106 18300 23112 18312
rect 23164 18300 23170 18352
rect 24136 18349 24164 18380
rect 24121 18343 24179 18349
rect 24121 18309 24133 18343
rect 24167 18309 24179 18343
rect 24121 18303 24179 18309
rect 9859 18275 9917 18281
rect 9859 18272 9871 18275
rect 8586 18244 9871 18272
rect 9859 18241 9871 18244
rect 9905 18272 9917 18275
rect 10318 18272 10324 18284
rect 9905 18244 10324 18272
rect 9905 18241 9917 18244
rect 9859 18235 9917 18241
rect 10318 18232 10324 18244
rect 10376 18232 10382 18284
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 11379 18244 11989 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 11977 18241 11989 18244
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 12216 18244 12449 18272
rect 12216 18232 12222 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 14148 18244 14197 18272
rect 14148 18232 14154 18244
rect 14185 18241 14197 18244
rect 14231 18241 14243 18275
rect 14185 18235 14243 18241
rect 14459 18275 14517 18281
rect 14459 18241 14471 18275
rect 14505 18272 14517 18275
rect 14505 18244 15516 18272
rect 14505 18241 14517 18244
rect 14459 18235 14517 18241
rect 1578 18164 1584 18216
rect 1636 18164 1642 18216
rect 4982 18164 4988 18216
rect 5040 18164 5046 18216
rect 9582 18164 9588 18216
rect 9640 18164 9646 18216
rect 12526 18164 12532 18216
rect 12584 18164 12590 18216
rect 12894 18164 12900 18216
rect 12952 18164 12958 18216
rect 1596 18136 1624 18164
rect 11146 18136 11152 18148
rect 1504 18108 1624 18136
rect 4908 18108 8340 18136
rect 1504 18080 1532 18108
rect 1486 18028 1492 18080
rect 1544 18028 1550 18080
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 3016 18040 3065 18068
rect 3016 18028 3022 18040
rect 3053 18037 3065 18040
rect 3099 18037 3111 18071
rect 3053 18031 3111 18037
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 4908 18068 4936 18108
rect 3651 18040 4936 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4982 18028 4988 18080
rect 5040 18028 5046 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 6454 18068 6460 18080
rect 5592 18040 6460 18068
rect 5592 18028 5598 18040
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 8312 18068 8340 18108
rect 10428 18108 11152 18136
rect 10428 18068 10456 18108
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 12912 18136 12940 18164
rect 12989 18139 13047 18145
rect 12989 18136 13001 18139
rect 12912 18108 13001 18136
rect 12989 18105 13001 18108
rect 13035 18136 13047 18139
rect 13078 18136 13084 18148
rect 13035 18108 13084 18136
rect 13035 18105 13047 18108
rect 12989 18099 13047 18105
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 15488 18136 15516 18244
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 17175 18244 17448 18272
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 15764 18204 15792 18232
rect 17420 18216 17448 18244
rect 18322 18232 18328 18284
rect 18380 18232 18386 18284
rect 19242 18232 19248 18284
rect 19300 18232 19306 18284
rect 22370 18232 22376 18284
rect 22428 18272 22434 18284
rect 22557 18275 22615 18281
rect 22557 18272 22569 18275
rect 22428 18244 22569 18272
rect 22428 18232 22434 18244
rect 22557 18241 22569 18244
rect 22603 18241 22615 18275
rect 22557 18235 22615 18241
rect 23290 18232 23296 18284
rect 23348 18272 23354 18284
rect 23348 18244 24440 18272
rect 23348 18232 23354 18244
rect 17034 18204 17040 18216
rect 15764 18176 17040 18204
rect 17034 18164 17040 18176
rect 17092 18204 17098 18216
rect 17313 18207 17371 18213
rect 17313 18204 17325 18207
rect 17092 18176 17325 18204
rect 17092 18164 17098 18176
rect 17313 18173 17325 18176
rect 17359 18173 17371 18207
rect 17313 18167 17371 18173
rect 17402 18164 17408 18216
rect 17460 18164 17466 18216
rect 18046 18164 18052 18216
rect 18104 18164 18110 18216
rect 18187 18207 18245 18213
rect 18187 18173 18199 18207
rect 18233 18204 18245 18207
rect 19260 18204 19288 18232
rect 24412 18216 24440 18244
rect 18233 18176 19288 18204
rect 18233 18173 18245 18176
rect 18187 18167 18245 18173
rect 17678 18136 17684 18148
rect 15488 18108 17684 18136
rect 17678 18096 17684 18108
rect 17736 18096 17742 18148
rect 17773 18139 17831 18145
rect 17773 18105 17785 18139
rect 17819 18136 17831 18139
rect 17862 18136 17868 18148
rect 17819 18108 17868 18136
rect 17819 18105 17831 18108
rect 17773 18099 17831 18105
rect 17862 18096 17868 18108
rect 17920 18096 17926 18148
rect 8312 18040 10456 18068
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10560 18040 10609 18068
rect 10560 18028 10566 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 10686 18028 10692 18080
rect 10744 18068 10750 18080
rect 11698 18068 11704 18080
rect 10744 18040 11704 18068
rect 10744 18028 10750 18040
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 13722 18028 13728 18080
rect 13780 18068 13786 18080
rect 14550 18068 14556 18080
rect 13780 18040 14556 18068
rect 13780 18028 13786 18040
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 18708 18068 18736 18176
rect 24394 18164 24400 18216
rect 24452 18164 24458 18216
rect 16172 18040 18736 18068
rect 16172 18028 16178 18040
rect 18966 18028 18972 18080
rect 19024 18028 19030 18080
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 23937 18071 23995 18077
rect 23937 18068 23949 18071
rect 23624 18040 23949 18068
rect 23624 18028 23630 18040
rect 23937 18037 23949 18040
rect 23983 18037 23995 18071
rect 23937 18031 23995 18037
rect 24394 18028 24400 18080
rect 24452 18028 24458 18080
rect 1104 17978 24840 18000
rect 1104 17926 3917 17978
rect 3969 17926 3981 17978
rect 4033 17926 4045 17978
rect 4097 17926 4109 17978
rect 4161 17926 4173 17978
rect 4225 17926 9851 17978
rect 9903 17926 9915 17978
rect 9967 17926 9979 17978
rect 10031 17926 10043 17978
rect 10095 17926 10107 17978
rect 10159 17926 15785 17978
rect 15837 17926 15849 17978
rect 15901 17926 15913 17978
rect 15965 17926 15977 17978
rect 16029 17926 16041 17978
rect 16093 17926 21719 17978
rect 21771 17926 21783 17978
rect 21835 17926 21847 17978
rect 21899 17926 21911 17978
rect 21963 17926 21975 17978
rect 22027 17926 24840 17978
rect 1104 17904 24840 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 2130 17864 2136 17876
rect 1912 17836 2136 17864
rect 1912 17824 1918 17836
rect 2130 17824 2136 17836
rect 2188 17824 2194 17876
rect 2682 17864 2688 17876
rect 2424 17836 2688 17864
rect 2424 17805 2452 17836
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 4798 17864 4804 17876
rect 4448 17836 4804 17864
rect 4448 17805 4476 17836
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 10778 17864 10784 17876
rect 5736 17836 8524 17864
rect 2409 17799 2467 17805
rect 2409 17765 2421 17799
rect 2455 17765 2467 17799
rect 2409 17759 2467 17765
rect 4433 17799 4491 17805
rect 4433 17765 4445 17799
rect 4479 17765 4491 17799
rect 4433 17759 4491 17765
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 1995 17700 3648 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 3620 17672 3648 17700
rect 3786 17688 3792 17740
rect 3844 17688 3850 17740
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 3896 17700 4721 17728
rect 1394 17620 1400 17672
rect 1452 17620 1458 17672
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 2130 17660 2136 17672
rect 1811 17632 2136 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2682 17620 2688 17672
rect 2740 17620 2746 17672
rect 2774 17620 2780 17672
rect 2832 17669 2838 17672
rect 2832 17663 2860 17669
rect 2848 17629 2860 17663
rect 2832 17623 2860 17629
rect 2832 17620 2838 17623
rect 2958 17620 2964 17672
rect 3016 17620 3022 17672
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 3896 17660 3924 17700
rect 4709 17697 4721 17700
rect 4755 17697 4767 17731
rect 4709 17691 4767 17697
rect 4847 17731 4905 17737
rect 4847 17697 4859 17731
rect 4893 17728 4905 17731
rect 5736 17728 5764 17836
rect 4893 17700 5764 17728
rect 6773 17700 8432 17728
rect 4893 17697 4905 17700
rect 4847 17691 4905 17697
rect 3660 17632 3924 17660
rect 3973 17663 4031 17669
rect 3660 17620 3666 17632
rect 3973 17629 3985 17663
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 3988 17592 4016 17623
rect 4982 17620 4988 17672
rect 5040 17620 5046 17672
rect 5721 17663 5779 17669
rect 5721 17629 5733 17663
rect 5767 17629 5779 17663
rect 5721 17623 5779 17629
rect 5979 17633 6037 17639
rect 5736 17592 5764 17623
rect 5979 17599 5991 17633
rect 6025 17630 6037 17633
rect 6025 17599 6040 17630
rect 5979 17593 6040 17599
rect 6012 17592 6040 17593
rect 6362 17592 6368 17604
rect 3568 17564 4016 17592
rect 3568 17552 3574 17564
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 3234 17524 3240 17536
rect 1627 17496 3240 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 3234 17484 3240 17496
rect 3292 17484 3298 17536
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3476 17496 3617 17524
rect 3476 17484 3482 17496
rect 3605 17493 3617 17496
rect 3651 17493 3663 17527
rect 3988 17524 4016 17564
rect 5460 17564 5948 17592
rect 6012 17564 6368 17592
rect 4614 17524 4620 17536
rect 3988 17496 4620 17524
rect 3605 17487 3663 17493
rect 4614 17484 4620 17496
rect 4672 17484 4678 17536
rect 4798 17484 4804 17536
rect 4856 17524 4862 17536
rect 5460 17524 5488 17564
rect 4856 17496 5488 17524
rect 4856 17484 4862 17496
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5629 17527 5687 17533
rect 5629 17524 5641 17527
rect 5592 17496 5641 17524
rect 5592 17484 5598 17496
rect 5629 17493 5641 17496
rect 5675 17493 5687 17527
rect 5920 17524 5948 17564
rect 6362 17552 6368 17564
rect 6420 17552 6426 17604
rect 6773 17592 6801 17700
rect 8404 17672 8432 17700
rect 6914 17620 6920 17672
rect 6972 17620 6978 17672
rect 8386 17620 8392 17672
rect 8444 17620 8450 17672
rect 6472 17564 6801 17592
rect 6472 17524 6500 17564
rect 5920 17496 6500 17524
rect 5629 17487 5687 17493
rect 6730 17484 6736 17536
rect 6788 17484 6794 17536
rect 6932 17524 6960 17620
rect 8496 17592 8524 17836
rect 9784 17836 10784 17864
rect 9784 17740 9812 17836
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11112 17836 17816 17864
rect 11112 17824 11118 17836
rect 10413 17799 10471 17805
rect 10413 17765 10425 17799
rect 10459 17796 10471 17799
rect 10502 17796 10508 17808
rect 10459 17768 10508 17796
rect 10459 17765 10471 17768
rect 10413 17759 10471 17765
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 12250 17796 12256 17808
rect 12084 17768 12256 17796
rect 9766 17688 9772 17740
rect 9824 17688 9830 17740
rect 10806 17731 10864 17737
rect 10806 17728 10818 17731
rect 9876 17700 10818 17728
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 9876 17660 9904 17700
rect 10806 17697 10818 17700
rect 10852 17697 10864 17731
rect 10806 17691 10864 17697
rect 11146 17688 11152 17740
rect 11204 17728 11210 17740
rect 12084 17737 12112 17768
rect 12250 17756 12256 17768
rect 12308 17756 12314 17808
rect 12069 17731 12127 17737
rect 11204 17700 11836 17728
rect 11204 17688 11210 17700
rect 9364 17632 9904 17660
rect 9953 17663 10011 17669
rect 9364 17620 9370 17632
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 10134 17660 10140 17672
rect 9999 17632 10140 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 9968 17592 9996 17623
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10686 17620 10692 17672
rect 10744 17620 10750 17672
rect 10962 17620 10968 17672
rect 11020 17620 11026 17672
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17660 11667 17663
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11655 17632 11713 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11701 17623 11759 17629
rect 8496 17564 9996 17592
rect 11808 17592 11836 17700
rect 12069 17697 12081 17731
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 12158 17688 12164 17740
rect 12216 17728 12222 17740
rect 12216 17700 12434 17728
rect 12216 17688 12222 17700
rect 12406 17672 12434 17700
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 12989 17731 13047 17737
rect 12989 17697 13001 17731
rect 13035 17728 13047 17731
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13035 17700 14289 17728
rect 13035 17697 13047 17700
rect 12989 17691 13047 17697
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14366 17700 16344 17728
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12406 17632 12440 17672
rect 12253 17623 12311 17629
rect 12268 17592 12296 17623
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 13078 17620 13084 17672
rect 13136 17669 13142 17672
rect 13136 17663 13164 17669
rect 13152 17629 13164 17663
rect 13136 17623 13164 17629
rect 13136 17620 13142 17623
rect 13262 17620 13268 17672
rect 13320 17620 13326 17672
rect 13906 17620 13912 17672
rect 13964 17660 13970 17672
rect 14366 17660 14394 17700
rect 16316 17672 16344 17700
rect 17126 17688 17132 17740
rect 17184 17688 17190 17740
rect 13964 17632 14394 17660
rect 13964 17620 13970 17632
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15286 17660 15292 17672
rect 14884 17632 15292 17660
rect 14884 17620 14890 17632
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 17371 17663 17429 17669
rect 17371 17660 17383 17663
rect 16356 17632 17383 17660
rect 16356 17620 16362 17632
rect 17371 17629 17383 17632
rect 17417 17629 17429 17663
rect 17788 17660 17816 17836
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 18141 17867 18199 17873
rect 18141 17864 18153 17867
rect 17920 17836 18153 17864
rect 17920 17824 17926 17836
rect 18141 17833 18153 17836
rect 18187 17833 18199 17867
rect 22370 17864 22376 17876
rect 18141 17827 18199 17833
rect 20732 17836 22376 17864
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 18693 17799 18751 17805
rect 18693 17796 18705 17799
rect 18104 17768 18705 17796
rect 18104 17756 18110 17768
rect 18693 17765 18705 17768
rect 18739 17765 18751 17799
rect 18693 17759 18751 17765
rect 20732 17737 20760 17836
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 22830 17824 22836 17876
rect 22888 17824 22894 17876
rect 23750 17824 23756 17876
rect 23808 17824 23814 17876
rect 22186 17756 22192 17808
rect 22244 17796 22250 17808
rect 22848 17796 22876 17824
rect 22244 17768 22876 17796
rect 22244 17756 22250 17768
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17697 20775 17731
rect 20717 17691 20775 17697
rect 17788 17632 18184 17660
rect 17371 17623 17429 17629
rect 18046 17592 18052 17604
rect 11808 17564 12296 17592
rect 13832 17564 18052 17592
rect 11885 17527 11943 17533
rect 11885 17524 11897 17527
rect 6932 17496 11897 17524
rect 11885 17493 11897 17496
rect 11931 17493 11943 17527
rect 11885 17487 11943 17493
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 13832 17524 13860 17564
rect 18046 17552 18052 17564
rect 18104 17552 18110 17604
rect 12124 17496 13860 17524
rect 13909 17527 13967 17533
rect 12124 17484 12130 17496
rect 13909 17493 13921 17527
rect 13955 17524 13967 17527
rect 17862 17524 17868 17536
rect 13955 17496 17868 17524
rect 13955 17493 13967 17496
rect 13909 17487 13967 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18156 17524 18184 17632
rect 18966 17620 18972 17672
rect 19024 17620 19030 17672
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17660 19303 17663
rect 20732 17660 20760 17691
rect 22094 17688 22100 17740
rect 22152 17728 22158 17740
rect 22462 17728 22468 17740
rect 22152 17700 22468 17728
rect 22152 17688 22158 17700
rect 22462 17688 22468 17700
rect 22520 17728 22526 17740
rect 22741 17731 22799 17737
rect 22741 17728 22753 17731
rect 22520 17700 22753 17728
rect 22520 17688 22526 17700
rect 22741 17697 22753 17700
rect 22787 17697 22799 17731
rect 22741 17691 22799 17697
rect 19291 17632 20760 17660
rect 19291 17629 19303 17632
rect 19245 17623 19303 17629
rect 22186 17620 22192 17672
rect 22244 17620 22250 17672
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 22999 17633 23057 17639
rect 18984 17592 19012 17620
rect 19426 17592 19432 17604
rect 18984 17564 19432 17592
rect 19426 17552 19432 17564
rect 19484 17601 19490 17604
rect 19484 17595 19548 17601
rect 19484 17561 19502 17595
rect 19536 17561 19548 17595
rect 20898 17592 20904 17604
rect 19484 17555 19548 17561
rect 19628 17564 20904 17592
rect 19484 17552 19490 17555
rect 19628 17524 19656 17564
rect 20898 17552 20904 17564
rect 20956 17601 20962 17604
rect 20956 17595 21020 17601
rect 20956 17561 20974 17595
rect 21008 17561 21020 17595
rect 22664 17592 22692 17623
rect 22999 17599 23011 17633
rect 23045 17630 23057 17633
rect 23045 17599 23060 17630
rect 22999 17593 23060 17599
rect 20956 17555 21020 17561
rect 22112 17564 22692 17592
rect 23032 17592 23060 17593
rect 23106 17592 23112 17604
rect 23032 17564 23112 17592
rect 20956 17552 20962 17555
rect 18156 17496 19656 17524
rect 20622 17484 20628 17536
rect 20680 17484 20686 17536
rect 22112 17533 22140 17564
rect 22097 17527 22155 17533
rect 22097 17493 22109 17527
rect 22143 17493 22155 17527
rect 22097 17487 22155 17493
rect 22278 17484 22284 17536
rect 22336 17484 22342 17536
rect 22462 17484 22468 17536
rect 22520 17484 22526 17536
rect 22646 17484 22652 17536
rect 22704 17524 22710 17536
rect 23032 17524 23060 17564
rect 23106 17552 23112 17564
rect 23164 17552 23170 17604
rect 22704 17496 23060 17524
rect 22704 17484 22710 17496
rect 24486 17484 24492 17536
rect 24544 17524 24550 17536
rect 25038 17524 25044 17536
rect 24544 17496 25044 17524
rect 24544 17484 24550 17496
rect 25038 17484 25044 17496
rect 25096 17484 25102 17536
rect 1104 17434 25000 17456
rect 1104 17382 6884 17434
rect 6936 17382 6948 17434
rect 7000 17382 7012 17434
rect 7064 17382 7076 17434
rect 7128 17382 7140 17434
rect 7192 17382 12818 17434
rect 12870 17382 12882 17434
rect 12934 17382 12946 17434
rect 12998 17382 13010 17434
rect 13062 17382 13074 17434
rect 13126 17382 18752 17434
rect 18804 17382 18816 17434
rect 18868 17382 18880 17434
rect 18932 17382 18944 17434
rect 18996 17382 19008 17434
rect 19060 17382 24686 17434
rect 24738 17382 24750 17434
rect 24802 17382 24814 17434
rect 24866 17382 24878 17434
rect 24930 17382 24942 17434
rect 24994 17382 25000 17434
rect 1104 17360 25000 17382
rect 3326 17320 3332 17332
rect 1596 17292 3332 17320
rect 382 17212 388 17264
rect 440 17252 446 17264
rect 1026 17252 1032 17264
rect 440 17224 1032 17252
rect 440 17212 446 17224
rect 1026 17212 1032 17224
rect 1084 17212 1090 17264
rect 1596 17193 1624 17292
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 4522 17280 4528 17332
rect 4580 17280 4586 17332
rect 6730 17280 6736 17332
rect 6788 17320 6794 17332
rect 6914 17320 6920 17332
rect 6788 17292 6920 17320
rect 6788 17280 6794 17292
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7116 17292 7849 17320
rect 3418 17212 3424 17264
rect 3476 17252 3482 17264
rect 3513 17255 3571 17261
rect 3513 17252 3525 17255
rect 3476 17224 3525 17252
rect 3476 17212 3482 17224
rect 3513 17221 3525 17224
rect 3559 17221 3571 17255
rect 4540 17252 4568 17280
rect 5166 17252 5172 17264
rect 4540 17224 5172 17252
rect 3513 17215 3571 17221
rect 5150 17217 5172 17224
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 2866 17144 2872 17196
rect 2924 17144 2930 17196
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 4798 17144 4804 17196
rect 4856 17184 4862 17196
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4856 17156 4905 17184
rect 4856 17144 4862 17156
rect 4893 17153 4905 17156
rect 4939 17153 4951 17187
rect 5150 17186 5163 17217
rect 5224 17212 5230 17264
rect 6549 17255 6607 17261
rect 6549 17221 6561 17255
rect 6595 17252 6607 17255
rect 6638 17252 6644 17264
rect 6595 17224 6644 17252
rect 6595 17221 6607 17224
rect 6549 17215 6607 17221
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 7116 17252 7144 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 8297 17323 8355 17329
rect 8297 17289 8309 17323
rect 8343 17320 8355 17323
rect 9122 17320 9128 17332
rect 8343 17292 9128 17320
rect 8343 17289 8355 17292
rect 8297 17283 8355 17289
rect 7653 17255 7711 17261
rect 7653 17252 7665 17255
rect 6748 17224 7144 17252
rect 7208 17224 7665 17252
rect 5151 17183 5163 17186
rect 5197 17183 5209 17212
rect 6748 17184 6776 17224
rect 7208 17196 7236 17224
rect 7653 17221 7665 17224
rect 7699 17221 7711 17255
rect 7653 17215 7711 17221
rect 7852 17196 7880 17283
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 10778 17320 10784 17332
rect 9824 17292 10784 17320
rect 9824 17280 9830 17292
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 11020 17292 11069 17320
rect 11020 17280 11026 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 12802 17320 12808 17332
rect 11057 17283 11115 17289
rect 12544 17292 12808 17320
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 8168 17224 8294 17252
rect 8168 17212 8174 17224
rect 5151 17177 5209 17183
rect 4893 17147 4951 17153
rect 6196 17156 6776 17184
rect 6196 17128 6224 17156
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 6914 17144 6920 17196
rect 6972 17144 6978 17196
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7331 17156 7696 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7668 17128 7696 17156
rect 7834 17144 7840 17196
rect 7892 17144 7898 17196
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17116 1915 17119
rect 2038 17116 2044 17128
rect 1903 17088 2044 17116
rect 1903 17085 1915 17088
rect 1857 17079 1915 17085
rect 1688 17048 1716 17079
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 2406 17116 2412 17128
rect 2363 17088 2412 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 2590 17076 2596 17128
rect 2648 17076 2654 17128
rect 2731 17119 2789 17125
rect 2731 17085 2743 17119
rect 2777 17116 2789 17119
rect 4338 17116 4344 17128
rect 2777 17088 4344 17116
rect 2777 17085 2789 17088
rect 2731 17079 2789 17085
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 6178 17076 6184 17128
rect 6236 17076 6242 17128
rect 2130 17048 2136 17060
rect 1688 17020 2136 17048
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 3605 17051 3663 17057
rect 3605 17017 3617 17051
rect 3651 17048 3663 17051
rect 3694 17048 3700 17060
rect 3651 17020 3700 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17048 5963 17051
rect 6380 17048 6408 17102
rect 7650 17076 7656 17128
rect 7708 17076 7714 17128
rect 5951 17020 6408 17048
rect 8266 17048 8294 17224
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 12544 17252 12572 17292
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 13262 17280 13268 17332
rect 13320 17320 13326 17332
rect 13633 17323 13691 17329
rect 13633 17320 13645 17323
rect 13320 17292 13645 17320
rect 13320 17280 13326 17292
rect 13633 17289 13645 17292
rect 13679 17289 13691 17323
rect 13633 17283 13691 17289
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 17034 17320 17040 17332
rect 14424 17292 17040 17320
rect 14424 17280 14430 17292
rect 17034 17280 17040 17292
rect 17092 17280 17098 17332
rect 17862 17280 17868 17332
rect 17920 17280 17926 17332
rect 19426 17280 19432 17332
rect 19484 17280 19490 17332
rect 19521 17323 19579 17329
rect 19521 17289 19533 17323
rect 19567 17289 19579 17323
rect 19521 17283 19579 17289
rect 17126 17252 17132 17264
rect 10652 17224 12572 17252
rect 12636 17224 17132 17252
rect 10652 17212 10658 17224
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 9582 17184 9588 17196
rect 9272 17156 9588 17184
rect 9272 17144 9278 17156
rect 9582 17144 9588 17156
rect 9640 17184 9646 17196
rect 10033 17187 10091 17193
rect 10033 17184 10045 17187
rect 9640 17156 10045 17184
rect 9640 17144 9646 17156
rect 10033 17153 10045 17156
rect 10079 17153 10091 17187
rect 10033 17147 10091 17153
rect 10318 17144 10324 17196
rect 10376 17184 10382 17196
rect 10376 17156 10419 17184
rect 10376 17144 10382 17156
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 12250 17184 12256 17196
rect 11112 17156 12256 17184
rect 11112 17144 11118 17156
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 12636 17193 12664 17224
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 12066 17116 12072 17128
rect 11756 17088 12072 17116
rect 11756 17076 11762 17088
rect 12066 17076 12072 17088
rect 12124 17116 12130 17128
rect 12636 17116 12664 17147
rect 12802 17144 12808 17196
rect 12860 17184 12866 17196
rect 12895 17187 12953 17193
rect 12895 17184 12907 17187
rect 12860 17156 12907 17184
rect 12860 17144 12866 17156
rect 12895 17153 12907 17156
rect 12941 17184 12953 17187
rect 13446 17184 13452 17196
rect 12941 17156 13452 17184
rect 12941 17153 12953 17156
rect 12895 17147 12953 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15439 17187 15497 17193
rect 15439 17184 15451 17187
rect 15068 17156 15451 17184
rect 15068 17144 15074 17156
rect 15439 17153 15451 17156
rect 15485 17184 15497 17187
rect 16298 17184 16304 17196
rect 15485 17156 16304 17184
rect 15485 17153 15497 17156
rect 15439 17147 15497 17153
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 16850 17184 16856 17196
rect 16684 17156 16856 17184
rect 12124 17088 12664 17116
rect 12124 17076 12130 17088
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 16684 17125 16712 17156
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 16943 17187 17001 17193
rect 16943 17153 16955 17187
rect 16989 17184 17001 17187
rect 17034 17184 17040 17196
rect 16989 17156 17040 17184
rect 16989 17153 17001 17156
rect 16943 17147 17001 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 15197 17119 15255 17125
rect 15197 17116 15209 17119
rect 14148 17088 15209 17116
rect 14148 17076 14154 17088
rect 15197 17085 15209 17088
rect 15243 17085 15255 17119
rect 15197 17079 15255 17085
rect 16669 17119 16727 17125
rect 16669 17085 16681 17119
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 9582 17048 9588 17060
rect 8266 17020 9588 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 9582 17008 9588 17020
rect 9640 17008 9646 17060
rect 1397 16983 1455 16989
rect 1397 16949 1409 16983
rect 1443 16980 1455 16983
rect 2590 16980 2596 16992
rect 1443 16952 2596 16980
rect 1443 16949 1455 16952
rect 1397 16943 1455 16949
rect 2590 16940 2596 16952
rect 2648 16940 2654 16992
rect 2682 16940 2688 16992
rect 2740 16980 2746 16992
rect 6178 16980 6184 16992
rect 2740 16952 6184 16980
rect 2740 16940 2746 16952
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 8386 16940 8392 16992
rect 8444 16980 8450 16992
rect 11238 16980 11244 16992
rect 8444 16952 11244 16980
rect 8444 16940 8450 16952
rect 11238 16940 11244 16952
rect 11296 16940 11302 16992
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12526 16980 12532 16992
rect 12483 16952 12532 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12526 16940 12532 16952
rect 12584 16940 12590 16992
rect 14458 16940 14464 16992
rect 14516 16940 14522 16992
rect 15212 16980 15240 17079
rect 16684 17048 16712 17079
rect 17678 17076 17684 17128
rect 17736 17076 17742 17128
rect 17880 17116 17908 17280
rect 19444 17184 19472 17280
rect 19536 17252 19564 17283
rect 20438 17280 20444 17332
rect 20496 17320 20502 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 20496 17292 20545 17320
rect 20496 17280 20502 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20533 17283 20591 17289
rect 20622 17280 20628 17332
rect 20680 17280 20686 17332
rect 20898 17280 20904 17332
rect 20956 17280 20962 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 22186 17320 22192 17332
rect 21039 17292 22192 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22462 17280 22468 17332
rect 22520 17280 22526 17332
rect 23014 17280 23020 17332
rect 23072 17280 23078 17332
rect 23569 17323 23627 17329
rect 23569 17289 23581 17323
rect 23615 17320 23627 17323
rect 25130 17320 25136 17332
rect 23615 17292 25136 17320
rect 23615 17289 23627 17292
rect 23569 17283 23627 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 19536 17224 20116 17252
rect 20088 17193 20116 17224
rect 19705 17187 19763 17193
rect 19705 17184 19717 17187
rect 19444 17156 19717 17184
rect 19705 17153 19717 17156
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20530 17144 20536 17196
rect 20588 17144 20594 17196
rect 20640 17184 20668 17280
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20640 17156 20729 17184
rect 20717 17153 20729 17156
rect 20763 17153 20775 17187
rect 20916 17184 20944 17280
rect 22480 17252 22508 17280
rect 21284 17224 21579 17252
rect 21177 17187 21235 17193
rect 21177 17184 21189 17187
rect 20916 17156 21189 17184
rect 20717 17147 20775 17153
rect 21177 17153 21189 17156
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 20346 17116 20352 17128
rect 17880 17088 20352 17116
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 20548 17116 20576 17144
rect 21284 17116 21312 17224
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17153 21511 17187
rect 21453 17147 21511 17153
rect 20548 17088 21312 17116
rect 15856 17020 16712 17048
rect 17696 17048 17724 17076
rect 21468 17048 21496 17147
rect 21551 17116 21579 17224
rect 21652 17224 22508 17252
rect 23032 17252 23060 17280
rect 23032 17224 24348 17252
rect 21652 17193 21680 17224
rect 21637 17187 21695 17193
rect 21637 17153 21649 17187
rect 21683 17153 21695 17187
rect 22063 17187 22121 17193
rect 22063 17184 22075 17187
rect 21637 17147 21695 17153
rect 21744 17156 22075 17184
rect 21744 17116 21772 17156
rect 22063 17153 22075 17156
rect 22109 17153 22121 17187
rect 22063 17147 22121 17153
rect 22830 17144 22836 17196
rect 22888 17184 22894 17196
rect 23385 17187 23443 17193
rect 23385 17184 23397 17187
rect 22888 17156 23397 17184
rect 22888 17144 22894 17156
rect 23385 17153 23397 17156
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23842 17144 23848 17196
rect 23900 17144 23906 17196
rect 24320 17193 24348 17224
rect 24305 17187 24363 17193
rect 24305 17153 24317 17187
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 21551 17088 21772 17116
rect 21818 17076 21824 17128
rect 21876 17076 21882 17128
rect 21634 17048 21640 17060
rect 17696 17020 18276 17048
rect 21468 17020 21640 17048
rect 15856 16980 15884 17020
rect 18248 16992 18276 17020
rect 21634 17008 21640 17020
rect 21692 17048 21698 17060
rect 21692 17020 21956 17048
rect 21692 17008 21698 17020
rect 15212 16952 15884 16980
rect 16206 16940 16212 16992
rect 16264 16940 16270 16992
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 18230 16940 18236 16992
rect 18288 16940 18294 16992
rect 20162 16940 20168 16992
rect 20220 16940 20226 16992
rect 21542 16940 21548 16992
rect 21600 16940 21606 16992
rect 21928 16980 21956 17020
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 21928 16952 22845 16980
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 24118 16940 24124 16992
rect 24176 16940 24182 16992
rect 24394 16940 24400 16992
rect 24452 16940 24458 16992
rect 1104 16890 24840 16912
rect 1104 16838 3917 16890
rect 3969 16838 3981 16890
rect 4033 16838 4045 16890
rect 4097 16838 4109 16890
rect 4161 16838 4173 16890
rect 4225 16838 9851 16890
rect 9903 16838 9915 16890
rect 9967 16838 9979 16890
rect 10031 16838 10043 16890
rect 10095 16838 10107 16890
rect 10159 16838 15785 16890
rect 15837 16838 15849 16890
rect 15901 16838 15913 16890
rect 15965 16838 15977 16890
rect 16029 16838 16041 16890
rect 16093 16838 21719 16890
rect 21771 16838 21783 16890
rect 21835 16838 21847 16890
rect 21899 16838 21911 16890
rect 21963 16838 21975 16890
rect 22027 16838 24840 16890
rect 1104 16816 24840 16838
rect 382 16736 388 16788
rect 440 16776 446 16788
rect 3510 16776 3516 16788
rect 440 16748 3516 16776
rect 440 16736 446 16748
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 3786 16736 3792 16788
rect 3844 16776 3850 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 3844 16748 8769 16776
rect 3844 16736 3850 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 10318 16776 10324 16788
rect 9640 16748 10324 16776
rect 9640 16736 9646 16748
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 11238 16736 11244 16788
rect 11296 16776 11302 16788
rect 13354 16776 13360 16788
rect 11296 16748 13360 16776
rect 11296 16736 11302 16748
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 6822 16708 6828 16720
rect 3292 16680 6828 16708
rect 3292 16668 3298 16680
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 7558 16668 7564 16720
rect 7616 16668 7622 16720
rect 1670 16600 1676 16652
rect 1728 16640 1734 16652
rect 1765 16643 1823 16649
rect 1765 16640 1777 16643
rect 1728 16612 1777 16640
rect 1728 16600 1734 16612
rect 1765 16609 1777 16612
rect 1811 16609 1823 16643
rect 1765 16603 1823 16609
rect 2041 16643 2099 16649
rect 2041 16609 2053 16643
rect 2087 16640 2099 16643
rect 2222 16640 2228 16652
rect 2087 16612 2228 16640
rect 2087 16609 2099 16612
rect 2041 16603 2099 16609
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 3142 16600 3148 16652
rect 3200 16640 3206 16652
rect 4522 16640 4528 16652
rect 3200 16612 4528 16640
rect 3200 16600 3206 16612
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 5902 16600 5908 16652
rect 5960 16600 5966 16652
rect 6362 16600 6368 16652
rect 6420 16640 6426 16652
rect 6730 16640 6736 16652
rect 6420 16612 6736 16640
rect 6420 16600 6426 16612
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 7006 16640 7012 16652
rect 6963 16612 7012 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16640 7159 16643
rect 7190 16640 7196 16652
rect 7147 16612 7196 16640
rect 7147 16609 7159 16612
rect 7101 16603 7159 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7300 16612 7997 16640
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 1578 16572 1584 16584
rect 1443 16544 1584 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 1578 16532 1584 16544
rect 1636 16532 1642 16584
rect 3510 16572 3516 16584
rect 2148 16544 3516 16572
rect 2148 16504 2176 16544
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 5350 16572 5356 16584
rect 3651 16544 5356 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 5920 16572 5948 16600
rect 6638 16572 6644 16584
rect 5920 16544 6644 16572
rect 6638 16532 6644 16544
rect 6696 16572 6702 16584
rect 7300 16572 7328 16612
rect 6696 16544 7328 16572
rect 6696 16532 6702 16544
rect 7834 16532 7840 16584
rect 7892 16532 7898 16584
rect 7969 16581 7997 16612
rect 8110 16600 8116 16652
rect 8168 16600 8174 16652
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 11974 16640 11980 16652
rect 8720 16612 11980 16640
rect 8720 16600 8726 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12636 16649 12664 16748
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 15565 16779 15623 16785
rect 15565 16745 15577 16779
rect 15611 16776 15623 16779
rect 16114 16776 16120 16788
rect 15611 16748 16120 16776
rect 15611 16745 15623 16748
rect 15565 16739 15623 16745
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 16206 16736 16212 16788
rect 16264 16736 16270 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16758 16776 16764 16788
rect 16356 16748 16764 16776
rect 16356 16736 16362 16748
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 17310 16776 17316 16788
rect 16908 16748 17316 16776
rect 16908 16736 16914 16748
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17678 16736 17684 16788
rect 17736 16736 17742 16788
rect 20162 16736 20168 16788
rect 20220 16776 20226 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 20220 16748 21281 16776
rect 20220 16736 20226 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 21542 16736 21548 16788
rect 21600 16736 21606 16788
rect 22005 16779 22063 16785
rect 22005 16745 22017 16779
rect 22051 16776 22063 16779
rect 22278 16776 22284 16788
rect 22051 16748 22284 16776
rect 22051 16745 22063 16748
rect 22005 16739 22063 16745
rect 22278 16736 22284 16748
rect 22336 16736 22342 16788
rect 13633 16711 13691 16717
rect 13633 16677 13645 16711
rect 13679 16677 13691 16711
rect 16224 16708 16252 16736
rect 16393 16711 16451 16717
rect 16393 16708 16405 16711
rect 16224 16680 16405 16708
rect 13633 16671 13691 16677
rect 16393 16677 16405 16680
rect 16439 16677 16451 16711
rect 16393 16671 16451 16677
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16609 12679 16643
rect 13648 16640 13676 16671
rect 13648 16612 14122 16640
rect 12621 16603 12679 16609
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 15712 16612 15976 16640
rect 15712 16600 15718 16612
rect 7969 16575 8033 16581
rect 7969 16544 7987 16575
rect 7975 16541 7987 16544
rect 8021 16541 8033 16575
rect 7975 16535 8033 16541
rect 12895 16575 12953 16581
rect 12895 16541 12907 16575
rect 12941 16572 12953 16575
rect 13630 16572 13636 16584
rect 12941 16544 13636 16572
rect 12941 16541 12953 16544
rect 12895 16535 12953 16541
rect 13188 16516 13216 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14516 16544 14565 16572
rect 14516 16532 14522 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15948 16581 15976 16612
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16080 16612 16712 16640
rect 16080 16600 16086 16612
rect 16684 16581 16712 16612
rect 16758 16600 16764 16652
rect 16816 16649 16822 16652
rect 16816 16643 16844 16649
rect 16832 16609 16844 16643
rect 16816 16603 16844 16609
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 17696 16640 17724 16736
rect 16991 16612 17724 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 16816 16600 16822 16603
rect 19610 16600 19616 16652
rect 19668 16640 19674 16652
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19668 16612 19809 16640
rect 19668 16600 19674 16612
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 21450 16600 21456 16652
rect 21508 16600 21514 16652
rect 21560 16640 21588 16736
rect 22097 16711 22155 16717
rect 22097 16677 22109 16711
rect 22143 16708 22155 16711
rect 22143 16680 23704 16708
rect 22143 16677 22155 16680
rect 22097 16671 22155 16677
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 21560 16612 22201 16640
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 22296 16612 23428 16640
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 15620 16544 15761 16572
rect 15620 16532 15626 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15933 16575 15991 16581
rect 15933 16541 15945 16575
rect 15979 16541 15991 16575
rect 15933 16535 15991 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 17681 16575 17739 16581
rect 17681 16572 17693 16575
rect 17635 16544 17693 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17681 16541 17693 16544
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 18230 16532 18236 16584
rect 18288 16572 18294 16584
rect 21177 16575 21235 16581
rect 18288 16551 20098 16572
rect 18288 16545 20113 16551
rect 18288 16544 20067 16545
rect 18288 16532 18294 16544
rect 1596 16476 2176 16504
rect 1596 16445 1624 16476
rect 2222 16464 2228 16516
rect 2280 16504 2286 16516
rect 2961 16507 3019 16513
rect 2961 16504 2973 16507
rect 2280 16476 2973 16504
rect 2280 16464 2286 16476
rect 2961 16473 2973 16476
rect 3007 16473 3019 16507
rect 3881 16507 3939 16513
rect 3881 16504 3893 16507
rect 2961 16467 3019 16473
rect 3436 16476 3893 16504
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 3050 16396 3056 16448
rect 3108 16396 3114 16448
rect 3436 16445 3464 16476
rect 3881 16473 3893 16476
rect 3927 16473 3939 16507
rect 3881 16467 3939 16473
rect 4614 16464 4620 16516
rect 4672 16504 4678 16516
rect 5258 16504 5264 16516
rect 4672 16476 5264 16504
rect 4672 16464 4678 16476
rect 5258 16464 5264 16476
rect 5316 16464 5322 16516
rect 13170 16464 13176 16516
rect 13228 16464 13234 16516
rect 13998 16464 14004 16516
rect 14056 16504 14062 16516
rect 14277 16507 14335 16513
rect 14277 16504 14289 16507
rect 14056 16476 14289 16504
rect 14056 16464 14062 16476
rect 14277 16473 14289 16476
rect 14323 16473 14335 16507
rect 14277 16467 14335 16473
rect 14645 16507 14703 16513
rect 14645 16473 14657 16507
rect 14691 16504 14703 16507
rect 14918 16504 14924 16516
rect 14691 16476 14924 16504
rect 14691 16473 14703 16476
rect 14645 16467 14703 16473
rect 14918 16464 14924 16476
rect 14976 16464 14982 16516
rect 15013 16507 15071 16513
rect 15013 16473 15025 16507
rect 15059 16504 15071 16507
rect 20055 16511 20067 16544
rect 20101 16511 20113 16545
rect 21177 16541 21189 16575
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 20055 16505 20113 16511
rect 15059 16476 15976 16504
rect 15059 16473 15071 16476
rect 15013 16467 15071 16473
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 3970 16396 3976 16448
rect 4028 16396 4034 16448
rect 4982 16396 4988 16448
rect 5040 16436 5046 16448
rect 6270 16436 6276 16448
rect 5040 16408 6276 16436
rect 5040 16396 5046 16408
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 12250 16436 12256 16448
rect 8444 16408 12256 16436
rect 8444 16396 8450 16408
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 15378 16396 15384 16448
rect 15436 16396 15442 16448
rect 15948 16436 15976 16476
rect 17402 16436 17408 16448
rect 15948 16408 17408 16436
rect 17402 16396 17408 16408
rect 17460 16396 17466 16448
rect 17862 16396 17868 16448
rect 17920 16396 17926 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 20809 16439 20867 16445
rect 20809 16436 20821 16439
rect 20772 16408 20821 16436
rect 20772 16396 20778 16408
rect 20809 16405 20821 16408
rect 20855 16436 20867 16439
rect 21192 16436 21220 16535
rect 21634 16532 21640 16584
rect 21692 16572 21698 16584
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 21692 16544 21925 16572
rect 21692 16532 21698 16544
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 21913 16535 21971 16541
rect 21453 16507 21511 16513
rect 21453 16473 21465 16507
rect 21499 16504 21511 16507
rect 22296 16504 22324 16612
rect 22922 16532 22928 16584
rect 22980 16532 22986 16584
rect 21499 16476 22324 16504
rect 21499 16473 21511 16476
rect 21453 16467 21511 16473
rect 20855 16408 21220 16436
rect 22940 16436 22968 16532
rect 23400 16504 23428 16612
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16572 23535 16575
rect 23566 16572 23572 16584
rect 23523 16544 23572 16572
rect 23523 16541 23535 16544
rect 23477 16535 23535 16541
rect 23566 16532 23572 16544
rect 23624 16532 23630 16584
rect 23676 16581 23704 16680
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 24029 16507 24087 16513
rect 23400 16476 23704 16504
rect 23676 16448 23704 16476
rect 24029 16473 24041 16507
rect 24075 16504 24087 16507
rect 25222 16504 25228 16516
rect 24075 16476 25228 16504
rect 24075 16473 24087 16476
rect 24029 16467 24087 16473
rect 25222 16464 25228 16476
rect 25280 16464 25286 16516
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22940 16408 23305 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 23658 16396 23664 16448
rect 23716 16396 23722 16448
rect 566 16328 572 16380
rect 624 16328 630 16380
rect 1104 16346 25000 16368
rect 584 16176 612 16328
rect 1104 16294 6884 16346
rect 6936 16294 6948 16346
rect 7000 16294 7012 16346
rect 7064 16294 7076 16346
rect 7128 16294 7140 16346
rect 7192 16294 12818 16346
rect 12870 16294 12882 16346
rect 12934 16294 12946 16346
rect 12998 16294 13010 16346
rect 13062 16294 13074 16346
rect 13126 16294 18752 16346
rect 18804 16294 18816 16346
rect 18868 16294 18880 16346
rect 18932 16294 18944 16346
rect 18996 16294 19008 16346
rect 19060 16294 24686 16346
rect 24738 16294 24750 16346
rect 24802 16294 24814 16346
rect 24866 16294 24878 16346
rect 24930 16294 24942 16346
rect 24994 16294 25000 16346
rect 1104 16272 25000 16294
rect 1688 16204 7604 16232
rect 566 16124 572 16176
rect 624 16124 630 16176
rect 1688 16173 1716 16204
rect 1673 16167 1731 16173
rect 1673 16133 1685 16167
rect 1719 16133 1731 16167
rect 1673 16127 1731 16133
rect 2038 16124 2044 16176
rect 2096 16124 2102 16176
rect 3326 16164 3332 16176
rect 2424 16136 3332 16164
rect 2424 16135 2452 16136
rect 2391 16129 2452 16135
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 2133 16099 2191 16105
rect 2133 16096 2145 16099
rect 1912 16068 2145 16096
rect 1912 16056 1918 16068
rect 2133 16065 2145 16068
rect 2179 16065 2191 16099
rect 2391 16095 2403 16129
rect 2437 16098 2452 16129
rect 3326 16124 3332 16136
rect 3384 16124 3390 16176
rect 5350 16124 5356 16176
rect 5408 16124 5414 16176
rect 6270 16124 6276 16176
rect 6328 16124 6334 16176
rect 7576 16164 7604 16204
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8481 16235 8539 16241
rect 8481 16232 8493 16235
rect 8168 16204 8493 16232
rect 8168 16192 8174 16204
rect 8481 16201 8493 16204
rect 8527 16201 8539 16235
rect 8481 16195 8539 16201
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13081 16235 13139 16241
rect 13081 16232 13093 16235
rect 12768 16204 13093 16232
rect 12768 16192 12774 16204
rect 13081 16201 13093 16204
rect 13127 16201 13139 16235
rect 13081 16195 13139 16201
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 15381 16235 15439 16241
rect 15381 16232 15393 16235
rect 14976 16204 15393 16232
rect 14976 16192 14982 16204
rect 15381 16201 15393 16204
rect 15427 16201 15439 16235
rect 15381 16195 15439 16201
rect 17862 16192 17868 16244
rect 17920 16192 17926 16244
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16201 19303 16235
rect 19245 16195 19303 16201
rect 17880 16164 17908 16192
rect 18138 16173 18144 16176
rect 18132 16164 18144 16173
rect 7576 16136 17908 16164
rect 18099 16136 18144 16164
rect 18132 16127 18144 16136
rect 18138 16124 18144 16127
rect 18196 16124 18202 16176
rect 19260 16164 19288 16195
rect 20438 16192 20444 16244
rect 20496 16192 20502 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21450 16232 21456 16244
rect 20855 16204 21456 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 21542 16192 21548 16244
rect 21600 16232 21606 16244
rect 23290 16232 23296 16244
rect 21600 16204 23296 16232
rect 21600 16192 21606 16204
rect 23290 16192 23296 16204
rect 23348 16192 23354 16244
rect 23750 16192 23756 16244
rect 23808 16192 23814 16244
rect 23842 16192 23848 16244
rect 23900 16232 23906 16244
rect 24305 16235 24363 16241
rect 24305 16232 24317 16235
rect 23900 16204 24317 16232
rect 23900 16192 23906 16204
rect 24305 16201 24317 16204
rect 24351 16201 24363 16235
rect 24305 16195 24363 16201
rect 20456 16164 20484 16192
rect 19260 16136 19840 16164
rect 20456 16136 20852 16164
rect 2437 16095 2449 16098
rect 2391 16089 2449 16095
rect 2133 16059 2191 16065
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 3513 16099 3571 16105
rect 3513 16096 3525 16099
rect 2832 16068 3525 16096
rect 2832 16056 2838 16068
rect 3513 16065 3525 16068
rect 3559 16065 3571 16099
rect 3513 16059 3571 16065
rect 4430 16056 4436 16108
rect 4488 16056 4494 16108
rect 6288 16096 6316 16124
rect 7711 16099 7769 16105
rect 7711 16096 7723 16099
rect 6288 16068 7723 16096
rect 7711 16065 7723 16068
rect 7757 16065 7769 16099
rect 7711 16059 7769 16065
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 9030 16096 9036 16108
rect 8895 16068 9036 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9123 16099 9181 16105
rect 9123 16065 9135 16099
rect 9169 16096 9181 16099
rect 9169 16068 10548 16096
rect 9169 16065 9181 16068
rect 9123 16059 9181 16065
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 4614 16037 4620 16040
rect 3697 16031 3755 16037
rect 3697 16028 3709 16031
rect 3660 16000 3709 16028
rect 3660 15988 3666 16000
rect 3697 15997 3709 16000
rect 3743 15997 3755 16031
rect 3697 15991 3755 15997
rect 4571 16031 4620 16037
rect 4571 15997 4583 16031
rect 4617 15997 4620 16031
rect 4571 15991 4620 15997
rect 4614 15988 4620 15991
rect 4672 15988 4678 16040
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 4890 15988 4896 16040
rect 4948 16028 4954 16040
rect 6270 16028 6276 16040
rect 4948 16000 6276 16028
rect 4948 15988 4954 16000
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7340 16000 7481 16028
rect 7340 15988 7346 16000
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 9674 16028 9680 16040
rect 7469 15991 7527 15997
rect 9600 16000 9680 16028
rect 3145 15963 3203 15969
rect 3145 15929 3157 15963
rect 3191 15960 3203 15963
rect 4157 15963 4215 15969
rect 4157 15960 4169 15963
rect 3191 15932 4169 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 4157 15929 4169 15932
rect 4203 15929 4215 15963
rect 4157 15923 4215 15929
rect 5092 15932 7604 15960
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 5092 15892 5120 15932
rect 3568 15864 5120 15892
rect 7576 15892 7604 15932
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 8662 15960 8668 15972
rect 8260 15932 8668 15960
rect 8260 15920 8266 15932
rect 8662 15920 8668 15932
rect 8720 15920 8726 15972
rect 9600 15892 9628 16000
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10520 15904 10548 16068
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 12066 16056 12072 16108
rect 12124 16056 12130 16108
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 12343 16099 12401 16105
rect 12343 16096 12355 16099
rect 12308 16068 12355 16096
rect 12308 16056 12314 16068
rect 12343 16065 12355 16068
rect 12389 16096 12401 16099
rect 13630 16096 13636 16108
rect 12389 16068 13636 16096
rect 12389 16065 12401 16068
rect 12343 16059 12401 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 14643 16099 14701 16105
rect 14643 16096 14655 16099
rect 14332 16068 14655 16096
rect 14332 16056 14338 16068
rect 14643 16065 14655 16068
rect 14689 16096 14701 16099
rect 15010 16096 15016 16108
rect 14689 16068 15016 16096
rect 14689 16065 14701 16068
rect 14643 16059 14701 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 19334 16056 19340 16108
rect 19392 16056 19398 16108
rect 19812 16105 19840 16136
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16096 20683 16099
rect 20714 16096 20720 16108
rect 20671 16068 20720 16096
rect 20671 16065 20683 16068
rect 20625 16059 20683 16065
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 20824 16105 20852 16136
rect 21266 16124 21272 16176
rect 21324 16164 21330 16176
rect 21324 16136 23336 16164
rect 21324 16124 21330 16136
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16065 20867 16099
rect 22891 16099 22949 16105
rect 22891 16096 22903 16099
rect 20809 16059 20867 16065
rect 22066 16068 22903 16096
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 13412 16000 14381 16028
rect 13412 15988 13418 16000
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 17862 15988 17868 16040
rect 17920 15988 17926 16040
rect 13906 15920 13912 15972
rect 13964 15920 13970 15972
rect 20162 15960 20168 15972
rect 19352 15932 20168 15960
rect 7576 15864 9628 15892
rect 3568 15852 3574 15864
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9732 15864 9873 15892
rect 9732 15852 9738 15864
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 9861 15855 9919 15861
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10376 15864 10425 15892
rect 10376 15852 10382 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 13924 15892 13952 15920
rect 10560 15864 13952 15892
rect 10560 15852 10566 15864
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 15746 15892 15752 15904
rect 14332 15864 15752 15892
rect 14332 15852 14338 15864
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 19352 15892 19380 15932
rect 20162 15920 20168 15932
rect 20220 15960 20226 15972
rect 22066 15960 22094 16068
rect 22891 16065 22903 16068
rect 22937 16065 22949 16099
rect 22891 16059 22949 16065
rect 22649 16031 22707 16037
rect 22649 15997 22661 16031
rect 22695 15997 22707 16031
rect 22649 15991 22707 15997
rect 20220 15932 22094 15960
rect 20220 15920 20226 15932
rect 16908 15864 19380 15892
rect 19429 15895 19487 15901
rect 16908 15852 16914 15864
rect 19429 15861 19441 15895
rect 19475 15892 19487 15895
rect 19518 15892 19524 15904
rect 19475 15864 19524 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 19978 15892 19984 15904
rect 19659 15864 19984 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22664 15892 22692 15991
rect 23308 15960 23336 16136
rect 23768 16096 23796 16192
rect 24029 16099 24087 16105
rect 24029 16096 24041 16099
rect 23768 16068 24041 16096
rect 24029 16065 24041 16068
rect 24075 16065 24087 16099
rect 24029 16059 24087 16065
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16096 24179 16099
rect 24394 16096 24400 16108
rect 24167 16068 24400 16096
rect 24167 16065 24179 16068
rect 24121 16059 24179 16065
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 24305 16031 24363 16037
rect 24305 16028 24317 16031
rect 23532 16000 24317 16028
rect 23532 15988 23538 16000
rect 24305 15997 24317 16000
rect 24351 15997 24363 16031
rect 24305 15991 24363 15997
rect 23308 15932 23888 15960
rect 23860 15904 23888 15932
rect 22152 15864 22692 15892
rect 22152 15852 22158 15864
rect 23566 15852 23572 15904
rect 23624 15892 23630 15904
rect 23661 15895 23719 15901
rect 23661 15892 23673 15895
rect 23624 15864 23673 15892
rect 23624 15852 23630 15864
rect 23661 15861 23673 15864
rect 23707 15861 23719 15895
rect 23661 15855 23719 15861
rect 23842 15852 23848 15904
rect 23900 15852 23906 15904
rect 1104 15802 24840 15824
rect 1104 15750 3917 15802
rect 3969 15750 3981 15802
rect 4033 15750 4045 15802
rect 4097 15750 4109 15802
rect 4161 15750 4173 15802
rect 4225 15750 9851 15802
rect 9903 15750 9915 15802
rect 9967 15750 9979 15802
rect 10031 15750 10043 15802
rect 10095 15750 10107 15802
rect 10159 15750 15785 15802
rect 15837 15750 15849 15802
rect 15901 15750 15913 15802
rect 15965 15750 15977 15802
rect 16029 15750 16041 15802
rect 16093 15750 21719 15802
rect 21771 15750 21783 15802
rect 21835 15750 21847 15802
rect 21899 15750 21911 15802
rect 21963 15750 21975 15802
rect 22027 15750 24840 15802
rect 1104 15728 24840 15750
rect 1762 15648 1768 15700
rect 1820 15648 1826 15700
rect 2130 15648 2136 15700
rect 2188 15688 2194 15700
rect 2774 15688 2780 15700
rect 2188 15660 2780 15688
rect 2188 15648 2194 15660
rect 2774 15648 2780 15660
rect 2832 15648 2838 15700
rect 2866 15648 2872 15700
rect 2924 15648 2930 15700
rect 3896 15660 4476 15688
rect 1578 15580 1584 15632
rect 1636 15620 1642 15632
rect 3694 15620 3700 15632
rect 1636 15592 3700 15620
rect 1636 15580 1642 15592
rect 3694 15580 3700 15592
rect 3752 15580 3758 15632
rect 3896 15620 3924 15660
rect 3804 15592 3924 15620
rect 4448 15620 4476 15660
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 4801 15691 4859 15697
rect 4801 15688 4813 15691
rect 4764 15660 4813 15688
rect 4764 15648 4770 15660
rect 4801 15657 4813 15660
rect 4847 15657 4859 15691
rect 7282 15688 7288 15700
rect 4801 15651 4859 15657
rect 5276 15660 7288 15688
rect 5276 15620 5304 15660
rect 4448 15592 5304 15620
rect 1854 15512 1860 15564
rect 1912 15552 1918 15564
rect 3804 15552 3832 15592
rect 1912 15524 3832 15552
rect 1912 15512 1918 15524
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 1946 15484 1952 15496
rect 1719 15456 1952 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15484 2283 15487
rect 2406 15484 2412 15496
rect 2271 15456 2412 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15453 2835 15487
rect 2777 15447 2835 15453
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15484 3479 15487
rect 3694 15484 3700 15496
rect 3467 15456 3700 15484
rect 3467 15453 3479 15456
rect 3421 15447 3479 15453
rect 2792 15416 2820 15447
rect 3694 15444 3700 15456
rect 3752 15444 3758 15496
rect 3804 15493 3832 15524
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 6840 15561 6868 15660
rect 7282 15648 7288 15660
rect 7340 15688 7346 15700
rect 7340 15660 7512 15688
rect 7340 15648 7346 15660
rect 7484 15620 7512 15660
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7616 15660 7849 15688
rect 7616 15648 7622 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 9674 15648 9680 15700
rect 9732 15648 9738 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10652 15660 10793 15688
rect 10652 15648 10658 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 10781 15651 10839 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 16850 15688 16856 15700
rect 12492 15660 16856 15688
rect 12492 15648 12498 15660
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 18325 15691 18383 15697
rect 18325 15657 18337 15691
rect 18371 15688 18383 15691
rect 19334 15688 19340 15700
rect 18371 15660 19340 15688
rect 18371 15657 18383 15660
rect 18325 15651 18383 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 22066 15660 23980 15688
rect 8202 15620 8208 15632
rect 7484 15592 8208 15620
rect 8202 15580 8208 15592
rect 8260 15620 8266 15632
rect 9214 15620 9220 15632
rect 8260 15592 9220 15620
rect 8260 15580 8266 15592
rect 9214 15580 9220 15592
rect 9272 15580 9278 15632
rect 9585 15623 9643 15629
rect 9585 15589 9597 15623
rect 9631 15620 9643 15623
rect 9692 15620 9720 15648
rect 9631 15592 9720 15620
rect 9631 15589 9643 15592
rect 9585 15583 9643 15589
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15521 6883 15555
rect 9674 15552 9680 15564
rect 6825 15515 6883 15521
rect 7438 15524 9680 15552
rect 3789 15487 3847 15493
rect 3789 15453 3801 15487
rect 3835 15453 3847 15487
rect 4062 15484 4068 15496
rect 4023 15456 4068 15484
rect 3789 15447 3847 15453
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 5258 15484 5264 15496
rect 4212 15456 5264 15484
rect 4212 15444 4218 15456
rect 5258 15444 5264 15456
rect 5316 15484 5322 15496
rect 5687 15487 5745 15493
rect 5687 15484 5699 15487
rect 5316 15456 5699 15484
rect 5316 15444 5322 15456
rect 5687 15453 5699 15456
rect 5733 15453 5745 15487
rect 5687 15447 5745 15453
rect 6270 15444 6276 15496
rect 6328 15484 6334 15496
rect 7067 15487 7125 15493
rect 7067 15484 7079 15487
rect 6328 15456 7079 15484
rect 6328 15444 6334 15456
rect 7067 15453 7079 15456
rect 7113 15453 7125 15487
rect 7067 15447 7125 15453
rect 7438 15416 7466 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9950 15512 9956 15564
rect 10008 15561 10014 15564
rect 10008 15555 10036 15561
rect 10024 15521 10036 15555
rect 10008 15515 10036 15521
rect 10008 15512 10014 15515
rect 10318 15512 10324 15564
rect 10376 15552 10382 15564
rect 10376 15524 10732 15552
rect 10376 15512 10382 15524
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 2792 15388 7466 15416
rect 2314 15308 2320 15360
rect 2372 15308 2378 15360
rect 3234 15308 3240 15360
rect 3292 15308 3298 15360
rect 6457 15351 6515 15357
rect 6457 15317 6469 15351
rect 6503 15348 6515 15351
rect 7282 15348 7288 15360
rect 6503 15320 7288 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8956 15348 8984 15447
rect 9122 15444 9128 15496
rect 9180 15444 9186 15496
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 9030 15348 9036 15360
rect 8956 15320 9036 15348
rect 9030 15308 9036 15320
rect 9088 15348 9094 15360
rect 9306 15348 9312 15360
rect 9088 15320 9312 15348
rect 9088 15308 9094 15320
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 9674 15308 9680 15360
rect 9732 15348 9738 15360
rect 10704 15348 10732 15524
rect 12066 15512 12072 15564
rect 12124 15512 12130 15564
rect 18322 15512 18328 15564
rect 18380 15552 18386 15564
rect 19150 15552 19156 15564
rect 18380 15524 19156 15552
rect 18380 15512 18386 15524
rect 19150 15512 19156 15524
rect 19208 15552 19214 15564
rect 19245 15555 19303 15561
rect 19245 15552 19257 15555
rect 19208 15524 19257 15552
rect 19208 15512 19214 15524
rect 19245 15521 19257 15524
rect 19291 15521 19303 15555
rect 19245 15515 19303 15521
rect 20806 15512 20812 15564
rect 20864 15552 20870 15564
rect 22066 15552 22094 15660
rect 20864 15524 22094 15552
rect 20864 15512 20870 15524
rect 22370 15512 22376 15564
rect 22428 15512 22434 15564
rect 10873 15487 10931 15493
rect 10873 15453 10885 15487
rect 10919 15453 10931 15487
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 10873 15447 10931 15453
rect 10888 15416 10916 15447
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11238 15416 11244 15428
rect 10888 15388 11244 15416
rect 11238 15376 11244 15388
rect 11296 15416 11302 15428
rect 12084 15416 12112 15512
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 17218 15484 17224 15496
rect 15068 15456 17224 15484
rect 15068 15444 15074 15456
rect 17218 15444 17224 15456
rect 17276 15484 17282 15496
rect 17678 15484 17684 15496
rect 17276 15456 17684 15484
rect 17276 15444 17282 15456
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18196 15456 18521 15484
rect 18196 15444 18202 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 19503 15457 19561 15463
rect 19503 15454 19515 15457
rect 18509 15447 18567 15453
rect 11296 15388 12112 15416
rect 11296 15376 11302 15388
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 14458 15416 14464 15428
rect 13320 15388 14464 15416
rect 13320 15376 13326 15388
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 17126 15376 17132 15428
rect 17184 15416 17190 15428
rect 17770 15416 17776 15428
rect 17184 15388 17776 15416
rect 17184 15376 17190 15388
rect 17770 15376 17776 15388
rect 17828 15376 17834 15428
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 19444 15426 19515 15454
rect 19444 15416 19472 15426
rect 19503 15423 19515 15426
rect 19549 15423 19561 15457
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 21726 15484 21732 15496
rect 19668 15456 21732 15484
rect 19668 15444 19674 15456
rect 21726 15444 21732 15456
rect 21784 15444 21790 15496
rect 22278 15444 22284 15496
rect 22336 15480 22342 15496
rect 23952 15493 23980 15660
rect 24118 15648 24124 15700
rect 24176 15648 24182 15700
rect 23937 15487 23995 15493
rect 22336 15452 22416 15480
rect 22336 15444 22342 15452
rect 19503 15417 19561 15423
rect 19392 15388 19472 15416
rect 22388 15416 22416 15452
rect 23937 15453 23949 15487
rect 23983 15453 23995 15487
rect 23937 15447 23995 15453
rect 22618 15419 22676 15425
rect 22618 15416 22630 15419
rect 22388 15388 22630 15416
rect 19392 15376 19398 15388
rect 22618 15385 22630 15388
rect 22664 15385 22676 15419
rect 22618 15379 22676 15385
rect 9732 15320 10732 15348
rect 9732 15308 9738 15320
rect 11882 15308 11888 15360
rect 11940 15308 11946 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 14274 15348 14280 15360
rect 12032 15320 14280 15348
rect 12032 15308 12038 15320
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17862 15348 17868 15360
rect 17276 15320 17868 15348
rect 17276 15308 17282 15320
rect 17862 15308 17868 15320
rect 17920 15348 17926 15360
rect 18138 15348 18144 15360
rect 17920 15320 18144 15348
rect 17920 15308 17926 15320
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 19852 15320 20269 15348
rect 19852 15308 19858 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 20438 15308 20444 15360
rect 20496 15348 20502 15360
rect 20990 15348 20996 15360
rect 20496 15320 20996 15348
rect 20496 15308 20502 15320
rect 20990 15308 20996 15320
rect 21048 15308 21054 15360
rect 22094 15308 22100 15360
rect 22152 15308 22158 15360
rect 23750 15308 23756 15360
rect 23808 15308 23814 15360
rect 1104 15258 25000 15280
rect 1104 15206 6884 15258
rect 6936 15206 6948 15258
rect 7000 15206 7012 15258
rect 7064 15206 7076 15258
rect 7128 15206 7140 15258
rect 7192 15206 12818 15258
rect 12870 15206 12882 15258
rect 12934 15206 12946 15258
rect 12998 15206 13010 15258
rect 13062 15206 13074 15258
rect 13126 15206 18752 15258
rect 18804 15206 18816 15258
rect 18868 15206 18880 15258
rect 18932 15206 18944 15258
rect 18996 15206 19008 15258
rect 19060 15206 24686 15258
rect 24738 15206 24750 15258
rect 24802 15206 24814 15258
rect 24866 15206 24878 15258
rect 24930 15206 24942 15258
rect 24994 15206 25000 15258
rect 1104 15184 25000 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 1581 15147 1639 15153
rect 1360 15116 1532 15144
rect 1360 15104 1366 15116
rect 1504 15076 1532 15116
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 2222 15144 2228 15156
rect 1627 15116 2228 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 2222 15104 2228 15116
rect 2280 15104 2286 15156
rect 2516 15116 2866 15144
rect 1504 15048 1900 15076
rect 1762 14968 1768 15020
rect 1820 14968 1826 15020
rect 1872 15017 1900 15048
rect 2131 15021 2189 15027
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 14977 1915 15011
rect 2131 14987 2143 15021
rect 2177 15008 2189 15021
rect 2516 15008 2544 15116
rect 2177 14987 2544 15008
rect 2131 14981 2544 14987
rect 2146 14980 2544 14981
rect 2608 15048 2774 15076
rect 1857 14971 1915 14977
rect 1872 14804 1900 14971
rect 2314 14804 2320 14816
rect 1872 14776 2320 14804
rect 2314 14764 2320 14776
rect 2372 14804 2378 14816
rect 2608 14804 2636 15048
rect 2746 14940 2774 15048
rect 2838 15008 2866 15116
rect 3050 15104 3056 15156
rect 3108 15144 3114 15156
rect 3421 15147 3479 15153
rect 3421 15144 3433 15147
rect 3108 15116 3433 15144
rect 3108 15104 3114 15116
rect 3421 15113 3433 15116
rect 3467 15113 3479 15147
rect 3421 15107 3479 15113
rect 3970 15104 3976 15156
rect 4028 15104 4034 15156
rect 4154 15104 4160 15156
rect 4212 15104 4218 15156
rect 6454 15144 6460 15156
rect 4356 15116 6460 15144
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 3329 15079 3387 15085
rect 3329 15076 3341 15079
rect 3292 15048 3341 15076
rect 3292 15036 3298 15048
rect 3329 15045 3341 15048
rect 3375 15045 3387 15079
rect 4172 15076 4200 15104
rect 4356 15088 4384 15116
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 7374 15144 7380 15156
rect 6564 15116 7380 15144
rect 3329 15039 3387 15045
rect 3712 15048 4200 15076
rect 3712 15008 3740 15048
rect 4338 15036 4344 15088
rect 4396 15036 4402 15088
rect 5258 15076 5264 15088
rect 4724 15048 5264 15076
rect 2838 14980 3740 15008
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 3844 14980 3893 15008
rect 3844 14968 3850 14980
rect 3881 14977 3893 14980
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 4615 15011 4673 15017
rect 4615 15008 4627 15011
rect 4304 14980 4627 15008
rect 4304 14968 4310 14980
rect 4615 14977 4627 14980
rect 4661 15008 4673 15011
rect 4724 15008 4752 15048
rect 5258 15036 5264 15048
rect 5316 15036 5322 15088
rect 4661 14980 4752 15008
rect 4661 14977 4673 14980
rect 4615 14971 4673 14977
rect 4982 14968 4988 15020
rect 5040 15008 5046 15020
rect 6564 15017 6592 15116
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 9398 15104 9404 15156
rect 9456 15104 9462 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 10192 15116 10241 15144
rect 10192 15104 10198 15116
rect 10229 15113 10241 15116
rect 10275 15113 10287 15147
rect 10229 15107 10287 15113
rect 11606 15104 11612 15156
rect 11664 15144 11670 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 11664 15116 11713 15144
rect 11664 15104 11670 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 11701 15107 11759 15113
rect 11790 15104 11796 15156
rect 11848 15104 11854 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12676 15116 12817 15144
rect 12676 15104 12682 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 16942 15144 16948 15156
rect 13504 15116 16948 15144
rect 13504 15104 13510 15116
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 19705 15147 19763 15153
rect 17050 15116 17908 15144
rect 7466 15017 7472 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5040 14980 6561 15008
rect 5040 14968 5046 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7423 15011 7472 15017
rect 7423 14977 7435 15011
rect 7469 14977 7472 15011
rect 7423 14971 7472 14977
rect 7466 14968 7472 14971
rect 7524 14968 7530 15020
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 9416 15008 9444 15104
rect 11146 15036 11152 15088
rect 11204 15076 11210 15088
rect 11808 15076 11836 15104
rect 17050 15076 17078 15116
rect 11204 15048 13584 15076
rect 11204 15036 11210 15048
rect 9475 15011 9533 15017
rect 9475 15008 9487 15011
rect 9416 14980 9487 15008
rect 9475 14977 9487 14980
rect 9521 14977 9533 15011
rect 9475 14971 9533 14977
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 11974 15008 11980 15020
rect 11848 14980 11980 15008
rect 11848 14968 11854 14980
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12066 14968 12072 15020
rect 12124 14968 12130 15020
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 13446 15008 13452 15020
rect 12492 14980 13452 15008
rect 12492 14968 12498 14980
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 13556 15008 13584 15048
rect 14292 15048 17078 15076
rect 14151 15021 14209 15027
rect 14151 15008 14163 15021
rect 13556 14987 14163 15008
rect 14197 15018 14209 15021
rect 14197 15008 14210 15018
rect 14292 15008 14320 15048
rect 17880 15020 17908 15116
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20806 15144 20812 15156
rect 19751 15116 20812 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 22094 15104 22100 15156
rect 22152 15104 22158 15156
rect 22738 15104 22744 15156
rect 22796 15144 22802 15156
rect 23566 15144 23572 15156
rect 22796 15116 23572 15144
rect 22796 15104 22802 15116
rect 23566 15104 23572 15116
rect 23624 15104 23630 15156
rect 18138 15036 18144 15088
rect 18196 15076 18202 15088
rect 19610 15076 19616 15088
rect 18196 15048 19616 15076
rect 18196 15036 18202 15048
rect 19610 15036 19616 15048
rect 19668 15076 19674 15088
rect 19668 15048 20300 15076
rect 19668 15036 19674 15048
rect 14197 14987 14320 15008
rect 13556 14980 14320 14987
rect 15286 14968 15292 15020
rect 15344 14968 15350 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17218 15008 17224 15020
rect 17175 14980 17224 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 17402 15017 17408 15020
rect 17396 15008 17408 15017
rect 17363 14980 17408 15008
rect 17396 14971 17408 14980
rect 17402 14968 17408 14971
rect 17460 14968 17466 15020
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 19334 15008 19340 15020
rect 17920 14980 19340 15008
rect 17920 14968 17926 14980
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 4341 14943 4399 14949
rect 4341 14940 4353 14943
rect 2746 14912 4353 14940
rect 4341 14909 4353 14912
rect 4387 14909 4399 14943
rect 4341 14903 4399 14909
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14940 6423 14943
rect 6638 14940 6644 14952
rect 6411 14912 6644 14940
rect 6411 14909 6423 14912
rect 6365 14903 6423 14909
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 2832 14844 3280 14872
rect 2832 14832 2838 14844
rect 3252 14816 3280 14844
rect 2372 14776 2636 14804
rect 2372 14764 2378 14776
rect 2866 14764 2872 14816
rect 2924 14764 2930 14816
rect 3234 14764 3240 14816
rect 3292 14764 3298 14816
rect 4356 14804 4384 14903
rect 6380 14872 6408 14903
rect 6638 14900 6644 14912
rect 6696 14900 6702 14952
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6748 14912 7297 14940
rect 5000 14844 6408 14872
rect 4706 14804 4712 14816
rect 4356 14776 4712 14804
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 4798 14764 4804 14816
rect 4856 14804 4862 14816
rect 5000 14804 5028 14844
rect 6454 14832 6460 14884
rect 6512 14872 6518 14884
rect 6748 14872 6776 14912
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 7558 14900 7564 14952
rect 7616 14900 7622 14952
rect 11882 14900 11888 14952
rect 11940 14900 11946 14952
rect 12802 14900 12808 14952
rect 12860 14940 12866 14952
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 12860 14912 13921 14940
rect 12860 14900 12866 14912
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 15304 14940 15332 14968
rect 13909 14903 13967 14909
rect 14568 14912 15332 14940
rect 19444 14940 19472 14971
rect 19518 14968 19524 15020
rect 19576 14968 19582 15020
rect 19794 15008 19800 15020
rect 19628 14980 19800 15008
rect 19628 14940 19656 14980
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20272 15017 20300 15048
rect 20346 15036 20352 15088
rect 20404 15076 20410 15088
rect 20524 15079 20582 15085
rect 20524 15076 20536 15079
rect 20404 15048 20536 15076
rect 20404 15036 20410 15048
rect 20524 15045 20536 15048
rect 20570 15045 20582 15079
rect 22112 15076 22140 15104
rect 22112 15048 23428 15076
rect 20524 15039 20582 15045
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 22063 15011 22121 15017
rect 22063 15008 22075 15011
rect 20257 14971 20315 14977
rect 20364 14980 22075 15008
rect 19444 14912 19656 14940
rect 19705 14943 19763 14949
rect 6512 14844 6776 14872
rect 7009 14875 7067 14881
rect 6512 14832 6518 14844
rect 7009 14841 7021 14875
rect 7055 14841 7067 14875
rect 7009 14835 7067 14841
rect 4856 14776 5028 14804
rect 4856 14764 4862 14776
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 5442 14764 5448 14816
rect 5500 14804 5506 14816
rect 5902 14804 5908 14816
rect 5500 14776 5908 14804
rect 5500 14764 5506 14776
rect 5902 14764 5908 14776
rect 5960 14804 5966 14816
rect 6822 14804 6828 14816
rect 5960 14776 6828 14804
rect 5960 14764 5966 14776
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 7024 14804 7052 14835
rect 7282 14804 7288 14816
rect 7024 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 8202 14764 8208 14816
rect 8260 14764 8266 14816
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13998 14804 14004 14816
rect 13035 14776 14004 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13998 14764 14004 14776
rect 14056 14804 14062 14816
rect 14568 14804 14596 14912
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19751 14912 19901 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 20364 14940 20392 14980
rect 22063 14977 22075 14980
rect 22109 14977 22121 15011
rect 22063 14971 22121 14977
rect 22186 14968 22192 15020
rect 22244 15008 22250 15020
rect 22462 15008 22468 15020
rect 22244 14980 22468 15008
rect 22244 14968 22250 14980
rect 22462 14968 22468 14980
rect 22520 15008 22526 15020
rect 23400 15017 23428 15048
rect 23385 15011 23443 15017
rect 22520 14980 22876 15008
rect 22520 14968 22526 14980
rect 19889 14903 19947 14909
rect 19996 14912 20392 14940
rect 14642 14832 14648 14884
rect 14700 14872 14706 14884
rect 14700 14844 15056 14872
rect 14700 14832 14706 14844
rect 14056 14776 14596 14804
rect 14056 14764 14062 14776
rect 14918 14764 14924 14816
rect 14976 14764 14982 14816
rect 15028 14804 15056 14844
rect 16206 14832 16212 14884
rect 16264 14872 16270 14884
rect 16666 14872 16672 14884
rect 16264 14844 16672 14872
rect 16264 14832 16270 14844
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 19996 14872 20024 14912
rect 21726 14900 21732 14952
rect 21784 14940 21790 14952
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21784 14912 21833 14940
rect 21784 14900 21790 14912
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 21821 14903 21879 14909
rect 18064 14844 20024 14872
rect 18064 14804 18092 14844
rect 15028 14776 18092 14804
rect 18506 14764 18512 14816
rect 18564 14764 18570 14816
rect 18690 14764 18696 14816
rect 18748 14804 18754 14816
rect 19886 14804 19892 14816
rect 18748 14776 19892 14804
rect 18748 14764 18754 14776
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 21634 14764 21640 14816
rect 21692 14764 21698 14816
rect 21836 14804 21864 14903
rect 22848 14881 22876 14980
rect 23385 14977 23397 15011
rect 23431 14977 23443 15011
rect 23584 15008 23612 15104
rect 23753 15079 23811 15085
rect 23753 15045 23765 15079
rect 23799 15076 23811 15079
rect 24302 15076 24308 15088
rect 23799 15048 24308 15076
rect 23799 15045 23811 15048
rect 23753 15039 23811 15045
rect 24302 15036 24308 15048
rect 24360 15036 24366 15088
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23584 14980 24225 15008
rect 23385 14971 23443 14977
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 23014 14900 23020 14952
rect 23072 14940 23078 14952
rect 24489 14943 24547 14949
rect 24489 14940 24501 14943
rect 23072 14912 24501 14940
rect 23072 14900 23078 14912
rect 24489 14909 24501 14912
rect 24535 14909 24547 14943
rect 24489 14903 24547 14909
rect 22833 14875 22891 14881
rect 22833 14841 22845 14875
rect 22879 14841 22891 14875
rect 22833 14835 22891 14841
rect 23477 14875 23535 14881
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 24305 14875 24363 14881
rect 24305 14872 24317 14875
rect 23523 14844 24317 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 24305 14841 24317 14844
rect 24351 14841 24363 14875
rect 24305 14835 24363 14841
rect 22278 14804 22284 14816
rect 21836 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 24026 14764 24032 14816
rect 24084 14764 24090 14816
rect 24397 14807 24455 14813
rect 24397 14773 24409 14807
rect 24443 14804 24455 14807
rect 24443 14776 24900 14804
rect 24443 14773 24455 14776
rect 24397 14767 24455 14773
rect 1104 14714 24840 14736
rect 1104 14662 3917 14714
rect 3969 14662 3981 14714
rect 4033 14662 4045 14714
rect 4097 14662 4109 14714
rect 4161 14662 4173 14714
rect 4225 14662 9851 14714
rect 9903 14662 9915 14714
rect 9967 14662 9979 14714
rect 10031 14662 10043 14714
rect 10095 14662 10107 14714
rect 10159 14662 15785 14714
rect 15837 14662 15849 14714
rect 15901 14662 15913 14714
rect 15965 14662 15977 14714
rect 16029 14662 16041 14714
rect 16093 14662 21719 14714
rect 21771 14662 21783 14714
rect 21835 14662 21847 14714
rect 21899 14662 21911 14714
rect 21963 14662 21975 14714
rect 22027 14662 24840 14714
rect 1104 14640 24840 14662
rect 2866 14600 2872 14612
rect 2424 14572 2872 14600
rect 2424 14541 2452 14572
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 3786 14560 3792 14612
rect 3844 14600 3850 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 3844 14572 4077 14600
rect 3844 14560 3850 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4065 14563 4123 14569
rect 4448 14572 7512 14600
rect 2409 14535 2467 14541
rect 2409 14501 2421 14535
rect 2455 14501 2467 14535
rect 4338 14532 4344 14544
rect 2409 14495 2467 14501
rect 3896 14504 4344 14532
rect 2866 14473 2872 14476
rect 2823 14467 2872 14473
rect 2823 14433 2835 14467
rect 2869 14433 2872 14467
rect 2823 14427 2872 14433
rect 2866 14424 2872 14427
rect 2924 14464 2930 14476
rect 3896 14464 3924 14504
rect 4338 14492 4344 14504
rect 4396 14492 4402 14544
rect 4448 14464 4476 14572
rect 5350 14492 5356 14544
rect 5408 14532 5414 14544
rect 5537 14535 5595 14541
rect 5537 14532 5549 14535
rect 5408 14504 5549 14532
rect 5408 14492 5414 14504
rect 5537 14501 5549 14504
rect 5583 14501 5595 14535
rect 7484 14532 7512 14572
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7616 14572 7849 14600
rect 7616 14560 7622 14572
rect 7837 14569 7849 14572
rect 7883 14569 7895 14603
rect 7837 14563 7895 14569
rect 8202 14560 8208 14612
rect 8260 14560 8266 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 11146 14600 11152 14612
rect 8904 14572 11152 14600
rect 8904 14560 8910 14572
rect 11146 14560 11152 14572
rect 11204 14560 11210 14612
rect 11256 14572 12020 14600
rect 8220 14532 8248 14560
rect 7484 14504 8248 14532
rect 5537 14495 5595 14501
rect 10134 14492 10140 14544
rect 10192 14532 10198 14544
rect 10502 14532 10508 14544
rect 10192 14504 10508 14532
rect 10192 14492 10198 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 11256 14532 11284 14572
rect 11164 14504 11284 14532
rect 2924 14436 3924 14464
rect 3988 14436 4476 14464
rect 4617 14467 4675 14473
rect 2924 14424 2930 14436
rect 934 14356 940 14408
rect 992 14396 998 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 992 14368 1777 14396
rect 992 14356 998 14368
rect 1765 14365 1777 14368
rect 1811 14396 1823 14399
rect 1854 14396 1860 14408
rect 1811 14368 1860 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 2682 14356 2688 14408
rect 2740 14356 2746 14408
rect 2958 14356 2964 14408
rect 3016 14356 3022 14408
rect 3988 14405 4016 14436
rect 4617 14433 4629 14467
rect 4663 14464 4675 14467
rect 5951 14467 6009 14473
rect 5951 14464 5963 14467
rect 4663 14436 5963 14464
rect 4663 14433 4675 14436
rect 4617 14427 4675 14433
rect 5951 14433 5963 14436
rect 5997 14464 6009 14467
rect 6454 14464 6460 14476
rect 5997 14436 6460 14464
rect 5997 14433 6009 14436
rect 5951 14427 6009 14433
rect 6454 14424 6460 14436
rect 6512 14424 6518 14476
rect 6822 14424 6828 14476
rect 6880 14424 6886 14476
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 10410 14464 10416 14476
rect 8168 14436 10416 14464
rect 8168 14424 8174 14436
rect 10410 14424 10416 14436
rect 10468 14424 10474 14476
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4246 14356 4252 14408
rect 4304 14356 4310 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4856 14368 4905 14396
rect 4856 14356 4862 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 4982 14356 4988 14408
rect 5040 14396 5046 14408
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 5040 14368 5089 14396
rect 5040 14356 5046 14368
rect 5077 14365 5089 14368
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 5810 14356 5816 14408
rect 5868 14356 5874 14408
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 7083 14369 7141 14375
rect 7083 14366 7095 14369
rect 6748 14328 6776 14356
rect 7082 14335 7095 14366
rect 7129 14335 7141 14369
rect 7650 14356 7656 14408
rect 7708 14396 7714 14408
rect 8018 14396 8024 14408
rect 7708 14368 8024 14396
rect 7708 14356 7714 14368
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 9398 14356 9404 14408
rect 9456 14396 9462 14408
rect 10042 14396 10048 14408
rect 9456 14368 10048 14396
rect 9456 14356 9462 14368
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 7082 14329 7141 14335
rect 7082 14328 7110 14329
rect 3436 14300 3832 14328
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 3436 14260 3464 14300
rect 2556 14232 3464 14260
rect 2556 14220 2562 14232
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 3804 14269 3832 14300
rect 6564 14300 7110 14328
rect 3605 14263 3663 14269
rect 3605 14260 3617 14263
rect 3568 14232 3617 14260
rect 3568 14220 3574 14232
rect 3605 14229 3617 14232
rect 3651 14229 3663 14263
rect 3605 14223 3663 14229
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 6564 14260 6592 14300
rect 7374 14288 7380 14340
rect 7432 14328 7438 14340
rect 11164 14328 11192 14504
rect 11238 14424 11244 14476
rect 11296 14424 11302 14476
rect 11422 14396 11428 14408
rect 7432 14300 11192 14328
rect 11348 14368 11428 14396
rect 7432 14288 7438 14300
rect 4856 14232 6592 14260
rect 4856 14220 4862 14232
rect 6730 14220 6736 14272
rect 6788 14220 6794 14272
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 11054 14260 11060 14272
rect 6972 14232 11060 14260
rect 6972 14220 6978 14232
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 11348 14260 11376 14368
rect 11422 14356 11428 14368
rect 11480 14405 11486 14408
rect 11480 14399 11541 14405
rect 11480 14365 11495 14399
rect 11529 14365 11541 14399
rect 11480 14359 11541 14365
rect 11480 14356 11486 14359
rect 11992 14328 12020 14572
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 12124 14572 12265 14600
rect 12124 14560 12130 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 13630 14560 13636 14612
rect 13688 14600 13694 14612
rect 14642 14600 14648 14612
rect 13688 14572 14648 14600
rect 13688 14560 13694 14572
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 14918 14560 14924 14612
rect 14976 14560 14982 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 18049 14603 18107 14609
rect 18049 14600 18061 14603
rect 15344 14572 18061 14600
rect 15344 14560 15350 14572
rect 18049 14569 18061 14572
rect 18095 14569 18107 14603
rect 18049 14563 18107 14569
rect 18506 14560 18512 14612
rect 18564 14560 18570 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 23290 14600 23296 14612
rect 20864 14572 23296 14600
rect 20864 14560 20870 14572
rect 23290 14560 23296 14572
rect 23348 14560 23354 14612
rect 24872 14600 24900 14776
rect 23492 14572 24900 14600
rect 13446 14492 13452 14544
rect 13504 14532 13510 14544
rect 13504 14504 14504 14532
rect 13504 14492 13510 14504
rect 14476 14473 14504 14504
rect 14936 14473 14964 14560
rect 16206 14532 16212 14544
rect 15948 14504 16212 14532
rect 14461 14467 14519 14473
rect 14461 14433 14473 14467
rect 14507 14433 14519 14467
rect 14461 14427 14519 14433
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14433 14979 14467
rect 14921 14427 14979 14433
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 15068 14436 15209 14464
rect 15068 14424 15074 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 15335 14467 15393 14473
rect 15335 14433 15347 14467
rect 15381 14464 15393 14467
rect 15948 14464 15976 14504
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 15381 14436 15976 14464
rect 15381 14433 15393 14436
rect 15335 14427 15393 14433
rect 16022 14424 16028 14476
rect 16080 14424 16086 14476
rect 16482 14430 16488 14476
rect 16408 14424 16488 14430
rect 16540 14424 16546 14476
rect 16850 14424 16856 14476
rect 16908 14424 16914 14476
rect 17126 14424 17132 14476
rect 17184 14424 17190 14476
rect 17218 14424 17224 14476
rect 17276 14473 17282 14476
rect 17276 14467 17304 14473
rect 17292 14433 17304 14467
rect 17276 14427 17304 14433
rect 17276 14424 17282 14427
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12618 14396 12624 14408
rect 12124 14368 12624 14396
rect 12124 14356 12130 14368
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 12894 14396 12900 14408
rect 12855 14368 12900 14396
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 14274 14356 14280 14408
rect 14332 14356 14338 14408
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 16040 14396 16068 14424
rect 16408 14405 16528 14424
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 16040 14368 16221 14396
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16393 14402 16528 14405
rect 16393 14399 16451 14402
rect 16393 14365 16405 14399
rect 16439 14365 16451 14399
rect 16393 14359 16451 14365
rect 17402 14356 17408 14408
rect 17460 14356 17466 14408
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 17972 14368 18337 14396
rect 16117 14331 16175 14337
rect 11992 14300 13768 14328
rect 11204 14232 11376 14260
rect 11204 14220 11210 14232
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13228 14232 13645 14260
rect 13228 14220 13234 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13740 14260 13768 14300
rect 16117 14297 16129 14331
rect 16163 14297 16175 14331
rect 16117 14291 16175 14297
rect 16132 14260 16160 14291
rect 13740 14232 16160 14260
rect 13633 14223 13691 14229
rect 17494 14220 17500 14272
rect 17552 14260 17558 14272
rect 17972 14260 18000 14368
rect 18325 14365 18337 14368
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18524 14396 18552 14560
rect 21545 14535 21603 14541
rect 21545 14501 21557 14535
rect 21591 14532 21603 14535
rect 21913 14535 21971 14541
rect 21913 14532 21925 14535
rect 21591 14504 21925 14532
rect 21591 14501 21603 14504
rect 21545 14495 21603 14501
rect 21913 14501 21925 14504
rect 21959 14501 21971 14535
rect 21913 14495 21971 14501
rect 21634 14424 21640 14476
rect 21692 14424 21698 14476
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 22557 14467 22615 14473
rect 22557 14464 22569 14467
rect 22143 14436 22569 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 22557 14433 22569 14436
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18524 14368 18889 14396
rect 18417 14359 18475 14365
rect 18877 14365 18889 14368
rect 18923 14365 18935 14399
rect 18877 14359 18935 14365
rect 18432 14328 18460 14359
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20404 14368 21097 14396
rect 20404 14356 20410 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 21468 14328 21496 14359
rect 18156 14300 18460 14328
rect 20916 14300 21496 14328
rect 21652 14328 21680 14424
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22186 14396 22192 14408
rect 21867 14368 22192 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22186 14356 22192 14368
rect 22244 14356 22250 14408
rect 22365 14399 22423 14405
rect 22365 14396 22377 14399
rect 22296 14368 22377 14396
rect 22296 14328 22324 14368
rect 22365 14365 22377 14368
rect 22411 14365 22423 14399
rect 22365 14359 22423 14365
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 22649 14399 22707 14405
rect 22649 14396 22661 14399
rect 22572 14368 22661 14396
rect 21652 14300 22324 14328
rect 18156 14269 18184 14300
rect 17552 14232 18000 14260
rect 18141 14263 18199 14269
rect 17552 14220 17558 14232
rect 18141 14229 18153 14263
rect 18187 14229 18199 14263
rect 18141 14223 18199 14229
rect 18506 14220 18512 14272
rect 18564 14220 18570 14272
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 19150 14260 19156 14272
rect 18739 14232 19156 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 20916 14269 20944 14300
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14229 20959 14263
rect 20901 14223 20959 14229
rect 22094 14220 22100 14272
rect 22152 14220 22158 14272
rect 22189 14263 22247 14269
rect 22189 14229 22201 14263
rect 22235 14260 22247 14263
rect 22572 14260 22600 14368
rect 22649 14365 22661 14368
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 23293 14399 23351 14405
rect 23293 14365 23305 14399
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 23385 14399 23443 14405
rect 23385 14365 23397 14399
rect 23431 14396 23443 14399
rect 23492 14396 23520 14572
rect 23569 14535 23627 14541
rect 23569 14501 23581 14535
rect 23615 14532 23627 14535
rect 25130 14532 25136 14544
rect 23615 14504 25136 14532
rect 23615 14501 23627 14504
rect 23569 14495 23627 14501
rect 25130 14492 25136 14504
rect 25188 14492 25194 14544
rect 23750 14424 23756 14476
rect 23808 14424 23814 14476
rect 23431 14368 23520 14396
rect 23431 14365 23443 14368
rect 23385 14359 23443 14365
rect 23308 14328 23336 14359
rect 23768 14328 23796 14424
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 24210 14396 24216 14408
rect 23891 14368 24216 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 24210 14356 24216 14368
rect 24268 14356 24274 14408
rect 23308 14300 23796 14328
rect 22235 14232 22600 14260
rect 22235 14229 22247 14232
rect 22189 14223 22247 14229
rect 23106 14220 23112 14272
rect 23164 14220 23170 14272
rect 24121 14263 24179 14269
rect 24121 14229 24133 14263
rect 24167 14260 24179 14263
rect 25314 14260 25320 14272
rect 24167 14232 25320 14260
rect 24167 14229 24179 14232
rect 24121 14223 24179 14229
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 1104 14170 25000 14192
rect 1104 14118 6884 14170
rect 6936 14118 6948 14170
rect 7000 14118 7012 14170
rect 7064 14118 7076 14170
rect 7128 14118 7140 14170
rect 7192 14118 12818 14170
rect 12870 14118 12882 14170
rect 12934 14118 12946 14170
rect 12998 14118 13010 14170
rect 13062 14118 13074 14170
rect 13126 14118 18752 14170
rect 18804 14118 18816 14170
rect 18868 14118 18880 14170
rect 18932 14118 18944 14170
rect 18996 14118 19008 14170
rect 19060 14118 24686 14170
rect 24738 14118 24750 14170
rect 24802 14118 24814 14170
rect 24866 14118 24878 14170
rect 24930 14118 24942 14170
rect 24994 14118 25000 14170
rect 1104 14096 25000 14118
rect 25314 14084 25320 14136
rect 25372 14124 25378 14136
rect 25866 14124 25872 14136
rect 25372 14096 25872 14124
rect 25372 14084 25378 14096
rect 25866 14084 25872 14096
rect 25924 14084 25930 14136
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 3016 14028 3249 14056
rect 3016 14016 3022 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 3326 14016 3332 14068
rect 3384 14056 3390 14068
rect 3789 14059 3847 14065
rect 3789 14056 3801 14059
rect 3384 14028 3801 14056
rect 3384 14016 3390 14028
rect 3789 14025 3801 14028
rect 3835 14025 3847 14059
rect 4798 14056 4804 14068
rect 3789 14019 3847 14025
rect 3896 14028 4804 14056
rect 1489 13991 1547 13997
rect 1489 13957 1501 13991
rect 1535 13988 1547 13991
rect 1578 13988 1584 14000
rect 1535 13960 1584 13988
rect 1535 13957 1547 13960
rect 1489 13951 1547 13957
rect 1578 13948 1584 13960
rect 1636 13948 1642 14000
rect 3896 13988 3924 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 6086 14056 6092 14068
rect 5951 14028 6092 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 7650 14056 7656 14068
rect 6932 14028 7656 14056
rect 6748 13988 6776 14016
rect 3620 13960 3924 13988
rect 4632 13960 6776 13988
rect 2130 13880 2136 13932
rect 2188 13880 2194 13932
rect 2499 13923 2557 13929
rect 2499 13889 2511 13923
rect 2545 13920 2557 13923
rect 3620 13920 3648 13960
rect 2545 13892 3648 13920
rect 3697 13923 3755 13929
rect 2545 13889 2557 13892
rect 2499 13883 2557 13889
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 1486 13812 1492 13864
rect 1544 13852 1550 13864
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 1544 13824 1777 13852
rect 1544 13812 1550 13824
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 2240 13784 2268 13815
rect 3712 13784 3740 13883
rect 4338 13880 4344 13932
rect 4396 13880 4402 13932
rect 4632 13929 4660 13960
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 4706 13880 4712 13932
rect 4764 13920 4770 13932
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4764 13892 4905 13920
rect 4764 13880 4770 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5167 13923 5225 13929
rect 5167 13920 5179 13923
rect 5132 13892 5179 13920
rect 5132 13880 5138 13892
rect 5167 13889 5179 13892
rect 5213 13889 5225 13923
rect 5167 13883 5225 13889
rect 5902 13880 5908 13932
rect 5960 13880 5966 13932
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 6932 13920 6960 14028
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 7834 14016 7840 14068
rect 7892 14056 7898 14068
rect 9766 14056 9772 14068
rect 7892 14028 9772 14056
rect 7892 14016 7898 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10042 14016 10048 14068
rect 10100 14016 10106 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10376 14028 10609 14056
rect 10376 14016 10382 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 10597 14019 10655 14025
rect 12406 14028 14289 14056
rect 7006 13948 7012 14000
rect 7064 13988 7070 14000
rect 7064 13960 7218 13988
rect 7064 13948 7070 13960
rect 7099 13923 7157 13929
rect 7099 13920 7111 13923
rect 6512 13892 7111 13920
rect 6512 13880 6518 13892
rect 7099 13889 7111 13892
rect 7145 13889 7157 13923
rect 7190 13920 7218 13960
rect 8018 13948 8024 14000
rect 8076 13988 8082 14000
rect 9674 13988 9680 14000
rect 8076 13960 9680 13988
rect 8076 13948 8082 13960
rect 9674 13948 9680 13960
rect 9732 13948 9738 14000
rect 9858 13959 9864 14000
rect 9843 13953 9864 13959
rect 8205 13923 8263 13929
rect 8205 13920 8217 13923
rect 7190 13892 8217 13920
rect 7099 13883 7157 13889
rect 8205 13889 8217 13892
rect 8251 13889 8263 13923
rect 8205 13883 8263 13889
rect 8479 13923 8537 13929
rect 8479 13889 8491 13923
rect 8525 13920 8537 13923
rect 9398 13920 9404 13932
rect 8525 13892 9404 13920
rect 8525 13889 8537 13892
rect 8479 13883 8537 13889
rect 5920 13852 5948 13880
rect 6822 13852 6828 13864
rect 5920 13824 6828 13852
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 8018 13784 8024 13796
rect 2240 13756 2360 13784
rect 3712 13756 5028 13784
rect 2332 13728 2360 13756
rect 1946 13676 1952 13728
rect 2004 13676 2010 13728
rect 2314 13676 2320 13728
rect 2372 13676 2378 13728
rect 3326 13676 3332 13728
rect 3384 13716 3390 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 3384 13688 4169 13716
rect 3384 13676 3390 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4157 13679 4215 13685
rect 4430 13676 4436 13728
rect 4488 13676 4494 13728
rect 5000 13716 5028 13756
rect 7760 13756 8024 13784
rect 7760 13716 7788 13756
rect 8018 13744 8024 13756
rect 8076 13744 8082 13796
rect 5000 13688 7788 13716
rect 7834 13676 7840 13728
rect 7892 13676 7898 13728
rect 8220 13716 8248 13883
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13889 9643 13923
rect 9843 13919 9855 13953
rect 9916 13948 9922 14000
rect 10060 13988 10088 14016
rect 12406 13988 12434 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 14277 14019 14335 14025
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 15528 14028 15669 14056
rect 15528 14016 15534 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17460 14028 17693 14056
rect 17460 14016 17466 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 19150 14016 19156 14068
rect 19208 14016 19214 14068
rect 19610 14016 19616 14068
rect 19668 14056 19674 14068
rect 21174 14056 21180 14068
rect 19668 14028 21180 14056
rect 19668 14016 19674 14028
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 23106 14056 23112 14068
rect 22940 14028 23112 14056
rect 10060 13960 12434 13988
rect 14458 13948 14464 14000
rect 14516 13988 14522 14000
rect 16666 13988 16672 14000
rect 14516 13960 16672 13988
rect 14516 13948 14522 13960
rect 16666 13948 16672 13960
rect 16724 13948 16730 14000
rect 9889 13922 9902 13948
rect 12437 13923 12495 13929
rect 9889 13919 9901 13922
rect 9843 13913 9901 13919
rect 9585 13883 9643 13889
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12483 13892 12848 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 9490 13784 9496 13796
rect 9140 13756 9496 13784
rect 9140 13716 9168 13756
rect 9490 13744 9496 13756
rect 9548 13784 9554 13796
rect 9600 13784 9628 13883
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12820 13852 12848 13892
rect 13630 13880 13636 13932
rect 13688 13880 13694 13932
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 14887 13923 14945 13929
rect 14887 13920 14899 13923
rect 14332 13892 14899 13920
rect 14332 13880 14338 13892
rect 14887 13889 14899 13892
rect 14933 13889 14945 13923
rect 16942 13920 16948 13932
rect 16903 13892 16948 13920
rect 14887 13883 14945 13889
rect 16942 13880 16948 13892
rect 17000 13920 17006 13932
rect 17402 13920 17408 13932
rect 17000 13892 17408 13920
rect 17000 13880 17006 13892
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 18064 13920 18092 14016
rect 19168 13988 19196 14016
rect 19168 13960 19656 13988
rect 18291 13923 18349 13929
rect 18291 13920 18303 13923
rect 18064 13892 18303 13920
rect 18291 13889 18303 13892
rect 18337 13889 18349 13923
rect 18291 13883 18349 13889
rect 19058 13880 19064 13932
rect 19116 13920 19122 13932
rect 19628 13929 19656 13960
rect 19978 13948 19984 14000
rect 20036 13988 20042 14000
rect 21634 13988 21640 14000
rect 20036 13960 21640 13988
rect 20036 13948 20042 13960
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 22940 13935 22968 14028
rect 23106 14016 23112 14028
rect 23164 14016 23170 14068
rect 23201 14059 23259 14065
rect 23201 14025 23213 14059
rect 23247 14025 23259 14059
rect 23201 14019 23259 14025
rect 23216 13988 23244 14019
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23348 14028 24164 14056
rect 23348 14016 23354 14028
rect 24136 13997 24164 14028
rect 25774 14016 25780 14068
rect 25832 14016 25838 14068
rect 23845 13991 23903 13997
rect 23845 13988 23857 13991
rect 23216 13960 23857 13988
rect 23845 13957 23857 13960
rect 23891 13957 23903 13991
rect 23845 13951 23903 13957
rect 24121 13991 24179 13997
rect 24121 13957 24133 13991
rect 24167 13957 24179 13991
rect 24121 13951 24179 13957
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 19116 13892 19441 13920
rect 19116 13880 19122 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 21542 13880 21548 13932
rect 21600 13880 21606 13932
rect 22738 13880 22744 13932
rect 22796 13880 22802 13932
rect 22916 13929 22974 13935
rect 22916 13895 22928 13929
rect 22962 13895 22974 13929
rect 22916 13889 22974 13895
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13889 23075 13923
rect 23017 13883 23075 13889
rect 12986 13852 12992 13864
rect 12820 13824 12992 13852
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13078 13812 13084 13864
rect 13136 13812 13142 13864
rect 13170 13812 13176 13864
rect 13228 13852 13234 13864
rect 13538 13861 13544 13864
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 13228 13824 13369 13852
rect 13228 13812 13234 13824
rect 13357 13821 13369 13824
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 13495 13855 13544 13861
rect 13495 13821 13507 13855
rect 13541 13821 13544 13855
rect 13495 13815 13544 13821
rect 13538 13812 13544 13815
rect 13596 13852 13602 13864
rect 13998 13852 14004 13864
rect 13596 13824 14004 13852
rect 13596 13812 13602 13824
rect 13998 13812 14004 13824
rect 14056 13812 14062 13864
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 16669 13855 16727 13861
rect 16669 13821 16681 13855
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 18049 13855 18107 13861
rect 18049 13821 18061 13855
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18984 13824 19748 13852
rect 9548 13756 9674 13784
rect 9548 13744 9554 13756
rect 8220 13688 9168 13716
rect 9214 13676 9220 13728
rect 9272 13676 9278 13728
rect 9646 13716 9674 13756
rect 11882 13716 11888 13728
rect 9646 13688 11888 13716
rect 11882 13676 11888 13688
rect 11940 13716 11946 13728
rect 14658 13716 14686 13815
rect 16684 13784 16712 13815
rect 16684 13756 16804 13784
rect 16776 13728 16804 13756
rect 14918 13716 14924 13728
rect 11940 13688 14924 13716
rect 11940 13676 11946 13688
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15470 13676 15476 13728
rect 15528 13716 15534 13728
rect 16022 13716 16028 13728
rect 15528 13688 16028 13716
rect 15528 13676 15534 13688
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 16758 13676 16764 13728
rect 16816 13676 16822 13728
rect 18064 13716 18092 13815
rect 18322 13716 18328 13728
rect 18064 13688 18328 13716
rect 18322 13676 18328 13688
rect 18380 13716 18386 13728
rect 18984 13716 19012 13824
rect 19150 13744 19156 13796
rect 19208 13784 19214 13796
rect 19720 13784 19748 13824
rect 19978 13812 19984 13864
rect 20036 13852 20042 13864
rect 21560 13852 21588 13880
rect 20036 13824 21588 13852
rect 22833 13855 22891 13861
rect 20036 13812 20042 13824
rect 22833 13821 22845 13855
rect 22879 13821 22891 13855
rect 23032 13852 23060 13883
rect 23198 13880 23204 13932
rect 23256 13880 23262 13932
rect 23474 13880 23480 13932
rect 23532 13880 23538 13932
rect 25792 13864 25820 14016
rect 23566 13852 23572 13864
rect 23032 13824 23572 13852
rect 22833 13815 22891 13821
rect 22186 13784 22192 13796
rect 19208 13756 19656 13784
rect 19720 13756 22192 13784
rect 19208 13744 19214 13756
rect 18380 13688 19012 13716
rect 18380 13676 18386 13688
rect 19058 13676 19064 13728
rect 19116 13676 19122 13728
rect 19518 13676 19524 13728
rect 19576 13676 19582 13728
rect 19628 13716 19656 13756
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 22848 13784 22876 13815
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 25774 13812 25780 13864
rect 25832 13812 25838 13864
rect 23014 13784 23020 13796
rect 22848 13756 23020 13784
rect 23014 13744 23020 13756
rect 23072 13744 23078 13796
rect 23477 13787 23535 13793
rect 23477 13753 23489 13787
rect 23523 13753 23535 13787
rect 23477 13747 23535 13753
rect 22094 13716 22100 13728
rect 19628 13688 22100 13716
rect 22094 13676 22100 13688
rect 22152 13676 22158 13728
rect 23290 13676 23296 13728
rect 23348 13716 23354 13728
rect 23492 13716 23520 13747
rect 23348 13688 23520 13716
rect 23348 13676 23354 13688
rect 24394 13676 24400 13728
rect 24452 13676 24458 13728
rect 1104 13626 24840 13648
rect 1104 13574 3917 13626
rect 3969 13574 3981 13626
rect 4033 13574 4045 13626
rect 4097 13574 4109 13626
rect 4161 13574 4173 13626
rect 4225 13574 9851 13626
rect 9903 13574 9915 13626
rect 9967 13574 9979 13626
rect 10031 13574 10043 13626
rect 10095 13574 10107 13626
rect 10159 13574 15785 13626
rect 15837 13574 15849 13626
rect 15901 13574 15913 13626
rect 15965 13574 15977 13626
rect 16029 13574 16041 13626
rect 16093 13574 21719 13626
rect 21771 13574 21783 13626
rect 21835 13574 21847 13626
rect 21899 13574 21911 13626
rect 21963 13574 21975 13626
rect 22027 13574 24840 13626
rect 1104 13552 24840 13574
rect 1210 13472 1216 13524
rect 1268 13512 1274 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 1268 13484 2697 13512
rect 1268 13472 1274 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 2685 13475 2743 13481
rect 3237 13515 3295 13521
rect 3237 13481 3249 13515
rect 3283 13481 3295 13515
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 3237 13475 3295 13481
rect 3804 13484 11621 13512
rect 1302 13404 1308 13456
rect 1360 13444 1366 13456
rect 3252 13444 3280 13475
rect 1360 13416 3280 13444
rect 1360 13404 1366 13416
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 1765 13379 1823 13385
rect 1765 13376 1777 13379
rect 1452 13348 1777 13376
rect 1452 13336 1458 13348
rect 1765 13345 1777 13348
rect 1811 13345 1823 13379
rect 1765 13339 1823 13345
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 3804 13376 3832 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 13446 13512 13452 13524
rect 11609 13475 11667 13481
rect 12544 13484 13452 13512
rect 5074 13404 5080 13456
rect 5132 13444 5138 13456
rect 5718 13444 5724 13456
rect 5132 13416 5724 13444
rect 5132 13404 5138 13416
rect 5718 13404 5724 13416
rect 5776 13404 5782 13456
rect 5902 13404 5908 13456
rect 5960 13404 5966 13456
rect 8386 13404 8392 13456
rect 8444 13444 8450 13456
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 8444 13416 9321 13444
rect 8444 13404 8450 13416
rect 9309 13413 9321 13416
rect 9355 13413 9367 13447
rect 9309 13407 9367 13413
rect 9490 13404 9496 13456
rect 9548 13444 9554 13456
rect 9858 13444 9864 13456
rect 9548 13416 9864 13444
rect 9548 13404 9554 13416
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 10226 13404 10232 13456
rect 10284 13404 10290 13456
rect 10318 13404 10324 13456
rect 10376 13444 10382 13456
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 10376 13416 10425 13444
rect 10376 13404 10382 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 5920 13376 5948 13404
rect 6086 13376 6092 13388
rect 2188 13348 3832 13376
rect 5460 13348 6092 13376
rect 2188 13336 2194 13348
rect 1486 13268 1492 13320
rect 1544 13268 1550 13320
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 3326 13308 3332 13320
rect 2087 13280 3332 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 2409 13243 2467 13249
rect 2409 13209 2421 13243
rect 2455 13209 2467 13243
rect 2409 13203 2467 13209
rect 2424 13172 2452 13203
rect 2590 13200 2596 13252
rect 2648 13200 2654 13252
rect 3142 13200 3148 13252
rect 3200 13200 3206 13252
rect 3804 13240 3832 13271
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 4063 13311 4121 13317
rect 4063 13308 4075 13311
rect 4028 13280 4075 13308
rect 4028 13268 4034 13280
rect 4063 13277 4075 13280
rect 4109 13277 4121 13311
rect 4063 13271 4121 13277
rect 5460 13240 5488 13348
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9180 13348 9965 13376
rect 9180 13336 9186 13348
rect 9953 13345 9965 13348
rect 9999 13376 10011 13379
rect 10134 13376 10140 13388
rect 9999 13348 10140 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10244 13376 10272 13404
rect 10827 13379 10885 13385
rect 10827 13376 10839 13379
rect 10244 13348 10839 13376
rect 10827 13345 10839 13348
rect 10873 13376 10885 13379
rect 12544 13376 12572 13484
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 13630 13472 13636 13524
rect 13688 13472 13694 13524
rect 16485 13515 16543 13521
rect 15488 13484 16160 13512
rect 10873 13348 12572 13376
rect 10873 13345 10885 13348
rect 10827 13339 10885 13345
rect 13630 13336 13636 13388
rect 13688 13376 13694 13388
rect 13906 13376 13912 13388
rect 13688 13348 13912 13376
rect 13688 13336 13694 13348
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 15488 13385 15516 13484
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 16132 13376 16160 13484
rect 16485 13481 16497 13515
rect 16531 13512 16543 13515
rect 16850 13512 16856 13524
rect 16531 13484 16856 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 18564 13484 18613 13512
rect 18564 13472 18570 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 20806 13512 20812 13524
rect 18601 13475 18659 13481
rect 18708 13484 20812 13512
rect 18708 13453 18736 13484
rect 20806 13472 20812 13484
rect 20864 13472 20870 13524
rect 22281 13515 22339 13521
rect 22281 13481 22293 13515
rect 22327 13512 22339 13515
rect 22554 13512 22560 13524
rect 22327 13484 22560 13512
rect 22327 13481 22339 13484
rect 22281 13475 22339 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 22649 13515 22707 13521
rect 22649 13481 22661 13515
rect 22695 13512 22707 13515
rect 23474 13512 23480 13524
rect 22695 13484 23480 13512
rect 22695 13481 22707 13484
rect 22649 13475 22707 13481
rect 23474 13472 23480 13484
rect 23532 13472 23538 13524
rect 18693 13447 18751 13453
rect 18693 13413 18705 13447
rect 18739 13413 18751 13447
rect 19978 13444 19984 13456
rect 18693 13407 18751 13413
rect 19628 13416 19984 13444
rect 16132 13348 16804 13376
rect 15473 13339 15531 13345
rect 16776 13320 16804 13348
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17678 13376 17684 13388
rect 17184 13348 17684 13376
rect 17184 13336 17190 13348
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 18785 13379 18843 13385
rect 18785 13345 18797 13379
rect 18831 13376 18843 13379
rect 19518 13376 19524 13388
rect 18831 13348 19524 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 5902 13308 5908 13320
rect 5592 13280 5908 13308
rect 5592 13268 5598 13280
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 9815 13280 9849 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 3804 13212 5488 13240
rect 8018 13200 8024 13252
rect 8076 13240 8082 13252
rect 9784 13240 9812 13271
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 11882 13268 11888 13320
rect 11940 13268 11946 13320
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12250 13308 12256 13320
rect 12032 13280 12256 13308
rect 12032 13268 12038 13280
rect 12250 13268 12256 13280
rect 12308 13268 12314 13320
rect 12621 13311 12679 13317
rect 12621 13277 12633 13311
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 12895 13311 12953 13317
rect 12895 13277 12907 13311
rect 12941 13308 12953 13311
rect 14366 13308 14372 13320
rect 12941 13280 14372 13308
rect 12941 13277 12953 13280
rect 12895 13271 12953 13277
rect 9950 13240 9956 13252
rect 8076 13212 9956 13240
rect 8076 13200 8082 13212
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 11900 13240 11928 13268
rect 12636 13240 12664 13271
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 14642 13268 14648 13320
rect 14700 13308 14706 13320
rect 15286 13308 15292 13320
rect 14700 13280 15292 13308
rect 14700 13268 14706 13280
rect 15286 13268 15292 13280
rect 15344 13308 15350 13320
rect 15715 13311 15773 13317
rect 15715 13308 15727 13311
rect 15344 13280 15727 13308
rect 15344 13268 15350 13280
rect 15715 13277 15727 13280
rect 15761 13277 15773 13311
rect 15715 13271 15773 13277
rect 16758 13268 16764 13320
rect 16816 13308 16822 13320
rect 18509 13311 18567 13317
rect 16816 13280 18350 13308
rect 16816 13268 16822 13280
rect 17678 13240 17684 13252
rect 11900 13212 12664 13240
rect 13096 13212 17684 13240
rect 2774 13172 2780 13184
rect 2424 13144 2780 13172
rect 2774 13132 2780 13144
rect 2832 13132 2838 13184
rect 4430 13132 4436 13184
rect 4488 13172 4494 13184
rect 4801 13175 4859 13181
rect 4801 13172 4813 13175
rect 4488 13144 4813 13172
rect 4488 13132 4494 13144
rect 4801 13141 4813 13144
rect 4847 13141 4859 13175
rect 4801 13135 4859 13141
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 6270 13172 6276 13184
rect 5408 13144 6276 13172
rect 5408 13132 5414 13144
rect 6270 13132 6276 13144
rect 6328 13132 6334 13184
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 13096 13172 13124 13212
rect 17678 13200 17684 13212
rect 17736 13240 17742 13252
rect 18230 13240 18236 13252
rect 17736 13212 18236 13240
rect 17736 13200 17742 13212
rect 18230 13200 18236 13212
rect 18288 13200 18294 13252
rect 18322 13240 18350 13280
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 19058 13308 19064 13320
rect 18555 13280 19064 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 19058 13268 19064 13280
rect 19116 13268 19122 13320
rect 19518 13240 19524 13252
rect 18322 13212 19524 13240
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 7340 13144 13124 13172
rect 7340 13132 7346 13144
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 14734 13172 14740 13184
rect 13228 13144 14740 13172
rect 13228 13132 13234 13144
rect 14734 13132 14740 13144
rect 14792 13132 14798 13184
rect 18046 13132 18052 13184
rect 18104 13172 18110 13184
rect 19628 13172 19656 13416
rect 19978 13404 19984 13416
rect 20036 13404 20042 13456
rect 21266 13404 21272 13456
rect 21324 13444 21330 13456
rect 22370 13444 22376 13456
rect 21324 13416 22376 13444
rect 21324 13404 21330 13416
rect 22370 13404 22376 13416
rect 22428 13444 22434 13456
rect 22428 13416 22876 13444
rect 22428 13404 22434 13416
rect 22848 13385 22876 13416
rect 20441 13379 20499 13385
rect 20441 13376 20453 13379
rect 19904 13348 20116 13376
rect 19904 13317 19932 13348
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 20088 13308 20116 13348
rect 20272 13348 20453 13376
rect 20272 13308 20300 13348
rect 20441 13345 20453 13348
rect 20487 13345 20499 13379
rect 20441 13339 20499 13345
rect 22833 13379 22891 13385
rect 22833 13345 22845 13379
rect 22879 13345 22891 13379
rect 22833 13339 22891 13345
rect 20088 13280 20300 13308
rect 19889 13271 19947 13277
rect 19720 13240 19748 13271
rect 20346 13268 20352 13320
rect 20404 13268 20410 13320
rect 20530 13268 20536 13320
rect 20588 13310 20594 13320
rect 20625 13311 20683 13317
rect 20625 13310 20637 13311
rect 20588 13282 20637 13310
rect 20588 13268 20594 13282
rect 20625 13277 20637 13282
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 21542 13308 21548 13320
rect 20855 13280 21548 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 21542 13268 21548 13280
rect 21600 13268 21606 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 19720 13212 19923 13240
rect 18104 13144 19656 13172
rect 19895 13172 19923 13212
rect 20162 13200 20168 13252
rect 20220 13200 20226 13252
rect 20257 13243 20315 13249
rect 20257 13209 20269 13243
rect 20303 13209 20315 13243
rect 20717 13243 20775 13249
rect 20717 13240 20729 13243
rect 20257 13203 20315 13209
rect 20456 13212 20729 13240
rect 19978 13172 19984 13184
rect 19895 13144 19984 13172
rect 18104 13132 18110 13144
rect 19978 13132 19984 13144
rect 20036 13132 20042 13184
rect 20272 13172 20300 13203
rect 20456 13172 20484 13212
rect 20717 13209 20729 13212
rect 20763 13209 20775 13243
rect 22480 13240 22508 13271
rect 22554 13268 22560 13320
rect 22612 13268 22618 13320
rect 23100 13243 23158 13249
rect 22480 13212 22784 13240
rect 20717 13203 20775 13209
rect 20272 13144 20484 13172
rect 22756 13172 22784 13212
rect 23100 13209 23112 13243
rect 23146 13240 23158 13243
rect 23474 13240 23480 13252
rect 23146 13212 23480 13240
rect 23146 13209 23158 13212
rect 23100 13203 23158 13209
rect 23474 13200 23480 13212
rect 23532 13200 23538 13252
rect 24213 13175 24271 13181
rect 24213 13172 24225 13175
rect 22756 13144 24225 13172
rect 24213 13141 24225 13144
rect 24259 13141 24271 13175
rect 24213 13135 24271 13141
rect 1104 13082 25000 13104
rect 1104 13030 6884 13082
rect 6936 13030 6948 13082
rect 7000 13030 7012 13082
rect 7064 13030 7076 13082
rect 7128 13030 7140 13082
rect 7192 13030 12818 13082
rect 12870 13030 12882 13082
rect 12934 13030 12946 13082
rect 12998 13030 13010 13082
rect 13062 13030 13074 13082
rect 13126 13030 18752 13082
rect 18804 13030 18816 13082
rect 18868 13030 18880 13082
rect 18932 13030 18944 13082
rect 18996 13030 19008 13082
rect 19060 13030 24686 13082
rect 24738 13030 24750 13082
rect 24802 13030 24814 13082
rect 24866 13030 24878 13082
rect 24930 13030 24942 13082
rect 24994 13030 25000 13082
rect 1104 13008 25000 13030
rect 1762 12928 1768 12980
rect 1820 12928 1826 12980
rect 6362 12968 6368 12980
rect 2608 12940 6368 12968
rect 2608 12851 2636 12940
rect 6362 12928 6368 12940
rect 6420 12968 6426 12980
rect 7282 12968 7288 12980
rect 6420 12940 7288 12968
rect 6420 12928 6426 12940
rect 6104 12872 6500 12900
rect 2591 12845 2649 12851
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2222 12832 2228 12844
rect 1719 12804 2228 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 2591 12811 2603 12845
rect 2637 12811 2649 12845
rect 6104 12844 6132 12872
rect 2591 12805 2649 12811
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3602 12832 3608 12844
rect 3292 12804 3608 12832
rect 3292 12792 3298 12804
rect 3602 12792 3608 12804
rect 3660 12832 3666 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3660 12804 3709 12832
rect 3660 12792 3666 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 6086 12792 6092 12844
rect 6144 12792 6150 12844
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12832 6423 12835
rect 6472 12832 6500 12872
rect 6622 12841 6650 12940
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7926 12968 7932 12980
rect 7432 12940 7932 12968
rect 7432 12928 7438 12940
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9122 12968 9128 12980
rect 8220 12940 9128 12968
rect 6411 12804 6500 12832
rect 6607 12835 6665 12841
rect 6411 12801 6423 12804
rect 6365 12795 6423 12801
rect 6607 12801 6619 12835
rect 6653 12801 6665 12835
rect 6607 12795 6665 12801
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 8220 12841 8248 12940
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 9490 12928 9496 12980
rect 9548 12968 9554 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9548 12940 9873 12968
rect 9548 12928 9554 12940
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 9861 12931 9919 12937
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 11020 12940 11069 12968
rect 11020 12928 11026 12940
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 11057 12931 11115 12937
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 20162 12968 20168 12980
rect 11664 12940 20168 12968
rect 11664 12928 11670 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20993 12971 21051 12977
rect 20993 12937 21005 12971
rect 21039 12968 21051 12971
rect 22189 12971 22247 12977
rect 21039 12940 21588 12968
rect 21039 12937 21051 12940
rect 20993 12931 21051 12937
rect 10502 12860 10508 12912
rect 10560 12860 10566 12912
rect 19150 12900 19156 12912
rect 11256 12872 19156 12900
rect 8205 12835 8263 12841
rect 6788 12804 7512 12832
rect 6788 12792 6794 12804
rect 1762 12724 1768 12776
rect 1820 12764 1826 12776
rect 2314 12764 2320 12776
rect 1820 12736 2320 12764
rect 1820 12724 1826 12736
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3786 12764 3792 12776
rect 3252 12736 3792 12764
rect 3252 12708 3280 12736
rect 3786 12724 3792 12736
rect 3844 12764 3850 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3844 12736 3893 12764
rect 3844 12724 3850 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4430 12764 4436 12776
rect 4387 12736 4436 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 4614 12724 4620 12776
rect 4672 12773 4678 12776
rect 4672 12767 4693 12773
rect 4681 12733 4693 12767
rect 4672 12727 4693 12733
rect 4672 12724 4678 12727
rect 4731 12724 4737 12776
rect 4789 12724 4795 12776
rect 3234 12656 3240 12708
rect 3292 12656 3298 12708
rect 3326 12588 3332 12640
rect 3384 12588 3390 12640
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 3844 12600 5549 12628
rect 3844 12588 3850 12600
rect 5537 12597 5549 12600
rect 5583 12597 5595 12631
rect 5537 12591 5595 12597
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 7377 12631 7435 12637
rect 7377 12628 7389 12631
rect 6144 12600 7389 12628
rect 6144 12588 6150 12600
rect 7377 12597 7389 12600
rect 7423 12597 7435 12631
rect 7484 12628 7512 12804
rect 8205 12801 8217 12835
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10045 12835 10103 12841
rect 10045 12832 10057 12835
rect 9916 12804 10057 12832
rect 9916 12792 9922 12804
rect 10045 12801 10057 12804
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10319 12835 10377 12841
rect 10319 12801 10331 12835
rect 10365 12832 10377 12835
rect 10520 12832 10548 12860
rect 11256 12832 11284 12872
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19978 12900 19984 12912
rect 19260 12872 19984 12900
rect 10365 12804 10548 12832
rect 10704 12804 11284 12832
rect 10365 12801 10377 12804
rect 10319 12795 10377 12801
rect 7834 12724 7840 12776
rect 7892 12724 7898 12776
rect 8018 12724 8024 12776
rect 8076 12724 8082 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8956 12764 8984 12792
rect 8444 12736 8984 12764
rect 8444 12724 8450 12736
rect 9030 12724 9036 12776
rect 9088 12773 9094 12776
rect 9088 12767 9116 12773
rect 9104 12733 9116 12767
rect 9088 12727 9116 12733
rect 9088 12724 9094 12727
rect 7852 12696 7880 12724
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 7852 12668 8677 12696
rect 8665 12665 8677 12668
rect 8711 12665 8723 12699
rect 8665 12659 8723 12665
rect 10704 12628 10732 12804
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11974 12832 11980 12844
rect 11388 12804 11980 12832
rect 11388 12792 11394 12804
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12066 12792 12072 12844
rect 12124 12832 12130 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 12124 12804 13921 12832
rect 12124 12792 12130 12804
rect 13909 12801 13921 12804
rect 13955 12801 13967 12835
rect 13909 12795 13967 12801
rect 14183 12835 14241 12841
rect 14183 12801 14195 12835
rect 14229 12832 14241 12835
rect 14826 12832 14832 12844
rect 14229 12804 14832 12832
rect 14229 12801 14241 12804
rect 14183 12795 14241 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 17034 12841 17040 12844
rect 17003 12835 17040 12841
rect 17003 12832 17015 12835
rect 14936 12804 17015 12832
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 14936 12764 14964 12804
rect 17003 12801 17015 12804
rect 17003 12795 17040 12801
rect 17034 12792 17040 12795
rect 17092 12792 17098 12844
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 18475 12835 18533 12841
rect 18475 12832 18487 12835
rect 17736 12804 18487 12832
rect 17736 12792 17742 12804
rect 18475 12801 18487 12804
rect 18521 12801 18533 12835
rect 18475 12795 18533 12801
rect 11701 12727 11759 12733
rect 14568 12736 14964 12764
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11606 12696 11612 12708
rect 11296 12668 11612 12696
rect 11296 12656 11302 12668
rect 11606 12656 11612 12668
rect 11664 12696 11670 12708
rect 11716 12696 11744 12727
rect 11664 12668 11744 12696
rect 11664 12656 11670 12668
rect 7484 12600 10732 12628
rect 11716 12628 11744 12668
rect 12636 12668 14044 12696
rect 11974 12628 11980 12640
rect 11716 12600 11980 12628
rect 7377 12591 7435 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 12636 12628 12664 12668
rect 12124 12600 12664 12628
rect 12124 12588 12130 12600
rect 12710 12588 12716 12640
rect 12768 12588 12774 12640
rect 14016 12628 14044 12668
rect 14568 12628 14596 12736
rect 16114 12724 16120 12776
rect 16172 12764 16178 12776
rect 16761 12767 16819 12773
rect 16761 12764 16773 12767
rect 16172 12736 16773 12764
rect 16172 12724 16178 12736
rect 16761 12733 16773 12736
rect 16807 12733 16819 12767
rect 16761 12727 16819 12733
rect 18233 12767 18291 12773
rect 18233 12733 18245 12767
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18248 12696 18276 12727
rect 19260 12705 19288 12872
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 20530 12900 20536 12912
rect 20272 12872 20536 12900
rect 19610 12792 19616 12844
rect 19668 12792 19674 12844
rect 19880 12835 19938 12841
rect 19880 12801 19892 12835
rect 19926 12832 19938 12835
rect 20272 12832 20300 12872
rect 20530 12860 20536 12872
rect 20588 12900 20594 12912
rect 20588 12872 21312 12900
rect 20588 12860 20594 12872
rect 21284 12841 21312 12872
rect 21560 12841 21588 12940
rect 22189 12937 22201 12971
rect 22235 12968 22247 12971
rect 22462 12968 22468 12980
rect 22235 12940 22468 12968
rect 22235 12937 22247 12940
rect 22189 12931 22247 12937
rect 22462 12928 22468 12940
rect 22520 12928 22526 12980
rect 22830 12928 22836 12980
rect 22888 12928 22894 12980
rect 23385 12971 23443 12977
rect 23385 12937 23397 12971
rect 23431 12968 23443 12971
rect 23566 12968 23572 12980
rect 23431 12940 23572 12968
rect 23431 12937 23443 12940
rect 23385 12931 23443 12937
rect 23566 12928 23572 12940
rect 23624 12928 23630 12980
rect 22848 12900 22876 12928
rect 22664 12872 22876 12900
rect 23937 12903 23995 12909
rect 22664 12871 22692 12872
rect 22631 12865 22692 12871
rect 19926 12804 20300 12832
rect 21269 12835 21327 12841
rect 19926 12801 19938 12804
rect 19880 12795 19938 12801
rect 21269 12801 21281 12835
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 21545 12835 21603 12841
rect 21545 12801 21557 12835
rect 21591 12801 21603 12835
rect 21545 12795 21603 12801
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12801 22155 12835
rect 22097 12795 22155 12801
rect 20990 12724 20996 12776
rect 21048 12764 21054 12776
rect 22112 12764 22140 12795
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 22244 12804 22385 12832
rect 22244 12792 22250 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22462 12802 22468 12854
rect 22520 12832 22526 12854
rect 22631 12832 22643 12865
rect 22520 12831 22643 12832
rect 22677 12831 22692 12865
rect 23937 12869 23949 12903
rect 23983 12900 23995 12903
rect 24486 12900 24492 12912
rect 23983 12872 24492 12900
rect 23983 12869 23995 12872
rect 23937 12863 23995 12869
rect 24486 12860 24492 12872
rect 24544 12860 24550 12912
rect 22520 12804 22692 12831
rect 22520 12802 22526 12804
rect 22373 12795 22431 12801
rect 21048 12736 22140 12764
rect 21048 12724 21054 12736
rect 19245 12699 19303 12705
rect 18248 12668 18368 12696
rect 18340 12640 18368 12668
rect 19245 12665 19257 12699
rect 19291 12665 19303 12699
rect 19245 12659 19303 12665
rect 21361 12699 21419 12705
rect 21361 12665 21373 12699
rect 21407 12696 21419 12699
rect 21542 12696 21548 12708
rect 21407 12668 21548 12696
rect 21407 12665 21419 12668
rect 21361 12659 21419 12665
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 14016 12600 14596 12628
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 14921 12631 14979 12637
rect 14921 12628 14933 12631
rect 14700 12600 14933 12628
rect 14700 12588 14706 12600
rect 14921 12597 14933 12600
rect 14967 12597 14979 12631
rect 14921 12591 14979 12597
rect 17770 12588 17776 12640
rect 17828 12588 17834 12640
rect 18322 12588 18328 12640
rect 18380 12588 18386 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20404 12600 21097 12628
rect 20404 12588 20410 12600
rect 21085 12597 21097 12600
rect 21131 12597 21143 12631
rect 21085 12591 21143 12597
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 22094 12628 22100 12640
rect 21232 12600 22100 12628
rect 21232 12588 21238 12600
rect 22094 12588 22100 12600
rect 22152 12588 22158 12640
rect 24210 12588 24216 12640
rect 24268 12588 24274 12640
rect 1104 12538 24840 12560
rect 1104 12486 3917 12538
rect 3969 12486 3981 12538
rect 4033 12486 4045 12538
rect 4097 12486 4109 12538
rect 4161 12486 4173 12538
rect 4225 12486 9851 12538
rect 9903 12486 9915 12538
rect 9967 12486 9979 12538
rect 10031 12486 10043 12538
rect 10095 12486 10107 12538
rect 10159 12486 15785 12538
rect 15837 12486 15849 12538
rect 15901 12486 15913 12538
rect 15965 12486 15977 12538
rect 16029 12486 16041 12538
rect 16093 12486 21719 12538
rect 21771 12486 21783 12538
rect 21835 12486 21847 12538
rect 21899 12486 21911 12538
rect 21963 12486 21975 12538
rect 22027 12486 24840 12538
rect 1104 12464 24840 12486
rect 3602 12384 3608 12436
rect 3660 12424 3666 12436
rect 4157 12427 4215 12433
rect 3660 12396 3740 12424
rect 3660 12384 3666 12396
rect 3712 12356 3740 12396
rect 4157 12393 4169 12427
rect 4203 12424 4215 12427
rect 4246 12424 4252 12436
rect 4203 12396 4252 12424
rect 4203 12393 4215 12396
rect 4157 12387 4215 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5350 12424 5356 12436
rect 4764 12396 5356 12424
rect 4764 12384 4770 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 6914 12424 6920 12436
rect 6564 12396 6920 12424
rect 4430 12356 4436 12368
rect 3712 12328 4436 12356
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 4816 12328 5672 12356
rect 934 12248 940 12300
rect 992 12288 998 12300
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 992 12260 1777 12288
rect 992 12248 998 12260
rect 1765 12257 1777 12260
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2038 12288 2044 12300
rect 1995 12260 2044 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2406 12248 2412 12300
rect 2464 12248 2470 12300
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2961 12291 3019 12297
rect 2832 12248 2845 12288
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3326 12288 3332 12300
rect 3007 12260 3332 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 3605 12291 3663 12297
rect 3605 12257 3617 12291
rect 3651 12288 3663 12291
rect 4246 12288 4252 12300
rect 3651 12260 4252 12288
rect 3651 12257 3663 12260
rect 3605 12251 3663 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 2682 12180 2688 12232
rect 2740 12180 2746 12232
rect 2817 12229 2845 12248
rect 4816 12232 4844 12328
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 2817 12223 2881 12229
rect 2817 12192 2835 12223
rect 2823 12189 2835 12192
rect 2869 12189 2881 12223
rect 2823 12183 2881 12189
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 3881 12223 3939 12229
rect 3881 12220 3893 12223
rect 3752 12192 3893 12220
rect 3752 12180 3758 12192
rect 3881 12189 3893 12192
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 4154 12180 4160 12232
rect 4212 12220 4218 12232
rect 4212 12192 4568 12220
rect 4212 12180 4218 12192
rect 4433 12155 4491 12161
rect 4433 12152 4445 12155
rect 3528 12124 4445 12152
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 3528 12084 3556 12124
rect 4433 12121 4445 12124
rect 4479 12121 4491 12155
rect 4540 12152 4568 12192
rect 4798 12180 4804 12232
rect 4856 12180 4862 12232
rect 4908 12220 4936 12251
rect 5534 12248 5540 12300
rect 5592 12248 5598 12300
rect 5644 12288 5672 12328
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5644 12260 5825 12288
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 5951 12291 6009 12297
rect 5951 12257 5963 12291
rect 5997 12288 6009 12291
rect 6564 12288 6592 12396
rect 6914 12384 6920 12396
rect 6972 12384 6978 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7432 12396 7604 12424
rect 7432 12384 7438 12396
rect 5997 12260 6592 12288
rect 5997 12257 6009 12260
rect 5951 12251 6009 12257
rect 6822 12248 6828 12300
rect 6880 12248 6886 12300
rect 7466 12248 7472 12300
rect 7524 12248 7530 12300
rect 7576 12288 7604 12396
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 7984 12396 8677 12424
rect 7984 12384 7990 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 8665 12387 8723 12393
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 15565 12427 15623 12433
rect 15565 12424 15577 12427
rect 15528 12396 15577 12424
rect 15528 12384 15534 12396
rect 15565 12393 15577 12396
rect 15611 12393 15623 12427
rect 20990 12424 20996 12436
rect 15565 12387 15623 12393
rect 19904 12396 20996 12424
rect 8478 12316 8484 12368
rect 8536 12316 8542 12368
rect 15580 12356 15608 12387
rect 15580 12328 17172 12356
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7576 12260 7757 12288
rect 7745 12257 7757 12260
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 7883 12291 7941 12297
rect 7883 12257 7895 12291
rect 7929 12288 7941 12291
rect 8496 12288 8524 12316
rect 7929 12260 8524 12288
rect 12532 12300 12584 12306
rect 7929 12257 7941 12260
rect 7883 12251 7941 12257
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 13964 12260 14122 12288
rect 13964 12248 13970 12260
rect 17034 12248 17040 12300
rect 17092 12248 17098 12300
rect 17144 12288 17172 12328
rect 17430 12291 17488 12297
rect 17430 12288 17442 12291
rect 17144 12260 17442 12288
rect 17430 12257 17442 12260
rect 17476 12257 17488 12291
rect 17430 12251 17488 12257
rect 17586 12248 17592 12300
rect 17644 12248 17650 12300
rect 18322 12248 18328 12300
rect 18380 12288 18386 12300
rect 18598 12288 18604 12300
rect 18380 12260 18604 12288
rect 18380 12248 18386 12260
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 19904 12297 19932 12396
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 22649 12427 22707 12433
rect 22649 12393 22661 12427
rect 22695 12424 22707 12427
rect 24121 12427 24179 12433
rect 22695 12396 23520 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 23293 12359 23351 12365
rect 23293 12325 23305 12359
rect 23339 12325 23351 12359
rect 23293 12319 23351 12325
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12257 19947 12291
rect 19889 12251 19947 12257
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 12532 12242 12584 12248
rect 4982 12220 4988 12232
rect 4908 12192 4988 12220
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5092 12152 5120 12183
rect 6086 12180 6092 12232
rect 6144 12180 6150 12232
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7024 12152 7052 12183
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12220 11943 12223
rect 12710 12220 12716 12232
rect 11931 12210 12480 12220
rect 12636 12210 12716 12220
rect 11931 12192 12716 12210
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 12452 12182 12664 12192
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 14366 12220 14372 12232
rect 12860 12192 14372 12220
rect 12860 12180 12866 12192
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14642 12180 14648 12232
rect 14700 12180 14706 12232
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 15378 12180 15384 12232
rect 15436 12180 15442 12232
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 15528 12192 16405 12220
rect 15528 12180 15534 12192
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16540 12192 16589 12220
rect 16540 12180 16546 12192
rect 16577 12189 16589 12192
rect 16623 12220 16635 12223
rect 16758 12220 16764 12232
rect 16623 12192 16764 12220
rect 16623 12189 16635 12192
rect 16577 12183 16635 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 20162 12229 20168 12232
rect 20131 12223 20168 12229
rect 20131 12189 20143 12223
rect 20131 12183 20168 12189
rect 20162 12180 20168 12183
rect 20220 12180 20226 12232
rect 20530 12180 20536 12232
rect 20588 12220 20594 12232
rect 20806 12220 20812 12232
rect 20588 12192 20812 12220
rect 20588 12180 20594 12192
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12220 23259 12223
rect 23308 12220 23336 12319
rect 23492 12229 23520 12396
rect 24121 12393 24133 12427
rect 24167 12424 24179 12427
rect 25130 12424 25136 12436
rect 24167 12396 25136 12424
rect 24167 12393 24179 12396
rect 24121 12387 24179 12393
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 23753 12359 23811 12365
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 25222 12356 25228 12368
rect 23799 12328 25228 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 25222 12316 25228 12328
rect 25280 12316 25286 12368
rect 23842 12288 23848 12300
rect 23584 12260 23848 12288
rect 23584 12229 23612 12260
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 23247 12192 23336 12220
rect 23477 12223 23535 12229
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 23477 12189 23489 12223
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 4540 12124 5120 12152
rect 4433 12115 4491 12121
rect 2004 12056 3556 12084
rect 2004 12044 2010 12056
rect 3786 12044 3792 12096
rect 3844 12084 3850 12096
rect 4525 12087 4583 12093
rect 4525 12084 4537 12087
rect 3844 12056 4537 12084
rect 3844 12044 3850 12056
rect 4525 12053 4537 12056
rect 4571 12053 4583 12087
rect 5092 12084 5120 12124
rect 6564 12124 7052 12152
rect 6086 12084 6092 12096
rect 5092 12056 6092 12084
rect 4525 12047 4583 12053
rect 6086 12044 6092 12056
rect 6144 12084 6150 12096
rect 6564 12084 6592 12124
rect 6144 12056 6592 12084
rect 6144 12044 6150 12056
rect 6730 12044 6736 12096
rect 6788 12044 6794 12096
rect 7024 12084 7052 12124
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 11793 12155 11851 12161
rect 9088 12124 11744 12152
rect 9088 12112 9094 12124
rect 9674 12084 9680 12096
rect 7024 12056 9680 12084
rect 9674 12044 9680 12056
rect 9732 12084 9738 12096
rect 11238 12084 11244 12096
rect 9732 12056 11244 12084
rect 9732 12044 9738 12056
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 11606 12084 11612 12096
rect 11563 12056 11612 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11716 12084 11744 12124
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 11974 12152 11980 12164
rect 11839 12124 11980 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 11974 12112 11980 12124
rect 12032 12112 12038 12164
rect 12158 12112 12164 12164
rect 12216 12152 12222 12164
rect 12253 12155 12311 12161
rect 12253 12152 12265 12155
rect 12216 12124 12265 12152
rect 12216 12112 12222 12124
rect 12253 12121 12265 12124
rect 12299 12121 12311 12155
rect 12253 12115 12311 12121
rect 12406 12124 12848 12152
rect 12406 12084 12434 12124
rect 11716 12056 12434 12084
rect 12618 12044 12624 12096
rect 12676 12044 12682 12096
rect 12820 12093 12848 12124
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 14240 12124 14565 12152
rect 14240 12112 14246 12124
rect 14553 12121 14565 12124
rect 14599 12152 14611 12155
rect 14752 12152 14780 12180
rect 14599 12124 14780 12152
rect 15013 12155 15071 12161
rect 14599 12121 14611 12124
rect 14553 12115 14611 12121
rect 15013 12121 15025 12155
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13722 12084 13728 12096
rect 13228 12056 13728 12084
rect 13228 12044 13234 12056
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 14274 12044 14280 12096
rect 14332 12044 14338 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14642 12084 14648 12096
rect 14424 12056 14648 12084
rect 14424 12044 14430 12056
rect 14642 12044 14648 12056
rect 14700 12084 14706 12096
rect 15028 12084 15056 12115
rect 14700 12056 15056 12084
rect 14700 12044 14706 12056
rect 15102 12044 15108 12096
rect 15160 12084 15166 12096
rect 15396 12093 15424 12180
rect 21542 12161 21548 12164
rect 21536 12152 21548 12161
rect 18064 12124 20760 12152
rect 21503 12124 21548 12152
rect 15381 12087 15439 12093
rect 15381 12084 15393 12087
rect 15160 12056 15393 12084
rect 15160 12044 15166 12056
rect 15381 12053 15393 12056
rect 15427 12053 15439 12087
rect 15381 12047 15439 12053
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 18064 12084 18092 12124
rect 20732 12096 20760 12124
rect 21536 12115 21548 12124
rect 21542 12112 21548 12115
rect 21600 12112 21606 12164
rect 23032 12152 23060 12183
rect 23658 12180 23664 12232
rect 23716 12220 23722 12232
rect 23937 12223 23995 12229
rect 23937 12220 23949 12223
rect 23716 12192 23949 12220
rect 23716 12180 23722 12192
rect 23937 12189 23949 12192
rect 23983 12189 23995 12223
rect 23937 12183 23995 12189
rect 22066 12124 23060 12152
rect 15804 12056 18092 12084
rect 15804 12044 15810 12056
rect 18230 12044 18236 12096
rect 18288 12044 18294 12096
rect 20714 12044 20720 12096
rect 20772 12044 20778 12096
rect 20901 12087 20959 12093
rect 20901 12053 20913 12087
rect 20947 12084 20959 12087
rect 21818 12084 21824 12096
rect 20947 12056 21824 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 21818 12044 21824 12056
rect 21876 12084 21882 12096
rect 22066 12084 22094 12124
rect 21876 12056 22094 12084
rect 21876 12044 21882 12056
rect 22830 12044 22836 12096
rect 22888 12044 22894 12096
rect 23106 12044 23112 12096
rect 23164 12044 23170 12096
rect 1104 11994 25000 12016
rect 1104 11942 6884 11994
rect 6936 11942 6948 11994
rect 7000 11942 7012 11994
rect 7064 11942 7076 11994
rect 7128 11942 7140 11994
rect 7192 11942 12818 11994
rect 12870 11942 12882 11994
rect 12934 11942 12946 11994
rect 12998 11942 13010 11994
rect 13062 11942 13074 11994
rect 13126 11942 18752 11994
rect 18804 11942 18816 11994
rect 18868 11942 18880 11994
rect 18932 11942 18944 11994
rect 18996 11942 19008 11994
rect 19060 11942 24686 11994
rect 24738 11942 24750 11994
rect 24802 11942 24814 11994
rect 24866 11942 24878 11994
rect 24930 11942 24942 11994
rect 24994 11942 25000 11994
rect 1104 11920 25000 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2464 11852 2881 11880
rect 2464 11840 2470 11852
rect 2869 11849 2881 11852
rect 2915 11849 2927 11883
rect 4154 11880 4160 11892
rect 2869 11843 2927 11849
rect 2976 11852 4160 11880
rect 2038 11772 2044 11824
rect 2096 11812 2102 11824
rect 2976 11812 3004 11852
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4525 11883 4583 11889
rect 4525 11849 4537 11883
rect 4571 11880 4583 11883
rect 4890 11880 4896 11892
rect 4571 11852 4896 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5905 11883 5963 11889
rect 5905 11880 5917 11883
rect 5592 11852 5917 11880
rect 5592 11840 5598 11852
rect 5905 11849 5917 11852
rect 5951 11849 5963 11883
rect 5905 11843 5963 11849
rect 6362 11840 6368 11892
rect 6420 11840 6426 11892
rect 7929 11883 7987 11889
rect 6472 11852 7328 11880
rect 2096 11784 3004 11812
rect 2096 11772 2102 11784
rect 3050 11772 3056 11824
rect 3108 11812 3114 11824
rect 3970 11812 3976 11824
rect 3108 11784 3556 11812
rect 3108 11772 3114 11784
rect 2131 11747 2189 11753
rect 2131 11713 2143 11747
rect 2177 11744 2189 11747
rect 2177 11716 3372 11744
rect 2177 11713 2189 11716
rect 2131 11707 2189 11713
rect 1762 11636 1768 11688
rect 1820 11676 1826 11688
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1820 11648 1869 11676
rect 1820 11636 1826 11648
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 2746 11580 3280 11608
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 2746 11540 2774 11580
rect 3252 11549 3280 11580
rect 1544 11512 2774 11540
rect 3237 11543 3295 11549
rect 1544 11500 1550 11512
rect 3237 11509 3249 11543
rect 3283 11509 3295 11543
rect 3344 11540 3372 11716
rect 3418 11704 3424 11756
rect 3476 11704 3482 11756
rect 3528 11753 3556 11784
rect 3896 11784 3976 11812
rect 3896 11774 3924 11784
rect 3804 11763 3924 11774
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 6380 11812 6408 11840
rect 5182 11784 6408 11812
rect 5182 11783 5210 11784
rect 5151 11777 5210 11783
rect 3787 11757 3924 11763
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11713 3571 11747
rect 3787 11723 3799 11757
rect 3833 11746 3924 11757
rect 3833 11723 3845 11746
rect 5151 11744 5163 11777
rect 3787 11717 3845 11723
rect 4448 11743 5163 11744
rect 5197 11743 5210 11777
rect 3513 11707 3571 11713
rect 4448 11716 5210 11743
rect 4448 11608 4476 11716
rect 4890 11636 4896 11688
rect 4948 11636 4954 11688
rect 4172 11580 4476 11608
rect 4172 11540 4200 11580
rect 3344 11512 4200 11540
rect 3237 11503 3295 11509
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 6472 11540 6500 11852
rect 7300 11812 7328 11852
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8018 11880 8024 11892
rect 7975 11852 8024 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 12434 11880 12440 11892
rect 12216 11852 12440 11880
rect 12216 11840 12222 11852
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 12526 11840 12532 11892
rect 12584 11840 12590 11892
rect 12820 11852 13860 11880
rect 12820 11812 12848 11852
rect 7300 11784 12848 11812
rect 13832 11812 13860 11852
rect 13906 11840 13912 11892
rect 13964 11840 13970 11892
rect 14936 11852 15148 11880
rect 14936 11812 14964 11852
rect 13832 11784 14964 11812
rect 15120 11812 15148 11852
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 15436 11852 15945 11880
rect 15436 11840 15442 11852
rect 15933 11849 15945 11852
rect 15979 11849 15991 11883
rect 15933 11843 15991 11849
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 17092 11852 17693 11880
rect 17092 11840 17098 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 21453 11883 21511 11889
rect 17681 11843 17739 11849
rect 18064 11852 18644 11880
rect 17862 11812 17868 11824
rect 15120 11784 17868 11812
rect 17862 11772 17868 11784
rect 17920 11772 17926 11824
rect 7191 11747 7249 11753
rect 7191 11713 7203 11747
rect 7237 11744 7249 11747
rect 7282 11744 7288 11756
rect 7237 11716 7288 11744
rect 7237 11713 7249 11716
rect 7191 11707 7249 11713
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 8570 11704 8576 11756
rect 8628 11744 8634 11756
rect 9030 11744 9036 11756
rect 8628 11716 9036 11744
rect 8628 11704 8634 11716
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 11514 11704 11520 11756
rect 11572 11704 11578 11756
rect 11791 11747 11849 11753
rect 11791 11713 11803 11747
rect 11837 11744 11849 11747
rect 12802 11744 12808 11756
rect 11837 11716 12808 11744
rect 11837 11713 11849 11716
rect 11791 11707 11849 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13170 11744 13176 11756
rect 13131 11716 13176 11744
rect 13170 11704 13176 11716
rect 13228 11704 13234 11756
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 15194 11744 15200 11756
rect 15155 11716 15200 11744
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 16298 11744 16304 11756
rect 15344 11716 16304 11744
rect 15344 11704 15350 11716
rect 16298 11704 16304 11716
rect 16356 11744 16362 11756
rect 18064 11753 18092 11852
rect 18616 11824 18644 11852
rect 21453 11849 21465 11883
rect 21499 11880 21511 11883
rect 22738 11880 22744 11892
rect 21499 11852 22744 11880
rect 21499 11849 21511 11852
rect 21453 11843 21511 11849
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 22830 11840 22836 11892
rect 22888 11840 22894 11892
rect 23106 11840 23112 11892
rect 23164 11840 23170 11892
rect 18322 11783 18328 11824
rect 18307 11777 18328 11783
rect 16911 11747 16969 11753
rect 16911 11744 16923 11747
rect 16356 11716 16923 11744
rect 16356 11704 16362 11716
rect 16911 11713 16923 11716
rect 16957 11713 16969 11747
rect 16911 11707 16969 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18307 11743 18319 11777
rect 18380 11772 18386 11824
rect 18598 11772 18604 11824
rect 18656 11772 18662 11824
rect 21818 11772 21824 11824
rect 21876 11812 21882 11824
rect 22848 11812 22876 11840
rect 23124 11812 23152 11840
rect 21876 11784 21956 11812
rect 21876 11772 21882 11784
rect 18353 11746 18368 11772
rect 18353 11743 18365 11746
rect 18307 11737 18365 11743
rect 18049 11707 18107 11713
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 21542 11744 21548 11756
rect 20404 11716 21548 11744
rect 20404 11704 20410 11716
rect 21542 11704 21548 11716
rect 21600 11744 21606 11756
rect 21928 11753 21956 11784
rect 22388 11784 22876 11812
rect 22940 11784 23152 11812
rect 22388 11753 22416 11784
rect 21637 11747 21695 11753
rect 21637 11744 21649 11747
rect 21600 11716 21649 11744
rect 21600 11704 21606 11716
rect 21637 11713 21649 11716
rect 21683 11713 21695 11747
rect 21637 11707 21695 11713
rect 21913 11747 21971 11753
rect 21913 11713 21925 11747
rect 21959 11713 21971 11747
rect 21913 11707 21971 11713
rect 22373 11747 22431 11753
rect 22373 11713 22385 11747
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 22741 11747 22799 11753
rect 22741 11713 22753 11747
rect 22787 11744 22799 11747
rect 22940 11744 22968 11784
rect 22787 11716 22968 11744
rect 23293 11747 23351 11753
rect 22787 11713 22799 11716
rect 22741 11707 22799 11713
rect 23293 11713 23305 11747
rect 23339 11744 23351 11747
rect 23474 11744 23480 11756
rect 23339 11716 23480 11744
rect 23339 11713 23351 11716
rect 23293 11707 23351 11713
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 23566 11704 23572 11756
rect 23624 11704 23630 11756
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11713 24179 11747
rect 24121 11707 24179 11713
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 4488 11512 6500 11540
rect 6932 11540 6960 11639
rect 8294 11636 8300 11688
rect 8352 11636 8358 11688
rect 11054 11608 11060 11620
rect 9140 11580 11060 11608
rect 9140 11552 9168 11580
rect 11054 11568 11060 11580
rect 11112 11608 11118 11620
rect 11422 11608 11428 11620
rect 11112 11580 11428 11608
rect 11112 11568 11118 11580
rect 11422 11568 11428 11580
rect 11480 11568 11486 11620
rect 7006 11540 7012 11552
rect 6932 11512 7012 11540
rect 4488 11500 4494 11512
rect 7006 11500 7012 11512
rect 7064 11540 7070 11552
rect 8202 11540 8208 11552
rect 7064 11512 8208 11540
rect 7064 11500 7070 11512
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 9122 11500 9128 11552
rect 9180 11500 9186 11552
rect 9306 11500 9312 11552
rect 9364 11500 9370 11552
rect 11532 11540 11560 11704
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 11882 11540 11888 11552
rect 11532 11512 11888 11540
rect 11882 11500 11888 11512
rect 11940 11540 11946 11552
rect 12912 11540 12940 11639
rect 13722 11636 13728 11688
rect 13780 11636 13786 11688
rect 15746 11676 15752 11688
rect 15580 11648 15752 11676
rect 11940 11512 12940 11540
rect 11940 11500 11946 11512
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13740 11540 13768 11636
rect 13044 11512 13768 11540
rect 13044 11500 13050 11512
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 15580 11540 15608 11648
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 16114 11676 16120 11688
rect 15896 11648 16120 11676
rect 15896 11636 15902 11648
rect 16114 11636 16120 11648
rect 16172 11676 16178 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16172 11648 16681 11676
rect 16172 11636 16178 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 13964 11512 15608 11540
rect 16684 11540 16712 11639
rect 22922 11636 22928 11688
rect 22980 11676 22986 11688
rect 23676 11676 23704 11707
rect 22980 11648 23704 11676
rect 22980 11636 22986 11648
rect 19150 11568 19156 11620
rect 19208 11608 19214 11620
rect 22649 11611 22707 11617
rect 22649 11608 22661 11611
rect 19208 11580 22661 11608
rect 19208 11568 19214 11580
rect 22649 11577 22661 11580
rect 22695 11577 22707 11611
rect 22649 11571 22707 11577
rect 23109 11611 23167 11617
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 24136 11608 24164 11707
rect 25038 11704 25044 11756
rect 25096 11744 25102 11756
rect 25314 11744 25320 11756
rect 25096 11716 25320 11744
rect 25096 11704 25102 11716
rect 25314 11704 25320 11716
rect 25372 11704 25378 11756
rect 23155 11580 24164 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 16942 11540 16948 11552
rect 16684 11512 16948 11540
rect 13964 11500 13970 11512
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 19058 11500 19064 11552
rect 19116 11500 19122 11552
rect 22554 11500 22560 11552
rect 22612 11540 22618 11552
rect 23385 11543 23443 11549
rect 23385 11540 23397 11543
rect 22612 11512 23397 11540
rect 22612 11500 22618 11512
rect 23385 11509 23397 11512
rect 23431 11509 23443 11543
rect 23385 11503 23443 11509
rect 23842 11500 23848 11552
rect 23900 11500 23906 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 25222 11540 25228 11552
rect 24443 11512 25228 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 1104 11450 24840 11472
rect 1104 11398 3917 11450
rect 3969 11398 3981 11450
rect 4033 11398 4045 11450
rect 4097 11398 4109 11450
rect 4161 11398 4173 11450
rect 4225 11398 9851 11450
rect 9903 11398 9915 11450
rect 9967 11398 9979 11450
rect 10031 11398 10043 11450
rect 10095 11398 10107 11450
rect 10159 11398 15785 11450
rect 15837 11398 15849 11450
rect 15901 11398 15913 11450
rect 15965 11398 15977 11450
rect 16029 11398 16041 11450
rect 16093 11398 21719 11450
rect 21771 11398 21783 11450
rect 21835 11398 21847 11450
rect 21899 11398 21911 11450
rect 21963 11398 21975 11450
rect 22027 11398 24840 11450
rect 1104 11376 24840 11398
rect 2130 11296 2136 11348
rect 2188 11296 2194 11348
rect 3050 11296 3056 11348
rect 3108 11336 3114 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3108 11308 3433 11336
rect 3108 11296 3114 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 3936 11308 4537 11336
rect 3936 11296 3942 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 5077 11339 5135 11345
rect 5077 11305 5089 11339
rect 5123 11305 5135 11339
rect 5077 11299 5135 11305
rect 1670 11228 1676 11280
rect 1728 11228 1734 11280
rect 1854 11228 1860 11280
rect 1912 11268 1918 11280
rect 2593 11271 2651 11277
rect 2593 11268 2605 11271
rect 1912 11240 2605 11268
rect 1912 11228 1918 11240
rect 2593 11237 2605 11240
rect 2639 11237 2651 11271
rect 2593 11231 2651 11237
rect 3234 11228 3240 11280
rect 3292 11268 3298 11280
rect 5092 11268 5120 11299
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7524 11308 7665 11336
rect 7524 11296 7530 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9364 11308 9628 11336
rect 9364 11296 9370 11308
rect 3292 11240 5120 11268
rect 5445 11271 5503 11277
rect 3292 11228 3298 11240
rect 5445 11237 5457 11271
rect 5491 11237 5503 11271
rect 6748 11268 6776 11296
rect 9600 11277 9628 11308
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 9858 11336 9864 11348
rect 9732 11308 9864 11336
rect 9732 11296 9738 11308
rect 9858 11296 9864 11308
rect 9916 11296 9922 11348
rect 11054 11296 11060 11348
rect 11112 11296 11118 11348
rect 11517 11339 11575 11345
rect 11517 11305 11529 11339
rect 11563 11336 11575 11339
rect 13814 11336 13820 11348
rect 11563 11308 13820 11336
rect 11563 11305 11575 11308
rect 11517 11299 11575 11305
rect 5445 11231 5503 11237
rect 5644 11240 6776 11268
rect 9585 11271 9643 11277
rect 3786 11200 3792 11212
rect 2792 11172 3792 11200
rect 1489 11135 1547 11141
rect 1489 11101 1501 11135
rect 1535 11132 1547 11135
rect 2498 11132 2504 11144
rect 1535 11104 2504 11132
rect 1535 11101 1547 11104
rect 1489 11095 1547 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 2792 11141 2820 11172
rect 3786 11160 3792 11172
rect 3844 11160 3850 11212
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4522 11200 4528 11212
rect 4028 11172 4528 11200
rect 4028 11160 4034 11172
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11101 2835 11135
rect 2777 11095 2835 11101
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 3384 11104 3617 11132
rect 3384 11092 3390 11104
rect 3605 11101 3617 11104
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 3881 11135 3939 11141
rect 3881 11101 3893 11135
rect 3927 11132 3939 11135
rect 4338 11132 4344 11144
rect 3927 11104 4344 11132
rect 3927 11101 3939 11104
rect 3881 11095 3939 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 5460 11132 5488 11231
rect 5644 11141 5672 11240
rect 9585 11237 9597 11271
rect 9631 11237 9643 11271
rect 9585 11231 9643 11237
rect 7742 11160 7748 11212
rect 7800 11160 7806 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 11532 11200 11560 11299
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 15378 11296 15384 11348
rect 15436 11296 15442 11348
rect 16758 11336 16764 11348
rect 15948 11308 16764 11336
rect 15396 11268 15424 11296
rect 15841 11271 15899 11277
rect 15841 11268 15853 11271
rect 15396 11240 15853 11268
rect 15841 11237 15853 11240
rect 15887 11237 15899 11271
rect 15841 11231 15899 11237
rect 8987 11172 11560 11200
rect 15381 11203 15439 11209
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 15381 11169 15393 11203
rect 15427 11200 15439 11203
rect 15948 11200 15976 11308
rect 16758 11296 16764 11308
rect 16816 11296 16822 11348
rect 18141 11339 18199 11345
rect 18141 11336 18153 11339
rect 17144 11308 18153 11336
rect 17034 11228 17040 11280
rect 17092 11228 17098 11280
rect 15427 11172 15976 11200
rect 15427 11169 15439 11172
rect 15381 11163 15439 11169
rect 16206 11160 16212 11212
rect 16264 11209 16270 11212
rect 16264 11203 16292 11209
rect 16280 11169 16292 11203
rect 16264 11163 16292 11169
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 17144 11200 17172 11308
rect 18141 11305 18153 11308
rect 18187 11305 18199 11339
rect 18141 11299 18199 11305
rect 18230 11296 18236 11348
rect 18288 11336 18294 11348
rect 18598 11336 18604 11348
rect 18288 11308 18604 11336
rect 18288 11296 18294 11308
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 19058 11296 19064 11348
rect 19116 11296 19122 11348
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 23753 11339 23811 11345
rect 23753 11336 23765 11339
rect 23532 11308 23765 11336
rect 23532 11296 23538 11308
rect 23753 11305 23765 11308
rect 23799 11305 23811 11339
rect 23753 11299 23811 11305
rect 17862 11228 17868 11280
rect 17920 11268 17926 11280
rect 18693 11271 18751 11277
rect 18693 11268 18705 11271
rect 17920 11240 18705 11268
rect 17920 11228 17926 11240
rect 18693 11237 18705 11240
rect 18739 11237 18751 11271
rect 18693 11231 18751 11237
rect 16439 11172 17172 11200
rect 18877 11203 18935 11209
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19076 11200 19104 11296
rect 20714 11228 20720 11280
rect 20772 11228 20778 11280
rect 22278 11228 22284 11280
rect 22336 11268 22342 11280
rect 22336 11240 22784 11268
rect 22336 11228 22342 11240
rect 22756 11212 22784 11240
rect 18923 11172 19104 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 16264 11160 16270 11163
rect 5031 11104 5488 11132
rect 5629 11135 5687 11141
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6915 11135 6973 11141
rect 6915 11101 6927 11135
rect 6961 11132 6973 11135
rect 7374 11132 7380 11144
rect 6961 11104 7380 11132
rect 6961 11101 6973 11104
rect 6915 11095 6973 11101
rect 2038 11024 2044 11076
rect 2096 11024 2102 11076
rect 2590 11024 2596 11076
rect 2648 11064 2654 11076
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2648 11036 2973 11064
rect 2648 11024 2654 11036
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 2961 11027 3019 11033
rect 3436 11036 4090 11064
rect 934 10956 940 11008
rect 992 10996 998 11008
rect 3053 10999 3111 11005
rect 3053 10996 3065 10999
rect 992 10968 3065 10996
rect 992 10956 998 10968
rect 3053 10965 3065 10968
rect 3099 10965 3111 10999
rect 3053 10959 3111 10965
rect 3326 10956 3332 11008
rect 3384 10996 3390 11008
rect 3436 10996 3464 11036
rect 3384 10968 3464 10996
rect 3384 10956 3390 10968
rect 3970 10956 3976 11008
rect 4028 10956 4034 11008
rect 4062 10996 4090 11036
rect 4430 11024 4436 11076
rect 4488 11024 4494 11076
rect 6656 11064 6684 11095
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7760 11132 7788 11160
rect 7484 11104 7788 11132
rect 7006 11064 7012 11076
rect 6656 11036 7012 11064
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7484 10996 7512 11104
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 7984 11104 8493 11132
rect 7984 11092 7990 11104
rect 8481 11101 8493 11104
rect 8527 11132 8539 11135
rect 9122 11132 9128 11144
rect 8527 11104 9128 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 9950 11092 9956 11144
rect 10008 11141 10014 11144
rect 10008 11135 10036 11141
rect 10024 11101 10036 11135
rect 10008 11095 10036 11101
rect 10008 11092 10014 11095
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 12710 11092 12716 11144
rect 12768 11132 12774 11144
rect 13170 11132 13176 11144
rect 12768 11104 13176 11132
rect 12768 11092 12774 11104
rect 13170 11092 13176 11104
rect 13228 11092 13234 11144
rect 15197 11135 15255 11141
rect 15197 11101 15209 11135
rect 15243 11101 15255 11135
rect 15197 11095 15255 11101
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 7800 11036 9168 11064
rect 7800 11024 7806 11036
rect 4062 10968 7512 10996
rect 9140 10996 9168 11036
rect 10612 11036 10793 11064
rect 10612 10996 10640 11036
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 15212 11064 15240 11095
rect 16114 11092 16120 11144
rect 16172 11092 16178 11144
rect 17129 11135 17187 11141
rect 17129 11132 17141 11135
rect 16960 11104 17141 11132
rect 16960 11076 16988 11104
rect 17129 11101 17141 11104
rect 17175 11101 17187 11135
rect 17402 11132 17408 11144
rect 17363 11104 17408 11132
rect 17129 11095 17187 11101
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 18656 11104 18705 11132
rect 18656 11092 18662 11104
rect 18693 11101 18705 11104
rect 18739 11101 18751 11135
rect 19076 11132 19104 11172
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 22370 11200 22376 11212
rect 19576 11172 22376 11200
rect 19576 11160 19582 11172
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 22738 11160 22744 11212
rect 22796 11160 22802 11212
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 19076 11104 19257 11132
rect 18693 11095 18751 11101
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 20254 11092 20260 11144
rect 20312 11092 20318 11144
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 21174 11092 21180 11144
rect 21232 11132 21238 11144
rect 22922 11132 22928 11144
rect 21232 11104 22928 11132
rect 21232 11092 21238 11104
rect 22922 11092 22928 11104
rect 22980 11141 22986 11144
rect 22980 11135 23041 11141
rect 22980 11101 22995 11135
rect 23029 11101 23041 11135
rect 22980 11095 23041 11101
rect 22980 11092 22986 11095
rect 15378 11064 15384 11076
rect 15212 11036 15384 11064
rect 10781 11027 10839 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 16942 11024 16948 11076
rect 17000 11064 17006 11076
rect 17218 11064 17224 11076
rect 17000 11036 17224 11064
rect 17000 11024 17006 11036
rect 17218 11024 17224 11036
rect 17276 11024 17282 11076
rect 17420 11064 17448 11092
rect 17586 11064 17592 11076
rect 17420 11036 17592 11064
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 19061 11067 19119 11073
rect 19061 11033 19073 11067
rect 19107 11064 19119 11067
rect 19337 11067 19395 11073
rect 19337 11064 19349 11067
rect 19107 11036 19349 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 19337 11033 19349 11036
rect 19383 11033 19395 11067
rect 19794 11064 19800 11076
rect 19337 11027 19395 11033
rect 19444 11036 19800 11064
rect 9140 10968 10640 10996
rect 13170 10956 13176 11008
rect 13228 10996 13234 11008
rect 15286 10996 15292 11008
rect 13228 10968 15292 10996
rect 13228 10956 13234 10968
rect 15286 10956 15292 10968
rect 15344 10956 15350 11008
rect 16298 10956 16304 11008
rect 16356 10996 16362 11008
rect 19444 10996 19472 11036
rect 19794 11024 19800 11036
rect 19852 11024 19858 11076
rect 16356 10968 19472 10996
rect 16356 10956 16362 10968
rect 19518 10956 19524 11008
rect 19576 10996 19582 11008
rect 20622 10996 20628 11008
rect 19576 10968 20628 10996
rect 19576 10956 19582 10968
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 21450 10956 21456 11008
rect 21508 10996 21514 11008
rect 23566 10996 23572 11008
rect 21508 10968 23572 10996
rect 21508 10956 21514 10968
rect 23566 10956 23572 10968
rect 23624 10956 23630 11008
rect 1104 10906 25000 10928
rect 1104 10854 6884 10906
rect 6936 10854 6948 10906
rect 7000 10854 7012 10906
rect 7064 10854 7076 10906
rect 7128 10854 7140 10906
rect 7192 10854 12818 10906
rect 12870 10854 12882 10906
rect 12934 10854 12946 10906
rect 12998 10854 13010 10906
rect 13062 10854 13074 10906
rect 13126 10854 18752 10906
rect 18804 10854 18816 10906
rect 18868 10854 18880 10906
rect 18932 10854 18944 10906
rect 18996 10854 19008 10906
rect 19060 10854 24686 10906
rect 24738 10854 24750 10906
rect 24802 10854 24814 10906
rect 24866 10854 24878 10906
rect 24930 10854 24942 10906
rect 24994 10854 25000 10906
rect 1104 10832 25000 10854
rect 1578 10752 1584 10804
rect 1636 10752 1642 10804
rect 2038 10752 2044 10804
rect 2096 10792 2102 10804
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 2096 10764 3801 10792
rect 2096 10752 2102 10764
rect 3789 10761 3801 10764
rect 3835 10761 3847 10795
rect 4338 10792 4344 10804
rect 3789 10755 3847 10761
rect 3896 10764 4344 10792
rect 1486 10684 1492 10736
rect 1544 10684 1550 10736
rect 3896 10724 3924 10764
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 5626 10792 5632 10804
rect 4580 10764 5632 10792
rect 4580 10752 4586 10764
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 6454 10792 6460 10804
rect 5868 10764 6460 10792
rect 5868 10752 5874 10764
rect 6454 10752 6460 10764
rect 6512 10752 6518 10804
rect 7466 10752 7472 10804
rect 7524 10792 7530 10804
rect 8662 10792 8668 10804
rect 7524 10764 8668 10792
rect 7524 10752 7530 10764
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 9766 10752 9772 10804
rect 9824 10752 9830 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 10192 10764 10241 10792
rect 10192 10752 10198 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 10229 10755 10287 10761
rect 10318 10764 10977 10792
rect 7558 10724 7564 10736
rect 2514 10696 3924 10724
rect 3988 10696 7564 10724
rect 2514 10695 2542 10696
rect 2483 10689 2542 10695
rect 2130 10616 2136 10668
rect 2188 10616 2194 10668
rect 2483 10655 2495 10689
rect 2529 10658 2542 10689
rect 3988 10665 4016 10696
rect 7558 10684 7564 10696
rect 7616 10684 7622 10736
rect 9784 10724 9812 10752
rect 10318 10724 10346 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 11790 10752 11796 10804
rect 11848 10792 11854 10804
rect 12250 10792 12256 10804
rect 11848 10764 12256 10792
rect 11848 10752 11854 10764
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 13262 10752 13268 10804
rect 13320 10752 13326 10804
rect 14274 10792 14280 10804
rect 13648 10764 14280 10792
rect 9784 10696 10346 10724
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 13170 10724 13176 10736
rect 10928 10696 13176 10724
rect 10928 10684 10934 10696
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 3973 10659 4031 10665
rect 2529 10655 2541 10658
rect 2483 10649 2541 10655
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 4338 10656 4344 10668
rect 4299 10628 4344 10656
rect 3973 10619 4031 10625
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6178 10656 6184 10668
rect 5868 10628 6184 10656
rect 5868 10616 5874 10628
rect 6178 10616 6184 10628
rect 6236 10656 6242 10668
rect 6607 10659 6665 10665
rect 6607 10656 6619 10659
rect 6236 10628 6619 10656
rect 6236 10616 6242 10628
rect 6607 10625 6619 10628
rect 6653 10625 6665 10659
rect 6607 10619 6665 10625
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 9398 10656 9404 10668
rect 8628 10628 9404 10656
rect 8628 10616 8634 10628
rect 9398 10616 9404 10628
rect 9456 10665 9462 10668
rect 9456 10659 9517 10665
rect 9456 10625 9471 10659
rect 9505 10625 9517 10659
rect 9456 10619 9517 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 11238 10656 11244 10668
rect 10827 10628 11244 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 9456 10616 9462 10619
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 12343 10659 12401 10665
rect 12343 10656 12355 10659
rect 11348 10628 12355 10656
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1762 10588 1768 10600
rect 1360 10560 1768 10588
rect 1360 10548 1366 10560
rect 1762 10548 1768 10560
rect 1820 10588 1826 10600
rect 2225 10591 2283 10597
rect 2225 10588 2237 10591
rect 1820 10560 2237 10588
rect 1820 10548 1826 10560
rect 2225 10557 2237 10560
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 4062 10548 4068 10600
rect 4120 10548 4126 10600
rect 4982 10548 4988 10600
rect 5040 10588 5046 10600
rect 5166 10588 5172 10600
rect 5040 10560 5172 10588
rect 5040 10548 5046 10560
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 1946 10412 1952 10464
rect 2004 10412 2010 10464
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 3016 10424 3249 10452
rect 3016 10412 3022 10424
rect 3237 10421 3249 10424
rect 3283 10421 3295 10455
rect 3237 10415 3295 10421
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 5077 10455 5135 10461
rect 5077 10452 5089 10455
rect 5040 10424 5089 10452
rect 5040 10412 5046 10424
rect 5077 10421 5089 10424
rect 5123 10421 5135 10455
rect 6380 10452 6408 10551
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 9214 10588 9220 10600
rect 8352 10560 9220 10588
rect 8352 10548 8358 10560
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 6822 10452 6828 10464
rect 6380 10424 6828 10452
rect 5077 10415 5135 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7374 10412 7380 10464
rect 7432 10412 7438 10464
rect 8018 10412 8024 10464
rect 8076 10452 8082 10464
rect 11348 10452 11376 10628
rect 12343 10625 12355 10628
rect 12389 10656 12401 10659
rect 13280 10656 13308 10752
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 13648 10733 13676 10764
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 16206 10792 16212 10804
rect 14967 10764 16212 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 17696 10764 19923 10792
rect 13633 10727 13691 10733
rect 13633 10724 13645 10727
rect 13504 10696 13645 10724
rect 13504 10684 13510 10696
rect 13633 10693 13645 10696
rect 13679 10693 13691 10727
rect 13633 10687 13691 10693
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 14182 10724 14188 10736
rect 13964 10696 14188 10724
rect 13964 10684 13970 10696
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 14369 10727 14427 10733
rect 14369 10693 14381 10727
rect 14415 10724 14427 10727
rect 14642 10724 14648 10736
rect 14415 10696 14648 10724
rect 14415 10693 14427 10696
rect 14369 10687 14427 10693
rect 14642 10684 14648 10696
rect 14700 10684 14706 10736
rect 14734 10684 14740 10736
rect 14792 10724 14798 10736
rect 15102 10724 15108 10736
rect 14792 10696 15108 10724
rect 14792 10684 14798 10696
rect 15102 10684 15108 10696
rect 15160 10684 15166 10736
rect 12389 10628 13308 10656
rect 12389 10625 12401 10628
rect 12343 10619 12401 10625
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 17696 10665 17724 10764
rect 17788 10696 19656 10724
rect 17788 10665 17816 10696
rect 19628 10668 19656 10696
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17773 10659 17831 10665
rect 17773 10625 17785 10659
rect 17819 10625 17831 10659
rect 18029 10659 18087 10665
rect 18029 10656 18041 10659
rect 17773 10619 17831 10625
rect 17880 10628 18041 10656
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 11882 10588 11888 10600
rect 11480 10560 11888 10588
rect 11480 10548 11486 10560
rect 11882 10548 11888 10560
rect 11940 10588 11946 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11940 10560 12081 10588
rect 11940 10548 11946 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 17696 10588 17724 10619
rect 17880 10588 17908 10628
rect 18029 10625 18041 10628
rect 18075 10625 18087 10659
rect 18029 10619 18087 10625
rect 18322 10616 18328 10668
rect 18380 10656 18386 10668
rect 19518 10656 19524 10668
rect 18380 10628 19288 10656
rect 19479 10628 19524 10656
rect 18380 10616 18386 10628
rect 19260 10597 19288 10628
rect 19518 10616 19524 10628
rect 19576 10616 19582 10668
rect 19610 10616 19616 10668
rect 19668 10616 19674 10668
rect 12069 10551 12127 10557
rect 13081 10523 13139 10529
rect 13081 10489 13093 10523
rect 13127 10520 13139 10523
rect 13464 10520 13492 10574
rect 17696 10560 17908 10588
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19895 10588 19923 10764
rect 20070 10752 20076 10804
rect 20128 10792 20134 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 20128 10764 20269 10792
rect 20128 10752 20134 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20257 10755 20315 10761
rect 20272 10656 20300 10755
rect 20714 10752 20720 10804
rect 20772 10752 20778 10804
rect 20990 10752 20996 10804
rect 21048 10752 21054 10804
rect 21008 10724 21036 10752
rect 23198 10724 23204 10736
rect 20732 10696 21036 10724
rect 22998 10696 23204 10724
rect 20732 10668 20760 10696
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 20272 10628 20637 10656
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20714 10616 20720 10668
rect 20772 10616 20778 10668
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 20855 10628 20944 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 19895 10560 20852 10588
rect 19245 10551 19303 10557
rect 13127 10492 13492 10520
rect 13127 10489 13139 10492
rect 13081 10483 13139 10489
rect 8076 10424 11376 10452
rect 8076 10412 8082 10424
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 13630 10452 13636 10464
rect 13228 10424 13636 10452
rect 13228 10412 13234 10424
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 17494 10412 17500 10464
rect 17552 10412 17558 10464
rect 19150 10412 19156 10464
rect 19208 10412 19214 10464
rect 19260 10452 19288 10551
rect 20714 10452 20720 10464
rect 19260 10424 20720 10452
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 20824 10452 20852 10560
rect 20916 10529 20944 10628
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 20901 10523 20959 10529
rect 20901 10489 20913 10523
rect 20947 10489 20959 10523
rect 20901 10483 20959 10489
rect 20990 10452 20996 10464
rect 20824 10424 20996 10452
rect 20990 10412 20996 10424
rect 21048 10412 21054 10464
rect 22465 10455 22523 10461
rect 22465 10421 22477 10455
rect 22511 10452 22523 10455
rect 22554 10452 22560 10464
rect 22511 10424 22560 10452
rect 22511 10421 22523 10424
rect 22465 10415 22523 10421
rect 22554 10412 22560 10424
rect 22612 10412 22618 10464
rect 22664 10452 22692 10619
rect 22738 10616 22744 10668
rect 22796 10616 22802 10668
rect 22998 10665 23026 10696
rect 23198 10684 23204 10696
rect 23256 10684 23262 10736
rect 22983 10659 23041 10665
rect 22983 10625 22995 10659
rect 23029 10625 23041 10659
rect 22983 10619 23041 10625
rect 23753 10455 23811 10461
rect 23753 10452 23765 10455
rect 22664 10424 23765 10452
rect 23753 10421 23765 10424
rect 23799 10421 23811 10455
rect 23753 10415 23811 10421
rect 1104 10362 24840 10384
rect 1104 10310 3917 10362
rect 3969 10310 3981 10362
rect 4033 10310 4045 10362
rect 4097 10310 4109 10362
rect 4161 10310 4173 10362
rect 4225 10310 9851 10362
rect 9903 10310 9915 10362
rect 9967 10310 9979 10362
rect 10031 10310 10043 10362
rect 10095 10310 10107 10362
rect 10159 10310 15785 10362
rect 15837 10310 15849 10362
rect 15901 10310 15913 10362
rect 15965 10310 15977 10362
rect 16029 10310 16041 10362
rect 16093 10310 21719 10362
rect 21771 10310 21783 10362
rect 21835 10310 21847 10362
rect 21899 10310 21911 10362
rect 21963 10310 21975 10362
rect 22027 10310 24840 10362
rect 1104 10288 24840 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 2188 10220 3617 10248
rect 2188 10208 2194 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 5994 10248 6000 10260
rect 4120 10220 6000 10248
rect 4120 10208 4126 10220
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 7282 10248 7288 10260
rect 6420 10220 7288 10248
rect 6420 10208 6426 10220
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 7374 10208 7380 10260
rect 7432 10208 7438 10260
rect 7558 10208 7564 10260
rect 7616 10208 7622 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 14056 10220 15117 10248
rect 14056 10208 14062 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 17494 10208 17500 10260
rect 17552 10208 17558 10260
rect 18417 10251 18475 10257
rect 18417 10217 18429 10251
rect 18463 10248 18475 10251
rect 18598 10248 18604 10260
rect 18463 10220 18604 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 19150 10208 19156 10260
rect 19208 10208 19214 10260
rect 20165 10251 20223 10257
rect 20165 10217 20177 10251
rect 20211 10248 20223 10251
rect 20254 10248 20260 10260
rect 20211 10220 20260 10248
rect 20211 10217 20223 10220
rect 20165 10211 20223 10217
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20714 10208 20720 10260
rect 20772 10248 20778 10260
rect 20772 10220 20852 10248
rect 20772 10208 20778 10220
rect 3896 10152 4568 10180
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2130 10112 2136 10124
rect 1995 10084 2136 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 2406 10072 2412 10124
rect 2464 10072 2470 10124
rect 2682 10072 2688 10124
rect 2740 10112 2746 10124
rect 3896 10112 3924 10152
rect 2740 10084 3924 10112
rect 2740 10072 2746 10084
rect 3970 10072 3976 10124
rect 4028 10072 4034 10124
rect 4430 10072 4436 10124
rect 4488 10072 4494 10124
rect 4540 10112 4568 10152
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 6236 10152 6500 10180
rect 6236 10140 6242 10152
rect 6472 10124 6500 10152
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4540 10084 4721 10112
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 4798 10072 4804 10124
rect 4856 10121 4862 10124
rect 4856 10115 4884 10121
rect 4872 10081 4884 10115
rect 4856 10075 4884 10081
rect 4856 10072 4862 10075
rect 4982 10072 4988 10124
rect 5040 10072 5046 10124
rect 5166 10072 5172 10124
rect 5224 10112 5230 10124
rect 5224 10084 5764 10112
rect 5224 10072 5230 10084
rect 474 10004 480 10056
rect 532 10044 538 10056
rect 2866 10053 2872 10056
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 532 10016 1777 10044
rect 532 10004 538 10016
rect 1765 10013 1777 10016
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 2823 10047 2872 10053
rect 2823 10013 2835 10047
rect 2869 10013 2872 10047
rect 2823 10007 2872 10013
rect 2866 10004 2872 10007
rect 2924 10004 2930 10056
rect 2958 10004 2964 10056
rect 3016 10004 3022 10056
rect 3602 10004 3608 10056
rect 3660 10044 3666 10056
rect 5736 10053 5764 10084
rect 6086 10072 6092 10124
rect 6144 10072 6150 10124
rect 6362 10072 6368 10124
rect 6420 10072 6426 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6512 10084 6653 10112
rect 6512 10072 6518 10084
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 6730 10072 6736 10124
rect 6788 10121 6794 10124
rect 6788 10115 6816 10121
rect 6804 10081 6816 10115
rect 6788 10075 6816 10081
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7392 10112 7420 10208
rect 10965 10183 11023 10189
rect 10965 10149 10977 10183
rect 11011 10149 11023 10183
rect 10965 10143 11023 10149
rect 10870 10112 10876 10124
rect 6963 10084 7420 10112
rect 10612 10084 10876 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 6788 10072 6794 10075
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3660 10016 3801 10044
rect 3660 10004 3666 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10044 5963 10047
rect 6104 10044 6132 10072
rect 5951 10016 6132 10044
rect 9953 10047 10011 10053
rect 5951 10013 5963 10016
rect 5905 10007 5963 10013
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10227 10047 10285 10053
rect 10227 10013 10239 10047
rect 10273 10044 10285 10047
rect 10612 10044 10640 10084
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10980 10112 11008 10143
rect 10980 10084 11362 10112
rect 10273 10016 10640 10044
rect 10273 10013 10285 10016
rect 10227 10007 10285 10013
rect 9968 9976 9996 10007
rect 10686 10004 10692 10056
rect 10744 10044 10750 10056
rect 11885 10047 11943 10053
rect 10744 10016 11744 10044
rect 10744 10004 10750 10016
rect 11422 9976 11428 9988
rect 5460 9948 5762 9976
rect 9968 9948 11428 9976
rect 4890 9868 4896 9920
rect 4948 9908 4954 9920
rect 5460 9908 5488 9948
rect 4948 9880 5488 9908
rect 4948 9868 4954 9880
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 5734 9908 5762 9948
rect 11422 9936 11428 9948
rect 11480 9936 11486 9988
rect 6822 9908 6828 9920
rect 5734 9880 6828 9908
rect 6822 9868 6828 9880
rect 6880 9908 6886 9920
rect 9030 9908 9036 9920
rect 6880 9880 9036 9908
rect 6880 9868 6886 9880
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10686 9908 10692 9920
rect 10560 9880 10692 9908
rect 10560 9868 10566 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 11606 9908 11612 9920
rect 11563 9880 11612 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 11716 9908 11744 10016
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12618 10044 12624 10056
rect 11931 10016 12624 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 14056 10016 14105 10044
rect 14056 10004 14062 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 17512 10044 17540 10208
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 14093 10007 14151 10013
rect 14351 10017 14409 10023
rect 11793 9979 11851 9985
rect 11793 9945 11805 9979
rect 11839 9976 11851 9979
rect 11974 9976 11980 9988
rect 11839 9948 11980 9976
rect 11839 9945 11851 9948
rect 11793 9939 11851 9945
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 12158 9936 12164 9988
rect 12216 9976 12222 9988
rect 12253 9979 12311 9985
rect 12253 9976 12265 9979
rect 12216 9948 12265 9976
rect 12216 9936 12222 9948
rect 12253 9945 12265 9948
rect 12299 9945 12311 9979
rect 14351 9983 14363 10017
rect 14397 10014 14409 10017
rect 17512 10016 18337 10044
rect 14397 9988 14412 10014
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10044 19119 10047
rect 19168 10044 19196 10208
rect 20349 10183 20407 10189
rect 20349 10149 20361 10183
rect 20395 10149 20407 10183
rect 20349 10143 20407 10149
rect 19107 10016 19196 10044
rect 19260 10084 19564 10112
rect 19107 10013 19119 10016
rect 19061 10007 19119 10013
rect 14351 9977 14372 9983
rect 12253 9939 12311 9945
rect 12406 9948 12848 9976
rect 12406 9908 12434 9948
rect 11716 9880 12434 9908
rect 12526 9868 12532 9920
rect 12584 9908 12590 9920
rect 12820 9917 12848 9948
rect 14366 9936 14372 9977
rect 14424 9976 14430 9988
rect 19260 9976 19288 10084
rect 19426 10004 19432 10056
rect 19484 10004 19490 10056
rect 14424 9948 19288 9976
rect 14424 9936 14430 9948
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12584 9880 12633 9908
rect 12584 9868 12590 9880
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 12621 9871 12679 9877
rect 12805 9911 12863 9917
rect 12805 9877 12817 9911
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 18877 9911 18935 9917
rect 18877 9877 18889 9911
rect 18923 9908 18935 9911
rect 19444 9908 19472 10004
rect 19536 9976 19564 10084
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10044 20131 10047
rect 20364 10044 20392 10143
rect 20438 10140 20444 10192
rect 20496 10180 20502 10192
rect 20496 10152 20760 10180
rect 20496 10140 20502 10152
rect 20119 10016 20392 10044
rect 20456 10084 20668 10112
rect 20119 10013 20131 10016
rect 20073 10007 20131 10013
rect 20456 9976 20484 10084
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 19536 9948 20484 9976
rect 20548 9920 20576 10007
rect 20640 9976 20668 10084
rect 20732 10044 20760 10152
rect 20824 10121 20852 10220
rect 22462 10208 22468 10260
rect 22520 10248 22526 10260
rect 22520 10220 23428 10248
rect 22520 10208 22526 10220
rect 22094 10140 22100 10192
rect 22152 10180 22158 10192
rect 22738 10180 22744 10192
rect 22152 10152 22744 10180
rect 22152 10140 22158 10152
rect 22738 10140 22744 10152
rect 22796 10140 22802 10192
rect 20809 10115 20867 10121
rect 20809 10081 20821 10115
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 22278 10072 22284 10124
rect 22336 10112 22342 10124
rect 22336 10084 22784 10112
rect 22336 10072 22342 10084
rect 21051 10047 21109 10053
rect 21051 10044 21063 10047
rect 20732 10016 21063 10044
rect 21051 10013 21063 10016
rect 21097 10013 21109 10047
rect 21051 10007 21109 10013
rect 22462 10004 22468 10056
rect 22520 10004 22526 10056
rect 22756 10053 22784 10084
rect 22741 10047 22799 10053
rect 22741 10013 22753 10047
rect 22787 10013 22799 10047
rect 22741 10007 22799 10013
rect 22983 10047 23041 10053
rect 22983 10013 22995 10047
rect 23029 10044 23041 10047
rect 23400 10044 23428 10220
rect 24578 10140 24584 10192
rect 24636 10180 24642 10192
rect 25130 10180 25136 10192
rect 24636 10152 25136 10180
rect 24636 10140 24642 10152
rect 25130 10140 25136 10152
rect 25188 10140 25194 10192
rect 23029 10016 23428 10044
rect 23029 10013 23041 10016
rect 22983 10007 23041 10013
rect 22756 9976 22784 10007
rect 20640 9948 22416 9976
rect 22756 9948 23060 9976
rect 18923 9880 19472 9908
rect 18923 9877 18935 9880
rect 18877 9871 18935 9877
rect 20530 9868 20536 9920
rect 20588 9868 20594 9920
rect 21821 9911 21879 9917
rect 21821 9877 21833 9911
rect 21867 9908 21879 9911
rect 22186 9908 22192 9920
rect 21867 9880 22192 9908
rect 21867 9877 21879 9880
rect 21821 9871 21879 9877
rect 22186 9868 22192 9880
rect 22244 9868 22250 9920
rect 22278 9868 22284 9920
rect 22336 9868 22342 9920
rect 22388 9908 22416 9948
rect 23032 9920 23060 9948
rect 22738 9908 22744 9920
rect 22388 9880 22744 9908
rect 22738 9868 22744 9880
rect 22796 9868 22802 9920
rect 23014 9868 23020 9920
rect 23072 9868 23078 9920
rect 23750 9868 23756 9920
rect 23808 9868 23814 9920
rect 1104 9818 25000 9840
rect 1104 9766 6884 9818
rect 6936 9766 6948 9818
rect 7000 9766 7012 9818
rect 7064 9766 7076 9818
rect 7128 9766 7140 9818
rect 7192 9766 12818 9818
rect 12870 9766 12882 9818
rect 12934 9766 12946 9818
rect 12998 9766 13010 9818
rect 13062 9766 13074 9818
rect 13126 9766 18752 9818
rect 18804 9766 18816 9818
rect 18868 9766 18880 9818
rect 18932 9766 18944 9818
rect 18996 9766 19008 9818
rect 19060 9766 24686 9818
rect 24738 9766 24750 9818
rect 24802 9766 24814 9818
rect 24866 9766 24878 9818
rect 24930 9766 24942 9818
rect 24994 9766 25000 9818
rect 1104 9744 25000 9766
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 2685 9707 2743 9713
rect 2685 9704 2697 9707
rect 2464 9676 2697 9704
rect 2464 9664 2470 9676
rect 2685 9673 2697 9676
rect 2731 9673 2743 9707
rect 4154 9704 4160 9716
rect 2685 9667 2743 9673
rect 3160 9676 4160 9704
rect 3160 9648 3188 9676
rect 4154 9664 4160 9676
rect 4212 9664 4218 9716
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 4525 9707 4583 9713
rect 4525 9704 4537 9707
rect 4488 9676 4537 9704
rect 4488 9664 4494 9676
rect 4525 9673 4537 9676
rect 4571 9673 4583 9707
rect 4525 9667 4583 9673
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6362 9704 6368 9716
rect 5951 9676 6368 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 7834 9704 7840 9716
rect 7432 9676 7840 9704
rect 7432 9664 7438 9676
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 10134 9664 10140 9716
rect 10192 9704 10198 9716
rect 10594 9704 10600 9716
rect 10192 9676 10600 9704
rect 10192 9664 10198 9676
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 10870 9704 10876 9716
rect 10744 9676 10876 9704
rect 10744 9664 10750 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11238 9664 11244 9716
rect 11296 9664 11302 9716
rect 11992 9676 12204 9704
rect 14 9596 20 9648
rect 72 9636 78 9648
rect 72 9608 1716 9636
rect 72 9596 78 9608
rect 1302 9528 1308 9580
rect 1360 9528 1366 9580
rect 1578 9528 1584 9580
rect 1636 9528 1642 9580
rect 1688 9568 1716 9608
rect 3142 9596 3148 9648
rect 3200 9596 3206 9648
rect 3510 9636 3516 9648
rect 3252 9608 3516 9636
rect 3252 9577 3280 9608
rect 3510 9596 3516 9608
rect 3568 9596 3574 9648
rect 11992 9636 12020 9676
rect 11164 9608 12020 9636
rect 1915 9571 1973 9577
rect 1915 9568 1927 9571
rect 1688 9540 1927 9568
rect 1915 9537 1927 9540
rect 1961 9568 1973 9571
rect 3237 9571 3295 9577
rect 1961 9540 2774 9568
rect 1961 9537 1973 9540
rect 1915 9531 1973 9537
rect 1320 9500 1348 9528
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1320 9472 1685 9500
rect 1596 9444 1624 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 2746 9500 2774 9540
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3755 9571 3813 9577
rect 3755 9568 3767 9571
rect 3237 9531 3295 9537
rect 3344 9540 3767 9568
rect 3344 9500 3372 9540
rect 3755 9537 3767 9540
rect 3801 9537 3813 9571
rect 3755 9531 3813 9537
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 5135 9571 5193 9577
rect 5135 9568 5147 9571
rect 4764 9540 5147 9568
rect 4764 9528 4770 9540
rect 5135 9537 5147 9540
rect 5181 9537 5193 9571
rect 7653 9571 7711 9577
rect 7653 9568 7665 9571
rect 5135 9531 5193 9537
rect 6380 9540 7665 9568
rect 6380 9512 6408 9540
rect 7653 9537 7665 9540
rect 7699 9568 7711 9571
rect 7834 9568 7840 9580
rect 7699 9540 7840 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8384 9528 8390 9580
rect 8442 9568 8448 9580
rect 8651 9571 8709 9577
rect 8442 9540 8487 9568
rect 8442 9528 8448 9540
rect 8651 9537 8663 9571
rect 8697 9537 8709 9571
rect 8651 9531 8709 9537
rect 3501 9503 3559 9509
rect 3501 9500 3513 9503
rect 2746 9472 3372 9500
rect 1673 9463 1731 9469
rect 3482 9469 3513 9500
rect 3547 9469 3559 9503
rect 3482 9463 3559 9469
rect 1578 9392 1584 9444
rect 1636 9392 1642 9444
rect 2774 9392 2780 9444
rect 2832 9392 2838 9444
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 3482 9432 3510 9463
rect 4890 9460 4896 9512
rect 4948 9460 4954 9512
rect 6362 9460 6368 9512
rect 6420 9460 6426 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 3200 9404 3510 9432
rect 3200 9392 3206 9404
rect 1397 9367 1455 9373
rect 1397 9333 1409 9367
rect 1443 9364 1455 9367
rect 2792 9364 2820 9392
rect 1443 9336 2820 9364
rect 1443 9333 1455 9336
rect 1397 9327 1455 9333
rect 3050 9324 3056 9376
rect 3108 9324 3114 9376
rect 7484 9364 7512 9463
rect 8478 9460 8484 9512
rect 8536 9509 8542 9512
rect 8536 9503 8585 9509
rect 8536 9469 8539 9503
rect 8573 9469 8585 9503
rect 8680 9500 8708 9531
rect 9306 9528 9312 9580
rect 9364 9528 9370 9580
rect 9398 9528 9404 9580
rect 9456 9528 9462 9580
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10502 9577 10508 9580
rect 10459 9571 10508 9577
rect 10459 9537 10471 9571
rect 10505 9537 10508 9571
rect 10459 9531 10508 9537
rect 10502 9528 10508 9531
rect 10560 9528 10566 9580
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 9582 9500 9588 9512
rect 8680 9472 9444 9500
rect 9543 9472 9588 9500
rect 8536 9463 8585 9469
rect 8536 9460 8542 9463
rect 8110 9392 8116 9444
rect 8168 9392 8174 9444
rect 9416 9432 9444 9472
rect 9582 9460 9588 9472
rect 9640 9500 9646 9512
rect 10134 9500 10140 9512
rect 9640 9472 10140 9500
rect 9640 9460 9646 9472
rect 10134 9460 10140 9472
rect 10192 9500 10198 9512
rect 11164 9500 11192 9608
rect 12176 9598 12204 9676
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12805 9707 12863 9713
rect 12805 9704 12817 9707
rect 12676 9676 12817 9704
rect 12676 9664 12682 9676
rect 12805 9673 12817 9676
rect 12851 9673 12863 9707
rect 13262 9704 13268 9716
rect 12805 9667 12863 9673
rect 13004 9676 13268 9704
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11480 9540 11805 9568
rect 11480 9528 11486 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 12066 9568 12072 9580
rect 12027 9540 12072 9568
rect 11793 9531 11851 9537
rect 10192 9472 11192 9500
rect 10192 9460 10198 9472
rect 10045 9435 10103 9441
rect 9416 9404 9628 9432
rect 9600 9376 9628 9404
rect 10045 9401 10057 9435
rect 10091 9401 10103 9435
rect 10045 9395 10103 9401
rect 9398 9364 9404 9376
rect 7484 9336 9404 9364
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9582 9324 9588 9376
rect 9640 9324 9646 9376
rect 10060 9364 10088 9395
rect 10318 9364 10324 9376
rect 10060 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 11808 9364 11836 9531
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 12176 9570 12296 9598
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 13004 9636 13032 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 15102 9704 15108 9716
rect 14056 9676 15108 9704
rect 14056 9664 14062 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 16298 9704 16304 9716
rect 15344 9676 16304 9704
rect 15344 9664 15350 9676
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 17954 9704 17960 9716
rect 16632 9676 17960 9704
rect 16632 9664 16638 9676
rect 17954 9664 17960 9676
rect 18012 9664 18018 9716
rect 21082 9664 21088 9716
rect 21140 9664 21146 9716
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 23658 9704 23664 9716
rect 22428 9676 23664 9704
rect 22428 9664 22434 9676
rect 23658 9664 23664 9676
rect 23716 9664 23722 9716
rect 12400 9608 13032 9636
rect 12400 9596 12406 9608
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 18196 9608 18451 9636
rect 18196 9596 18202 9608
rect 12268 9568 12296 9570
rect 12268 9540 14136 9568
rect 12618 9364 12624 9376
rect 11808 9336 12624 9364
rect 12618 9324 12624 9336
rect 12676 9364 12682 9376
rect 13998 9364 14004 9376
rect 12676 9336 14004 9364
rect 12676 9324 12682 9336
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14108 9364 14136 9540
rect 18322 9528 18328 9580
rect 18380 9528 18386 9580
rect 18423 9568 18451 9608
rect 18583 9601 18641 9607
rect 18583 9568 18595 9601
rect 18423 9567 18595 9568
rect 18629 9567 18641 9601
rect 19794 9596 19800 9648
rect 19852 9636 19858 9648
rect 19852 9608 20760 9636
rect 19852 9596 19858 9608
rect 18423 9561 18641 9567
rect 19972 9571 20030 9577
rect 18423 9540 18626 9561
rect 19972 9537 19984 9571
rect 20018 9568 20030 9571
rect 20530 9568 20536 9580
rect 20018 9540 20536 9568
rect 20018 9537 20030 9540
rect 19972 9531 20030 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 19518 9500 19524 9512
rect 19392 9472 19524 9500
rect 19392 9460 19398 9472
rect 19518 9460 19524 9472
rect 19576 9460 19582 9512
rect 19610 9460 19616 9512
rect 19668 9500 19674 9512
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 19668 9472 19717 9500
rect 19668 9460 19674 9472
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 17954 9432 17960 9444
rect 15160 9404 17960 9432
rect 15160 9392 15166 9404
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 20732 9432 20760 9608
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9568 22155 9571
rect 22186 9568 22192 9580
rect 22143 9540 22192 9568
rect 22143 9537 22155 9540
rect 22097 9531 22155 9537
rect 21836 9500 21864 9531
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 22296 9577 22324 9664
rect 23842 9596 23848 9648
rect 23900 9636 23906 9648
rect 25682 9636 25688 9648
rect 23900 9608 25688 9636
rect 23900 9596 23906 9608
rect 25682 9596 25688 9608
rect 25740 9596 25746 9648
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 22370 9528 22376 9580
rect 22428 9568 22434 9580
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22428 9540 22569 9568
rect 22428 9528 22434 9540
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 22983 9571 23041 9577
rect 22983 9568 22995 9571
rect 22557 9531 22615 9537
rect 22664 9540 22995 9568
rect 21836 9472 22416 9500
rect 22388 9441 22416 9472
rect 22373 9435 22431 9441
rect 18984 9404 19748 9432
rect 20732 9404 22324 9432
rect 18984 9364 19012 9404
rect 19720 9376 19748 9404
rect 14108 9336 19012 9364
rect 19337 9367 19395 9373
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 19518 9364 19524 9376
rect 19383 9336 19524 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19702 9324 19708 9376
rect 19760 9324 19766 9376
rect 21913 9367 21971 9373
rect 21913 9333 21925 9367
rect 21959 9364 21971 9367
rect 22094 9364 22100 9376
rect 21959 9336 22100 9364
rect 21959 9333 21971 9336
rect 21913 9327 21971 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 22186 9324 22192 9376
rect 22244 9324 22250 9376
rect 22296 9364 22324 9404
rect 22373 9401 22385 9435
rect 22419 9401 22431 9435
rect 22373 9395 22431 9401
rect 22664 9364 22692 9540
rect 22983 9537 22995 9540
rect 23029 9537 23041 9571
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 22983 9531 23041 9537
rect 23768 9540 24317 9568
rect 22741 9503 22799 9509
rect 22741 9469 22753 9503
rect 22787 9469 22799 9503
rect 22741 9463 22799 9469
rect 22296 9336 22692 9364
rect 22756 9364 22784 9463
rect 23768 9441 23796 9540
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 24578 9460 24584 9512
rect 24636 9460 24642 9512
rect 23753 9435 23811 9441
rect 23753 9401 23765 9435
rect 23799 9401 23811 9435
rect 24596 9432 24624 9460
rect 23753 9395 23811 9401
rect 23860 9404 24624 9432
rect 23014 9364 23020 9376
rect 22756 9336 23020 9364
rect 23014 9324 23020 9336
rect 23072 9364 23078 9376
rect 23860 9364 23888 9404
rect 23072 9336 23888 9364
rect 23072 9324 23078 9336
rect 24118 9324 24124 9376
rect 24176 9324 24182 9376
rect 1104 9274 24840 9296
rect 1104 9222 3917 9274
rect 3969 9222 3981 9274
rect 4033 9222 4045 9274
rect 4097 9222 4109 9274
rect 4161 9222 4173 9274
rect 4225 9222 9851 9274
rect 9903 9222 9915 9274
rect 9967 9222 9979 9274
rect 10031 9222 10043 9274
rect 10095 9222 10107 9274
rect 10159 9222 15785 9274
rect 15837 9222 15849 9274
rect 15901 9222 15913 9274
rect 15965 9222 15977 9274
rect 16029 9222 16041 9274
rect 16093 9222 21719 9274
rect 21771 9222 21783 9274
rect 21835 9222 21847 9274
rect 21899 9222 21911 9274
rect 21963 9222 21975 9274
rect 22027 9222 24840 9274
rect 1104 9200 24840 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 1360 9132 2697 9160
rect 1360 9120 1366 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 2685 9123 2743 9129
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 3108 9132 3188 9160
rect 3108 9120 3114 9132
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 1673 9095 1731 9101
rect 1673 9092 1685 9095
rect 1544 9064 1685 9092
rect 1544 9052 1550 9064
rect 1673 9061 1685 9064
rect 1719 9061 1731 9095
rect 1673 9055 1731 9061
rect 2222 9052 2228 9104
rect 2280 9052 2286 9104
rect 934 8984 940 9036
rect 992 9024 998 9036
rect 992 8996 2268 9024
rect 992 8984 998 8996
rect 1946 8916 1952 8968
rect 2004 8956 2010 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 2004 8928 2053 8956
rect 2004 8916 2010 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 1489 8891 1547 8897
rect 1489 8857 1501 8891
rect 1535 8888 1547 8891
rect 1854 8888 1860 8900
rect 1535 8860 1860 8888
rect 1535 8857 1547 8860
rect 1489 8851 1547 8857
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 2240 8820 2268 8996
rect 3160 8965 3188 9132
rect 3234 9120 3240 9172
rect 3292 9160 3298 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3292 9132 4077 9160
rect 3292 9120 3298 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 7834 9160 7840 9172
rect 7524 9132 7840 9160
rect 7524 9120 7530 9132
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 9582 9160 9588 9172
rect 8527 9132 9588 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9784 9132 10548 9160
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9784 9033 9812 9132
rect 10520 9092 10548 9132
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10781 9163 10839 9169
rect 10781 9160 10793 9163
rect 10652 9132 10793 9160
rect 10652 9120 10658 9132
rect 10781 9129 10793 9132
rect 10827 9129 10839 9163
rect 17218 9160 17224 9172
rect 10781 9123 10839 9129
rect 16868 9132 17224 9160
rect 10520 9064 13952 9092
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 9088 8996 9781 9024
rect 9088 8984 9094 8996
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 11256 8996 13676 9024
rect 3145 8959 3203 8965
rect 2424 8928 2774 8956
rect 2424 8900 2452 8928
rect 2406 8848 2412 8900
rect 2464 8848 2470 8900
rect 2590 8848 2596 8900
rect 2648 8848 2654 8900
rect 2746 8888 2774 8928
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3476 8928 3985 8956
rect 3476 8916 3482 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4264 8888 4292 8919
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 7743 8959 7801 8965
rect 7743 8925 7755 8959
rect 7789 8956 7801 8959
rect 7834 8956 7840 8968
rect 7789 8928 7840 8956
rect 7789 8925 7801 8928
rect 7743 8919 7801 8925
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 10043 8959 10101 8965
rect 10043 8925 10055 8959
rect 10089 8956 10101 8959
rect 11256 8956 11284 8996
rect 10089 8928 11284 8956
rect 10089 8925 10101 8928
rect 10043 8919 10101 8925
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 13538 8956 13544 8968
rect 12492 8928 13544 8956
rect 12492 8916 12498 8928
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13262 8888 13268 8900
rect 2746 8860 3832 8888
rect 4264 8860 13268 8888
rect 3804 8829 3832 8860
rect 13262 8848 13268 8860
rect 13320 8848 13326 8900
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 2240 8792 3249 8820
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 8478 8780 8484 8832
rect 8536 8820 8542 8832
rect 12434 8820 12440 8832
rect 8536 8792 12440 8820
rect 8536 8780 8542 8792
rect 12434 8780 12440 8792
rect 12492 8780 12498 8832
rect 13648 8820 13676 8996
rect 13924 8888 13952 9064
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14093 9027 14151 9033
rect 14093 9024 14105 9027
rect 14056 8996 14105 9024
rect 14056 8984 14062 8996
rect 14093 8993 14105 8996
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 14366 8965 14372 8968
rect 14335 8959 14372 8965
rect 14335 8925 14347 8959
rect 14335 8919 14372 8925
rect 14366 8916 14372 8919
rect 14424 8916 14430 8968
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8925 15531 8959
rect 15746 8956 15752 8968
rect 15707 8928 15752 8956
rect 15473 8919 15531 8925
rect 15488 8888 15516 8919
rect 15746 8916 15752 8928
rect 15804 8916 15810 8968
rect 16868 8965 16896 9132
rect 17218 9120 17224 9132
rect 17276 9160 17282 9172
rect 17276 9132 17632 9160
rect 17276 9120 17282 9132
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 15856 8928 16865 8956
rect 15856 8888 15884 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 17095 8959 17153 8965
rect 17095 8925 17107 8959
rect 17141 8925 17153 8959
rect 17095 8919 17153 8925
rect 17110 8888 17138 8919
rect 13924 8860 15884 8888
rect 16132 8860 17138 8888
rect 17604 8888 17632 9132
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 17736 9132 22416 9160
rect 17736 9120 17742 9132
rect 22388 9092 22416 9132
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22520 9132 22661 9160
rect 22520 9120 22526 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 23290 9120 23296 9172
rect 23348 9160 23354 9172
rect 23385 9163 23443 9169
rect 23385 9160 23397 9163
rect 23348 9132 23397 9160
rect 23348 9120 23354 9132
rect 23385 9129 23397 9132
rect 23431 9129 23443 9163
rect 23385 9123 23443 9129
rect 23937 9163 23995 9169
rect 23937 9129 23949 9163
rect 23983 9160 23995 9163
rect 24026 9160 24032 9172
rect 23983 9132 24032 9160
rect 23983 9129 23995 9132
rect 23937 9123 23995 9129
rect 24026 9120 24032 9132
rect 24084 9120 24090 9172
rect 24118 9120 24124 9172
rect 24176 9120 24182 9172
rect 22388 9064 23980 9092
rect 23952 9036 23980 9064
rect 19610 8984 19616 9036
rect 19668 9024 19674 9036
rect 21266 9024 21272 9036
rect 19668 8996 21272 9024
rect 19668 8984 19674 8996
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 23842 9024 23848 9036
rect 22480 8996 23848 9024
rect 19150 8916 19156 8968
rect 19208 8956 19214 8968
rect 22480 8956 22508 8996
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 23934 8984 23940 9036
rect 23992 8984 23998 9036
rect 19208 8928 22508 8956
rect 19208 8916 19214 8928
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23566 8956 23572 8968
rect 22971 8928 23572 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8956 23719 8959
rect 24136 8956 24164 9120
rect 23707 8928 24164 8956
rect 23707 8925 23719 8928
rect 23661 8919 23719 8925
rect 20438 8888 20444 8900
rect 17604 8860 20444 8888
rect 16132 8832 16160 8860
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 21536 8891 21594 8897
rect 21536 8857 21548 8891
rect 21582 8888 21594 8891
rect 22370 8888 22376 8900
rect 21582 8860 22376 8888
rect 21582 8857 21594 8860
rect 21536 8851 21594 8857
rect 22370 8848 22376 8860
rect 22428 8888 22434 8900
rect 22572 8888 22600 8916
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 22428 8860 22508 8888
rect 22572 8860 23121 8888
rect 22428 8848 22434 8860
rect 14826 8820 14832 8832
rect 13648 8792 14832 8820
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 15102 8780 15108 8832
rect 15160 8780 15166 8832
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 16482 8780 16488 8832
rect 16540 8780 16546 8832
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17184 8792 17877 8820
rect 17184 8780 17190 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 17865 8783 17923 8789
rect 17954 8780 17960 8832
rect 18012 8820 18018 8832
rect 22002 8820 22008 8832
rect 18012 8792 22008 8820
rect 18012 8780 18018 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 22480 8820 22508 8860
rect 23109 8857 23121 8860
rect 23155 8857 23167 8891
rect 23109 8851 23167 8857
rect 22741 8823 22799 8829
rect 22741 8820 22753 8823
rect 22480 8792 22753 8820
rect 22741 8789 22753 8792
rect 22787 8789 22799 8823
rect 22741 8783 22799 8789
rect 1104 8730 25000 8752
rect 1104 8678 6884 8730
rect 6936 8678 6948 8730
rect 7000 8678 7012 8730
rect 7064 8678 7076 8730
rect 7128 8678 7140 8730
rect 7192 8678 12818 8730
rect 12870 8678 12882 8730
rect 12934 8678 12946 8730
rect 12998 8678 13010 8730
rect 13062 8678 13074 8730
rect 13126 8678 18752 8730
rect 18804 8678 18816 8730
rect 18868 8678 18880 8730
rect 18932 8678 18944 8730
rect 18996 8678 19008 8730
rect 19060 8678 24686 8730
rect 24738 8678 24750 8730
rect 24802 8678 24814 8730
rect 24866 8678 24878 8730
rect 24930 8678 24942 8730
rect 24994 8678 25000 8730
rect 1104 8656 25000 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 1268 8588 2697 8616
rect 1268 8576 1274 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 7101 8619 7159 8625
rect 7101 8585 7113 8619
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 1486 8508 1492 8560
rect 1544 8508 1550 8560
rect 1670 8508 1676 8560
rect 1728 8548 1734 8560
rect 2409 8551 2467 8557
rect 2409 8548 2421 8551
rect 1728 8520 2421 8548
rect 1728 8508 1734 8520
rect 2409 8517 2421 8520
rect 2455 8517 2467 8551
rect 2409 8511 2467 8517
rect 2593 8551 2651 8557
rect 2593 8517 2605 8551
rect 2639 8548 2651 8551
rect 7116 8548 7144 8579
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 8168 8588 8401 8616
rect 8168 8576 8174 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8389 8579 8447 8585
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10318 8616 10324 8628
rect 10183 8588 10324 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 12066 8616 12072 8628
rect 10928 8588 12072 8616
rect 10928 8576 10934 8588
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 12989 8619 13047 8625
rect 12989 8616 13001 8619
rect 12492 8588 13001 8616
rect 12492 8576 12498 8588
rect 12989 8585 13001 8588
rect 13035 8585 13047 8619
rect 12989 8579 13047 8585
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 13722 8616 13728 8628
rect 13596 8588 13728 8616
rect 13596 8576 13602 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 15102 8616 15108 8628
rect 14200 8588 15108 8616
rect 7466 8548 7472 8560
rect 2639 8520 7144 8548
rect 7392 8520 7472 8548
rect 2639 8517 2651 8520
rect 2593 8511 2651 8517
rect 1854 8440 1860 8492
rect 1912 8440 1918 8492
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2056 8276 2084 8443
rect 2222 8440 2228 8492
rect 2280 8480 2286 8492
rect 3145 8483 3203 8489
rect 3145 8480 3157 8483
rect 2280 8452 3157 8480
rect 2280 8440 2286 8452
rect 3145 8449 3157 8452
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 2372 8384 3924 8412
rect 2372 8372 2378 8384
rect 3326 8304 3332 8356
rect 3384 8304 3390 8356
rect 3896 8353 3924 8384
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 7392 8421 7420 8520
rect 7466 8508 7472 8520
rect 7524 8508 7530 8560
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11664 8520 11713 8548
rect 11664 8508 11670 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 12710 8548 12716 8560
rect 11701 8511 11759 8517
rect 11806 8520 12716 8548
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7651 8483 7709 8489
rect 7651 8480 7663 8483
rect 7616 8452 7663 8480
rect 7616 8440 7622 8452
rect 7651 8449 7663 8452
rect 7697 8480 7709 8483
rect 8018 8480 8024 8492
rect 7697 8452 8024 8480
rect 7697 8449 7709 8452
rect 7651 8443 7709 8449
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8294 8440 8300 8492
rect 8352 8480 8358 8492
rect 9367 8483 9425 8489
rect 9367 8480 9379 8483
rect 8352 8452 9379 8480
rect 8352 8440 8358 8452
rect 9367 8449 9379 8452
rect 9413 8480 9425 8483
rect 11806 8480 11834 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8517 12863 8551
rect 12805 8511 12863 8517
rect 9413 8452 11834 8480
rect 9413 8449 9425 8452
rect 9367 8443 9425 8449
rect 11974 8440 11980 8492
rect 12032 8440 12038 8492
rect 12066 8440 12072 8492
rect 12124 8440 12130 8492
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12342 8480 12348 8492
rect 12216 8452 12348 8480
rect 12216 8440 12222 8452
rect 12342 8440 12348 8452
rect 12400 8480 12406 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12400 8452 12449 8480
rect 12400 8440 12406 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12820 8480 12848 8511
rect 13446 8508 13452 8560
rect 13504 8548 13510 8560
rect 14200 8557 14228 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 17034 8616 17040 8628
rect 16356 8588 17040 8616
rect 16356 8576 16362 8588
rect 17034 8576 17040 8588
rect 17092 8616 17098 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 17092 8588 17141 8616
rect 17092 8576 17098 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 17129 8579 17187 8585
rect 17512 8588 19625 8616
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13504 8520 13829 8548
rect 13504 8508 13510 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 14185 8551 14243 8557
rect 14185 8517 14197 8551
rect 14231 8517 14243 8551
rect 14185 8511 14243 8517
rect 14921 8551 14979 8557
rect 14921 8517 14933 8551
rect 14967 8517 14979 8551
rect 14921 8511 14979 8517
rect 12584 8452 12848 8480
rect 12584 8440 12590 8452
rect 13906 8440 13912 8492
rect 13964 8480 13970 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13964 8452 14105 8480
rect 13964 8440 13970 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14642 8480 14648 8492
rect 14599 8452 14648 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 14936 8480 14964 8511
rect 15654 8508 15660 8560
rect 15712 8508 15718 8560
rect 17310 8508 17316 8560
rect 17368 8548 17374 8560
rect 17512 8557 17540 8588
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19613 8579 19671 8585
rect 22094 8576 22100 8628
rect 22152 8576 22158 8628
rect 22186 8576 22192 8628
rect 22244 8576 22250 8628
rect 23750 8576 23756 8628
rect 23808 8576 23814 8628
rect 17405 8551 17463 8557
rect 17405 8548 17417 8551
rect 17368 8520 17417 8548
rect 17368 8508 17374 8520
rect 17405 8517 17417 8520
rect 17451 8517 17463 8551
rect 17405 8511 17463 8517
rect 17497 8551 17555 8557
rect 17497 8517 17509 8551
rect 17543 8517 17555 8551
rect 18233 8551 18291 8557
rect 18233 8548 18245 8551
rect 17497 8511 17555 8517
rect 17604 8520 18245 8548
rect 14792 8452 14964 8480
rect 15672 8480 15700 8508
rect 17604 8480 17632 8520
rect 18233 8517 18245 8520
rect 18279 8548 18291 8551
rect 18598 8548 18604 8560
rect 18279 8520 18604 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 15672 8452 17632 8480
rect 14792 8440 14798 8452
rect 17862 8440 17868 8492
rect 17920 8440 17926 8492
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 18843 8483 18901 8489
rect 18843 8480 18855 8483
rect 18380 8452 18855 8480
rect 18380 8440 18386 8452
rect 18843 8449 18855 8452
rect 18889 8480 18901 8483
rect 19334 8480 19340 8492
rect 18889 8452 19340 8480
rect 18889 8449 18901 8452
rect 18843 8443 18901 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19576 8452 19993 8480
rect 19576 8440 19582 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 20162 8440 20168 8492
rect 20220 8440 20226 8492
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 22112 8480 22140 8576
rect 22204 8548 22232 8576
rect 23768 8548 23796 8576
rect 22204 8520 22692 8548
rect 23768 8520 24532 8548
rect 22664 8489 22692 8520
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22112 8452 22201 8480
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22189 8443 22247 8449
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 23014 8440 23020 8492
rect 23072 8480 23078 8492
rect 23477 8483 23535 8489
rect 23477 8480 23489 8483
rect 23072 8452 23489 8480
rect 23072 8440 23078 8452
rect 23477 8449 23489 8452
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 24504 8489 24532 8520
rect 24489 8483 24547 8489
rect 24489 8449 24501 8483
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 13820 8424 13872 8430
rect 18144 8424 18196 8430
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 6144 8384 7389 8412
rect 6144 8372 6150 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7377 8375 7435 8381
rect 9030 8372 9036 8424
rect 9088 8412 9094 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 9088 8384 9137 8412
rect 9088 8372 9094 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 11146 8372 11152 8424
rect 11204 8412 11210 8424
rect 11204 8384 11546 8412
rect 11204 8372 11210 8384
rect 15562 8372 15568 8424
rect 15620 8372 15626 8424
rect 18601 8415 18659 8421
rect 18601 8381 18613 8415
rect 18647 8381 18659 8415
rect 21100 8412 21128 8440
rect 18601 8375 18659 8381
rect 19306 8384 21128 8412
rect 22005 8415 22063 8421
rect 13820 8366 13872 8372
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 8110 8304 8116 8356
rect 8168 8344 8174 8356
rect 8386 8344 8392 8356
rect 8168 8316 8392 8344
rect 8168 8304 8174 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 15105 8347 15163 8353
rect 15105 8313 15117 8347
rect 15151 8344 15163 8347
rect 15580 8344 15608 8372
rect 18144 8366 18196 8372
rect 15151 8316 15608 8344
rect 18616 8344 18644 8375
rect 18616 8316 18736 8344
rect 15151 8313 15163 8316
rect 15105 8307 15163 8313
rect 18708 8288 18736 8316
rect 2314 8276 2320 8288
rect 2056 8248 2320 8276
rect 2314 8236 2320 8248
rect 2372 8236 2378 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 4890 8276 4896 8288
rect 2740 8248 4896 8276
rect 2740 8236 2746 8248
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 11238 8276 11244 8288
rect 7248 8248 11244 8276
rect 7248 8236 7254 8248
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13262 8276 13268 8288
rect 13044 8248 13268 8276
rect 13044 8236 13050 8248
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 18414 8236 18420 8288
rect 18472 8236 18478 8288
rect 18690 8236 18696 8288
rect 18748 8276 18754 8288
rect 19306 8276 19334 8384
rect 22005 8381 22017 8415
rect 22051 8412 22063 8415
rect 22278 8412 22284 8424
rect 22051 8384 22284 8412
rect 22051 8381 22063 8384
rect 22005 8375 22063 8381
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23339 8384 23520 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23492 8356 23520 8384
rect 23934 8372 23940 8424
rect 23992 8372 23998 8424
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 22649 8347 22707 8353
rect 22649 8344 22661 8347
rect 19760 8316 22661 8344
rect 19760 8304 19766 8316
rect 22649 8313 22661 8316
rect 22695 8313 22707 8347
rect 22649 8307 22707 8313
rect 23474 8304 23480 8356
rect 23532 8304 23538 8356
rect 18748 8248 19334 8276
rect 18748 8236 18754 8248
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20073 8279 20131 8285
rect 20073 8276 20085 8279
rect 20036 8248 20085 8276
rect 20036 8236 20042 8248
rect 20073 8245 20085 8248
rect 20119 8245 20131 8279
rect 20073 8239 20131 8245
rect 22922 8236 22928 8288
rect 22980 8276 22986 8288
rect 23198 8276 23204 8288
rect 22980 8248 23204 8276
rect 22980 8236 22986 8248
rect 23198 8236 23204 8248
rect 23256 8236 23262 8288
rect 24302 8236 24308 8288
rect 24360 8236 24366 8288
rect 1104 8186 24840 8208
rect 1104 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 9851 8186
rect 9903 8134 9915 8186
rect 9967 8134 9979 8186
rect 10031 8134 10043 8186
rect 10095 8134 10107 8186
rect 10159 8134 15785 8186
rect 15837 8134 15849 8186
rect 15901 8134 15913 8186
rect 15965 8134 15977 8186
rect 16029 8134 16041 8186
rect 16093 8134 21719 8186
rect 21771 8134 21783 8186
rect 21835 8134 21847 8186
rect 21899 8134 21911 8186
rect 21963 8134 21975 8186
rect 22027 8134 24840 8186
rect 1104 8112 24840 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1452 8044 1593 8072
rect 1452 8032 1458 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2222 8072 2228 8084
rect 1912 8044 2228 8072
rect 1912 8032 1918 8044
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 2372 8044 3341 8072
rect 2372 8032 2378 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 5350 8072 5356 8084
rect 3329 8035 3387 8041
rect 3896 8044 5356 8072
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 2832 7976 3801 8004
rect 2832 7964 2838 7976
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 2682 7896 2688 7948
rect 2740 7896 2746 7948
rect 3896 7936 3924 8044
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 7190 8072 7196 8084
rect 5828 8044 7196 8072
rect 3344 7908 3924 7936
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 1949 7831 2007 7837
rect 1486 7760 1492 7812
rect 1544 7760 1550 7812
rect 1670 7760 1676 7812
rect 1728 7760 1734 7812
rect 1964 7800 1992 7831
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2314 7800 2320 7812
rect 1964 7772 2320 7800
rect 2314 7760 2320 7772
rect 2372 7800 2378 7812
rect 2700 7800 2728 7896
rect 3344 7880 3372 7908
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4154 7868 4160 7880
rect 4019 7840 4160 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 2372 7772 2728 7800
rect 3528 7800 3556 7831
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4246 7828 4252 7880
rect 4304 7828 4310 7880
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4396 7840 4905 7868
rect 4396 7828 4402 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5167 7871 5225 7877
rect 5167 7837 5179 7871
rect 5213 7868 5225 7871
rect 5828 7868 5856 8044
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7340 8044 8125 8072
rect 7340 8032 7346 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11146 8072 11152 8084
rect 10919 8044 11152 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11296 8044 11928 8072
rect 11296 8032 11302 8044
rect 5905 8007 5963 8013
rect 5905 7973 5917 8007
rect 5951 8004 5963 8007
rect 6917 8007 6975 8013
rect 6917 8004 6929 8007
rect 5951 7976 6929 8004
rect 5951 7973 5963 7976
rect 5905 7967 5963 7973
rect 6917 7973 6929 7976
rect 6963 7973 6975 8007
rect 6917 7967 6975 7973
rect 6270 7896 6276 7948
rect 6328 7896 6334 7948
rect 7190 7896 7196 7948
rect 7248 7896 7254 7948
rect 9766 7936 9772 7948
rect 7392 7908 9772 7936
rect 7392 7880 7420 7908
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 11900 7936 11928 8044
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 12124 8044 12265 8072
rect 12124 8032 12130 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13814 8072 13820 8084
rect 13679 8044 13820 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 16482 8072 16488 8084
rect 15948 8044 16488 8072
rect 15948 8013 15976 8044
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 16908 8044 17908 8072
rect 16908 8032 16914 8044
rect 15933 8007 15991 8013
rect 15933 7973 15945 8007
rect 15979 7973 15991 8007
rect 17880 8004 17908 8044
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 18196 8044 18245 8072
rect 18196 8032 18202 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 18233 8035 18291 8041
rect 18598 8032 18604 8084
rect 18656 8072 18662 8084
rect 19889 8075 19947 8081
rect 18656 8044 19564 8072
rect 18656 8032 18662 8044
rect 19429 8007 19487 8013
rect 19429 8004 19441 8007
rect 17880 7976 19441 8004
rect 15933 7967 15991 7973
rect 19429 7973 19441 7976
rect 19475 7973 19487 8007
rect 19536 8004 19564 8044
rect 19889 8041 19901 8075
rect 19935 8072 19947 8075
rect 20162 8072 20168 8084
rect 19935 8044 20168 8072
rect 19935 8041 19947 8044
rect 19889 8035 19947 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 22649 8075 22707 8081
rect 22649 8041 22661 8075
rect 22695 8072 22707 8075
rect 23014 8072 23020 8084
rect 22695 8044 23020 8072
rect 22695 8041 22707 8044
rect 22649 8035 22707 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 21085 8007 21143 8013
rect 21085 8004 21097 8007
rect 19536 7976 21097 8004
rect 19429 7967 19487 7973
rect 21085 7973 21097 7976
rect 21131 7973 21143 8007
rect 21085 7967 21143 7973
rect 11900 7908 12388 7936
rect 5213 7840 5856 7868
rect 5213 7837 5225 7840
rect 5167 7831 5225 7837
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 7374 7877 7380 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6420 7840 6469 7868
rect 6420 7828 6426 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 7331 7871 7380 7877
rect 7331 7837 7343 7871
rect 7377 7837 7380 7871
rect 7331 7831 7380 7837
rect 7374 7828 7380 7831
rect 7432 7828 7438 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 10135 7871 10193 7877
rect 10135 7837 10147 7871
rect 10181 7868 10193 7871
rect 10778 7868 10784 7880
rect 10181 7840 10784 7868
rect 10181 7837 10193 7840
rect 10135 7831 10193 7837
rect 3528 7772 6500 7800
rect 2372 7760 2378 7772
rect 1688 7732 1716 7760
rect 2406 7732 2412 7744
rect 1688 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3200 7704 4077 7732
rect 3200 7692 3206 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4065 7695 4123 7701
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 5166 7732 5172 7744
rect 4488 7704 5172 7732
rect 4488 7692 4494 7704
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 6472 7732 6500 7772
rect 8018 7760 8024 7812
rect 8076 7800 8082 7812
rect 9214 7800 9220 7812
rect 8076 7772 9220 7800
rect 8076 7760 8082 7772
rect 9214 7760 9220 7772
rect 9272 7760 9278 7812
rect 9876 7800 9904 7831
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 11515 7871 11573 7877
rect 11515 7837 11527 7871
rect 11561 7868 11573 7871
rect 12250 7868 12256 7880
rect 11561 7840 12256 7868
rect 11561 7837 11573 7840
rect 11515 7831 11573 7837
rect 11256 7800 11284 7831
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 12360 7868 12388 7908
rect 12618 7896 12624 7948
rect 12676 7896 12682 7948
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 16326 7939 16384 7945
rect 16326 7936 16338 7939
rect 15620 7908 16338 7936
rect 15620 7896 15626 7908
rect 16326 7905 16338 7908
rect 16372 7905 16384 7939
rect 16326 7899 16384 7905
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 17126 7936 17132 7948
rect 16531 7908 17132 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 18923 7908 19472 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 12863 7871 12921 7877
rect 12863 7868 12875 7871
rect 12360 7840 12875 7868
rect 12863 7837 12875 7840
rect 12909 7837 12921 7871
rect 12863 7831 12921 7837
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 15289 7871 15347 7877
rect 13044 7840 14780 7868
rect 13044 7828 13050 7840
rect 13354 7800 13360 7812
rect 9876 7772 13360 7800
rect 11716 7744 11744 7772
rect 13354 7760 13360 7772
rect 13412 7760 13418 7812
rect 8478 7732 8484 7744
rect 6472 7704 8484 7732
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 11698 7692 11704 7744
rect 11756 7692 11762 7744
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 13722 7732 13728 7744
rect 12124 7704 13728 7732
rect 12124 7692 12130 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14752 7732 14780 7840
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15378 7868 15384 7880
rect 15335 7840 15384 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 15473 7871 15531 7877
rect 15473 7837 15485 7871
rect 15519 7868 15531 7871
rect 15654 7868 15660 7880
rect 15519 7840 15660 7868
rect 15519 7837 15531 7840
rect 15473 7831 15531 7837
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 16206 7828 16212 7880
rect 16264 7828 16270 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7837 17279 7871
rect 17221 7831 17279 7837
rect 17479 7841 17537 7847
rect 17236 7744 17264 7831
rect 17479 7807 17491 7841
rect 17525 7838 17537 7841
rect 17525 7807 17540 7838
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 19444 7877 19472 7908
rect 21266 7896 21272 7948
rect 21324 7936 21330 7948
rect 21324 7908 22876 7936
rect 21324 7896 21330 7908
rect 22848 7880 22876 7908
rect 18785 7871 18843 7877
rect 18785 7868 18797 7871
rect 18656 7840 18797 7868
rect 18656 7828 18662 7840
rect 18785 7837 18797 7840
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19576 7840 19625 7868
rect 19576 7828 19582 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19944 7840 20085 7868
rect 19944 7828 19950 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 22465 7871 22523 7877
rect 22465 7837 22477 7871
rect 22511 7837 22523 7871
rect 22465 7831 22523 7837
rect 17479 7801 17540 7807
rect 17512 7800 17540 7801
rect 17770 7800 17776 7812
rect 17512 7772 17776 7800
rect 17770 7760 17776 7772
rect 17828 7760 17834 7812
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7800 19855 7803
rect 19978 7800 19984 7812
rect 19843 7772 19984 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 22480 7800 22508 7831
rect 22554 7828 22560 7880
rect 22612 7828 22618 7880
rect 22830 7828 22836 7880
rect 22888 7828 22894 7880
rect 23100 7803 23158 7809
rect 22480 7772 22784 7800
rect 17129 7735 17187 7741
rect 17129 7732 17141 7735
rect 14752 7704 17141 7732
rect 17129 7701 17141 7704
rect 17175 7701 17187 7735
rect 17129 7695 17187 7701
rect 17218 7692 17224 7744
rect 17276 7732 17282 7744
rect 18690 7732 18696 7744
rect 17276 7704 18696 7732
rect 17276 7692 17282 7704
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 20898 7692 20904 7744
rect 20956 7732 20962 7744
rect 21358 7732 21364 7744
rect 20956 7704 21364 7732
rect 20956 7692 20962 7704
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 22094 7692 22100 7744
rect 22152 7732 22158 7744
rect 22281 7735 22339 7741
rect 22281 7732 22293 7735
rect 22152 7704 22293 7732
rect 22152 7692 22158 7704
rect 22281 7701 22293 7704
rect 22327 7701 22339 7735
rect 22756 7732 22784 7772
rect 23100 7769 23112 7803
rect 23146 7800 23158 7803
rect 23750 7800 23756 7812
rect 23146 7772 23756 7800
rect 23146 7769 23158 7772
rect 23100 7763 23158 7769
rect 23750 7760 23756 7772
rect 23808 7760 23814 7812
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 22756 7704 24225 7732
rect 22281 7695 22339 7701
rect 24213 7701 24225 7704
rect 24259 7701 24271 7735
rect 24213 7695 24271 7701
rect 1104 7642 25000 7664
rect 1104 7590 6884 7642
rect 6936 7590 6948 7642
rect 7000 7590 7012 7642
rect 7064 7590 7076 7642
rect 7128 7590 7140 7642
rect 7192 7590 12818 7642
rect 12870 7590 12882 7642
rect 12934 7590 12946 7642
rect 12998 7590 13010 7642
rect 13062 7590 13074 7642
rect 13126 7590 18752 7642
rect 18804 7590 18816 7642
rect 18868 7590 18880 7642
rect 18932 7590 18944 7642
rect 18996 7590 19008 7642
rect 19060 7590 24686 7642
rect 24738 7590 24750 7642
rect 24802 7590 24814 7642
rect 24866 7590 24878 7642
rect 24930 7590 24942 7642
rect 24994 7590 25000 7642
rect 1104 7568 25000 7590
rect 750 7488 756 7540
rect 808 7528 814 7540
rect 1118 7528 1124 7540
rect 808 7500 1124 7528
rect 808 7488 814 7500
rect 1118 7488 1124 7500
rect 1176 7488 1182 7540
rect 1762 7488 1768 7540
rect 1820 7488 1826 7540
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2590 7528 2596 7540
rect 2179 7500 2596 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 2832 7500 4108 7528
rect 2832 7488 2838 7500
rect 1670 7420 1676 7472
rect 1728 7420 1734 7472
rect 4080 7460 4108 7500
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4249 7531 4307 7537
rect 4249 7528 4261 7531
rect 4212 7500 4261 7528
rect 4212 7488 4218 7500
rect 4249 7497 4261 7500
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 4356 7500 6040 7528
rect 4356 7460 4384 7500
rect 1780 7432 2452 7460
rect 4080 7432 4384 7460
rect 6012 7460 6040 7500
rect 7466 7488 7472 7540
rect 7524 7488 7530 7540
rect 7576 7500 8432 7528
rect 7576 7460 7604 7500
rect 6012 7432 7604 7460
rect 8404 7460 8432 7500
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 18414 7528 18420 7540
rect 8536 7500 18420 7528
rect 8536 7488 8542 7500
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 19521 7531 19579 7537
rect 19521 7497 19533 7531
rect 19567 7528 19579 7531
rect 19886 7528 19892 7540
rect 19567 7500 19892 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7528 20039 7531
rect 20622 7528 20628 7540
rect 20027 7500 20628 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 21545 7531 21603 7537
rect 21545 7497 21557 7531
rect 21591 7528 21603 7531
rect 21591 7500 22048 7528
rect 21591 7497 21603 7500
rect 21545 7491 21603 7497
rect 8404 7432 12572 7460
rect 474 7352 480 7404
rect 532 7392 538 7404
rect 1780 7392 1808 7432
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 532 7364 1808 7392
rect 2056 7364 2329 7392
rect 532 7352 538 7364
rect 2056 7188 2084 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 2424 7336 2452 7432
rect 8279 7425 8337 7431
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2774 7392 2780 7404
rect 2593 7355 2651 7361
rect 2406 7284 2412 7336
rect 2464 7284 2470 7336
rect 2130 7216 2136 7268
rect 2188 7256 2194 7268
rect 2608 7256 2636 7355
rect 2746 7352 2780 7392
rect 2832 7352 2838 7404
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 5442 7401 5448 7404
rect 5399 7395 5448 7401
rect 5399 7361 5411 7395
rect 5445 7361 5448 7395
rect 5399 7355 5448 7361
rect 5442 7352 5448 7355
rect 5500 7352 5506 7404
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6731 7395 6789 7401
rect 6731 7361 6743 7395
rect 6777 7392 6789 7395
rect 6777 7364 7972 7392
rect 8279 7391 8291 7425
rect 8325 7422 8337 7425
rect 8325 7392 8340 7422
rect 8846 7392 8852 7404
rect 8325 7391 8852 7392
rect 8279 7385 8852 7391
rect 8312 7364 8852 7385
rect 6777 7361 6789 7364
rect 6731 7355 6789 7361
rect 2746 7256 2774 7352
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 3016 7296 3065 7324
rect 3016 7284 3022 7296
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 3467 7327 3525 7333
rect 3467 7293 3479 7327
rect 3513 7324 3525 7327
rect 3786 7324 3792 7336
rect 3513 7296 3792 7324
rect 3513 7293 3525 7296
rect 3467 7287 3525 7293
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 4430 7324 4436 7336
rect 4387 7296 4436 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7324 4583 7327
rect 4614 7324 4620 7336
rect 4571 7296 4620 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4614 7284 4620 7296
rect 4672 7284 4678 7336
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 5132 7296 5273 7324
rect 5132 7284 5138 7296
rect 5261 7293 5273 7296
rect 5307 7324 5319 7327
rect 6196 7324 6224 7352
rect 5307 7296 6224 7324
rect 6457 7327 6515 7333
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 6457 7293 6469 7327
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 2188 7228 2774 7256
rect 2188 7216 2194 7228
rect 4982 7216 4988 7268
rect 5040 7216 5046 7268
rect 6086 7216 6092 7268
rect 6144 7256 6150 7268
rect 6472 7256 6500 7287
rect 6144 7228 6500 7256
rect 6144 7216 6150 7228
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 2056 7160 6193 7188
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 7944 7188 7972 7364
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9272 7364 9413 7392
rect 9272 7352 9278 7364
rect 9401 7361 9413 7364
rect 9447 7392 9459 7395
rect 9582 7392 9588 7404
rect 9447 7364 9588 7392
rect 9447 7361 9459 7364
rect 9401 7355 9459 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 9675 7395 9733 7401
rect 9675 7361 9687 7395
rect 9721 7392 9733 7395
rect 10962 7392 10968 7404
rect 9721 7364 10968 7392
rect 9721 7361 9733 7364
rect 9675 7355 9733 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 8018 7284 8024 7336
rect 8076 7284 8082 7336
rect 10226 7284 10232 7336
rect 10284 7324 10290 7336
rect 12434 7324 12440 7336
rect 10284 7296 12440 7324
rect 10284 7284 10290 7296
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 11054 7256 11060 7268
rect 10060 7228 11060 7256
rect 8938 7188 8944 7200
rect 7944 7160 8944 7188
rect 6181 7151 6239 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 9030 7148 9036 7200
rect 9088 7148 9094 7200
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 10060 7188 10088 7228
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 12544 7256 12572 7432
rect 12618 7420 12624 7472
rect 12676 7460 12682 7472
rect 13265 7463 13323 7469
rect 13265 7460 13277 7463
rect 12676 7432 13277 7460
rect 12676 7420 12682 7432
rect 13265 7429 13277 7432
rect 13311 7460 13323 7463
rect 13446 7460 13452 7472
rect 13311 7432 13452 7460
rect 13311 7429 13323 7432
rect 13265 7423 13323 7429
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 13541 7463 13599 7469
rect 13541 7429 13553 7463
rect 13587 7460 13599 7463
rect 13814 7460 13820 7472
rect 13587 7432 13820 7460
rect 13587 7429 13599 7432
rect 13541 7423 13599 7429
rect 13814 7420 13820 7432
rect 13872 7420 13878 7472
rect 14369 7463 14427 7469
rect 14369 7429 14381 7463
rect 14415 7460 14427 7463
rect 14734 7460 14740 7472
rect 14415 7432 14740 7460
rect 14415 7429 14427 7432
rect 14369 7423 14427 7429
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 18156 7432 19334 7460
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13906 7392 13912 7404
rect 13679 7364 13912 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 14642 7392 14648 7404
rect 14056 7364 14648 7392
rect 14056 7352 14062 7364
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 13446 7284 13452 7336
rect 13504 7284 13510 7336
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 14752 7324 14780 7420
rect 18156 7401 18184 7432
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18408 7395 18466 7401
rect 18408 7361 18420 7395
rect 18454 7392 18466 7395
rect 18782 7392 18788 7404
rect 18454 7364 18788 7392
rect 18454 7361 18466 7364
rect 18408 7355 18466 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 14424 7296 14780 7324
rect 19306 7336 19334 7432
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7392 19947 7395
rect 20254 7392 20260 7404
rect 19935 7364 20260 7392
rect 19935 7361 19947 7364
rect 19889 7355 19947 7361
rect 20254 7352 20260 7364
rect 20312 7352 20318 7404
rect 20438 7401 20444 7404
rect 20432 7392 20444 7401
rect 20399 7364 20444 7392
rect 20432 7355 20444 7364
rect 20438 7352 20444 7355
rect 20496 7352 20502 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 22020 7401 22048 7500
rect 22554 7488 22560 7540
rect 22612 7488 22618 7540
rect 23293 7531 23351 7537
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 23474 7528 23480 7540
rect 23339 7500 23480 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 24121 7531 24179 7537
rect 24121 7497 24133 7531
rect 24167 7528 24179 7531
rect 25130 7528 25136 7540
rect 24167 7500 25136 7528
rect 24167 7497 24179 7500
rect 24121 7491 24179 7497
rect 25130 7488 25136 7500
rect 25188 7488 25194 7540
rect 22572 7460 22600 7488
rect 22572 7432 23520 7460
rect 22005 7395 22063 7401
rect 20772 7364 21220 7392
rect 20772 7352 20778 7364
rect 19306 7296 19340 7336
rect 14424 7284 14430 7296
rect 19334 7284 19340 7296
rect 19392 7324 19398 7336
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 19392 7296 20177 7324
rect 19392 7284 19398 7296
rect 20165 7293 20177 7296
rect 20211 7293 20223 7327
rect 21192 7324 21220 7364
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22555 7395 22613 7401
rect 22555 7361 22567 7395
rect 22601 7392 22613 7395
rect 22646 7392 22652 7404
rect 22601 7364 22652 7392
rect 22601 7361 22613 7364
rect 22555 7355 22613 7361
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 22186 7324 22192 7336
rect 21192 7296 22192 7324
rect 20165 7287 20223 7293
rect 22186 7284 22192 7296
rect 22244 7324 22250 7336
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 22244 7296 22293 7324
rect 22244 7284 22250 7296
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 14553 7259 14611 7265
rect 12544 7228 13308 7256
rect 13280 7200 13308 7228
rect 14553 7225 14565 7259
rect 14599 7256 14611 7259
rect 16298 7256 16304 7268
rect 14599 7228 16304 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 16298 7216 16304 7228
rect 16356 7216 16362 7268
rect 21266 7256 21272 7268
rect 21100 7228 21272 7256
rect 9272 7160 10088 7188
rect 9272 7148 9278 7160
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10376 7160 10425 7188
rect 10376 7148 10382 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 10413 7151 10471 7157
rect 13262 7148 13268 7200
rect 13320 7148 13326 7200
rect 14458 7148 14464 7200
rect 14516 7188 14522 7200
rect 21100 7188 21128 7228
rect 21266 7216 21272 7228
rect 21324 7216 21330 7268
rect 23492 7256 23520 7432
rect 23750 7420 23756 7472
rect 23808 7420 23814 7472
rect 23845 7463 23903 7469
rect 23845 7429 23857 7463
rect 23891 7460 23903 7463
rect 24302 7460 24308 7472
rect 23891 7432 24308 7460
rect 23891 7429 23903 7432
rect 23845 7423 23903 7429
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 23768 7392 23796 7420
rect 24210 7392 24216 7404
rect 23768 7364 24216 7392
rect 24210 7352 24216 7364
rect 24268 7392 24274 7404
rect 24489 7395 24547 7401
rect 24489 7392 24501 7395
rect 24268 7364 24501 7392
rect 24268 7352 24274 7364
rect 24489 7361 24501 7364
rect 24535 7361 24547 7395
rect 24489 7355 24547 7361
rect 24305 7259 24363 7265
rect 24305 7256 24317 7259
rect 23492 7228 24317 7256
rect 24305 7225 24317 7228
rect 24351 7225 24363 7259
rect 24305 7219 24363 7225
rect 14516 7160 21128 7188
rect 14516 7148 14522 7160
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21232 7160 21833 7188
rect 21232 7148 21238 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 21821 7151 21879 7157
rect 1104 7098 24840 7120
rect 1104 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 9851 7098
rect 9903 7046 9915 7098
rect 9967 7046 9979 7098
rect 10031 7046 10043 7098
rect 10095 7046 10107 7098
rect 10159 7046 15785 7098
rect 15837 7046 15849 7098
rect 15901 7046 15913 7098
rect 15965 7046 15977 7098
rect 16029 7046 16041 7098
rect 16093 7046 21719 7098
rect 21771 7046 21783 7098
rect 21835 7046 21847 7098
rect 21899 7046 21911 7098
rect 21963 7046 21975 7098
rect 22027 7046 24840 7098
rect 1104 7024 24840 7046
rect 1578 6944 1584 6996
rect 1636 6944 1642 6996
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3602 6984 3608 6996
rect 3375 6956 3608 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 3988 6956 5488 6984
rect 2314 6808 2320 6860
rect 2372 6808 2378 6860
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6749 2283 6783
rect 2225 6743 2283 6749
rect 2591 6783 2649 6789
rect 2591 6749 2603 6783
rect 2637 6780 2649 6783
rect 3326 6780 3332 6792
rect 2637 6752 3332 6780
rect 2637 6749 2649 6752
rect 2591 6743 2649 6749
rect 1489 6715 1547 6721
rect 1489 6681 1501 6715
rect 1535 6712 1547 6715
rect 2240 6712 2268 6743
rect 3326 6740 3332 6752
rect 3384 6780 3390 6792
rect 3602 6780 3608 6792
rect 3384 6752 3608 6780
rect 3384 6740 3390 6752
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 3988 6789 4016 6956
rect 4338 6916 4344 6928
rect 4080 6888 4344 6916
rect 4080 6792 4108 6888
rect 4338 6876 4344 6888
rect 4396 6916 4402 6928
rect 4396 6888 4568 6916
rect 4396 6876 4402 6888
rect 4540 6857 4568 6888
rect 4525 6851 4583 6857
rect 4172 6820 4476 6848
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4062 6740 4068 6792
rect 4120 6740 4126 6792
rect 4172 6712 4200 6820
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 1535 6684 2084 6712
rect 2240 6684 4200 6712
rect 1535 6681 1547 6684
rect 1489 6675 1547 6681
rect 2056 6653 2084 6684
rect 2041 6647 2099 6653
rect 2041 6613 2053 6647
rect 2087 6613 2099 6647
rect 2041 6607 2099 6613
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3418 6644 3424 6656
rect 2832 6616 3424 6644
rect 2832 6604 2838 6616
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3752 6616 3801 6644
rect 3752 6604 3758 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3936 6616 4077 6644
rect 3936 6604 3942 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4264 6644 4292 6743
rect 4448 6712 4476 6820
rect 4525 6817 4537 6851
rect 4571 6817 4583 6851
rect 5460 6848 5488 6956
rect 5534 6944 5540 6996
rect 5592 6944 5598 6996
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 7834 6984 7840 6996
rect 6696 6956 7840 6984
rect 6696 6944 6702 6956
rect 7834 6944 7840 6956
rect 7892 6944 7898 6996
rect 9692 6956 13216 6984
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9585 6919 9643 6925
rect 9585 6916 9597 6919
rect 9088 6888 9597 6916
rect 9088 6876 9094 6888
rect 9585 6885 9597 6888
rect 9631 6885 9643 6919
rect 9585 6879 9643 6885
rect 8662 6848 8668 6860
rect 5460 6820 8668 6848
rect 4525 6811 4583 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 9692 6848 9720 6956
rect 13188 6916 13216 6956
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13504 6956 13553 6984
rect 13504 6944 13510 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 18598 6944 18604 6996
rect 18656 6944 18662 6996
rect 19610 6984 19616 6996
rect 19444 6956 19616 6984
rect 15470 6916 15476 6928
rect 13188 6888 15476 6916
rect 15470 6876 15476 6888
rect 15528 6876 15534 6928
rect 17788 6916 17816 6944
rect 19444 6916 19472 6956
rect 19610 6944 19616 6956
rect 19668 6944 19674 6996
rect 20254 6944 20260 6996
rect 20312 6984 20318 6996
rect 20717 6987 20775 6993
rect 20717 6984 20729 6987
rect 20312 6956 20729 6984
rect 20312 6944 20318 6956
rect 20717 6953 20729 6956
rect 20763 6953 20775 6987
rect 20717 6947 20775 6953
rect 21082 6944 21088 6996
rect 21140 6944 21146 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 21324 6956 22692 6984
rect 21324 6944 21330 6956
rect 17788 6888 19472 6916
rect 20346 6876 20352 6928
rect 20404 6876 20410 6928
rect 20530 6876 20536 6928
rect 20588 6916 20594 6928
rect 21729 6919 21787 6925
rect 21729 6916 21741 6919
rect 20588 6888 21741 6916
rect 20588 6876 20594 6888
rect 21729 6885 21741 6888
rect 21775 6885 21787 6919
rect 22370 6916 22376 6928
rect 21729 6879 21787 6885
rect 22112 6888 22376 6916
rect 8996 6820 9720 6848
rect 10137 6851 10195 6857
rect 8996 6808 9002 6820
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10318 6848 10324 6860
rect 10183 6820 10324 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 17862 6848 17868 6860
rect 15436 6820 17868 6848
rect 15436 6808 15442 6820
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 20364 6848 20392 6876
rect 21361 6851 21419 6857
rect 20364 6820 21036 6848
rect 4799 6783 4857 6789
rect 4799 6749 4811 6783
rect 4845 6780 4857 6783
rect 5810 6780 5816 6792
rect 4845 6752 5816 6780
rect 4845 6749 4857 6752
rect 4799 6743 4857 6749
rect 5810 6740 5816 6752
rect 5868 6740 5874 6792
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9306 6780 9312 6792
rect 9171 6752 9312 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 9950 6740 9956 6792
rect 10008 6789 10014 6792
rect 10008 6783 10036 6789
rect 10024 6749 10036 6783
rect 10008 6743 10036 6749
rect 10008 6740 10014 6743
rect 11698 6740 11704 6792
rect 11756 6780 11762 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 11756 6752 12541 6780
rect 11756 6740 11762 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12787 6753 12845 6759
rect 12787 6750 12799 6753
rect 12529 6743 12587 6749
rect 9030 6712 9036 6724
rect 4448 6684 9036 6712
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 12728 6722 12799 6750
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 4264 6616 10793 6644
rect 4065 6607 4123 6613
rect 10781 6613 10793 6616
rect 10827 6613 10839 6647
rect 12728 6644 12756 6722
rect 12787 6719 12799 6722
rect 12833 6719 12845 6753
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 17770 6780 17776 6792
rect 15528 6752 17776 6780
rect 15528 6740 15534 6752
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 19337 6783 19395 6789
rect 18840 6752 19196 6780
rect 18840 6740 18846 6752
rect 12787 6713 12845 6719
rect 19168 6656 19196 6752
rect 19337 6749 19349 6783
rect 19383 6749 19395 6783
rect 19337 6743 19395 6749
rect 19352 6712 19380 6743
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 19668 6752 19711 6780
rect 19668 6740 19674 6752
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 21008 6789 21036 6820
rect 21361 6817 21373 6851
rect 21407 6848 21419 6851
rect 22112 6848 22140 6888
rect 22370 6876 22376 6888
rect 22428 6876 22434 6928
rect 22664 6925 22692 6956
rect 23474 6944 23480 6996
rect 23532 6944 23538 6996
rect 22649 6919 22707 6925
rect 22649 6885 22661 6919
rect 22695 6885 22707 6919
rect 22649 6879 22707 6885
rect 22922 6876 22928 6928
rect 22980 6916 22986 6928
rect 23198 6916 23204 6928
rect 22980 6888 23204 6916
rect 22980 6876 22986 6888
rect 23198 6876 23204 6888
rect 23256 6876 23262 6928
rect 23290 6848 23296 6860
rect 21407 6820 22140 6848
rect 22204 6820 23296 6848
rect 21407 6817 21419 6820
rect 21361 6811 21419 6817
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20496 6752 20913 6780
rect 20496 6740 20502 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 20714 6712 20720 6724
rect 19352 6684 20720 6712
rect 20714 6672 20720 6684
rect 20772 6672 20778 6724
rect 13170 6644 13176 6656
rect 12728 6616 13176 6644
rect 10781 6607 10839 6613
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 15102 6604 15108 6656
rect 15160 6644 15166 6656
rect 17218 6644 17224 6656
rect 15160 6616 17224 6644
rect 15160 6604 15166 6616
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 19150 6604 19156 6656
rect 19208 6604 19214 6656
rect 20916 6644 20944 6743
rect 21174 6740 21180 6792
rect 21232 6740 21238 6792
rect 21266 6740 21272 6792
rect 21324 6740 21330 6792
rect 21542 6740 21548 6792
rect 21600 6740 21606 6792
rect 22204 6790 22232 6820
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 23492 6848 23520 6944
rect 23492 6820 23980 6848
rect 22005 6783 22063 6789
rect 22005 6749 22017 6783
rect 22051 6780 22063 6783
rect 22112 6780 22232 6790
rect 22051 6762 22232 6780
rect 22373 6783 22431 6789
rect 22051 6752 22140 6762
rect 22051 6749 22063 6752
rect 22005 6743 22063 6749
rect 22373 6749 22385 6783
rect 22419 6749 22431 6783
rect 22373 6743 22431 6749
rect 21082 6672 21088 6724
rect 21140 6712 21146 6724
rect 22388 6712 22416 6743
rect 22738 6740 22744 6792
rect 22796 6740 22802 6792
rect 23382 6740 23388 6792
rect 23440 6740 23446 6792
rect 23474 6740 23480 6792
rect 23532 6740 23538 6792
rect 23952 6789 23980 6820
rect 24026 6808 24032 6860
rect 24084 6808 24090 6860
rect 23937 6783 23995 6789
rect 23937 6749 23949 6783
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 24121 6783 24179 6789
rect 24121 6749 24133 6783
rect 24167 6749 24179 6783
rect 24121 6743 24179 6749
rect 24136 6712 24164 6743
rect 21140 6684 22416 6712
rect 22480 6684 24164 6712
rect 21140 6672 21146 6684
rect 21910 6644 21916 6656
rect 20916 6616 21916 6644
rect 21910 6604 21916 6616
rect 21968 6604 21974 6656
rect 22094 6604 22100 6656
rect 22152 6644 22158 6656
rect 22480 6644 22508 6684
rect 22152 6616 22508 6644
rect 22152 6604 22158 6616
rect 22554 6604 22560 6656
rect 22612 6644 22618 6656
rect 23201 6647 23259 6653
rect 23201 6644 23213 6647
rect 22612 6616 23213 6644
rect 22612 6604 22618 6616
rect 23201 6613 23213 6616
rect 23247 6613 23259 6647
rect 23201 6607 23259 6613
rect 23566 6604 23572 6656
rect 23624 6604 23630 6656
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 1360 6412 3433 6440
rect 1360 6400 1366 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3421 6403 3479 6409
rect 4982 6400 4988 6452
rect 5040 6400 5046 6452
rect 5626 6400 5632 6452
rect 5684 6400 5690 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 5776 6412 8309 6440
rect 5776 6400 5782 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 8938 6440 8944 6452
rect 8297 6403 8355 6409
rect 8864 6412 8944 6440
rect 1210 6332 1216 6384
rect 1268 6372 1274 6384
rect 2225 6375 2283 6381
rect 1268 6344 1808 6372
rect 1268 6332 1274 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1780 6304 1808 6344
rect 2225 6341 2237 6375
rect 2271 6372 2283 6375
rect 2958 6372 2964 6384
rect 2271 6344 2964 6372
rect 2271 6341 2283 6344
rect 2225 6335 2283 6341
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3329 6375 3387 6381
rect 3329 6341 3341 6375
rect 3375 6372 3387 6375
rect 5442 6372 5448 6384
rect 3375 6344 5448 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 1780 6276 2605 6304
rect 1673 6267 1731 6273
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 2593 6267 2651 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 4247 6307 4305 6313
rect 2823 6276 3280 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 1688 6236 1716 6267
rect 3142 6236 3148 6248
rect 1688 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 1302 6128 1308 6180
rect 1360 6168 1366 6180
rect 3252 6168 3280 6276
rect 4247 6273 4259 6307
rect 4293 6304 4305 6307
rect 4706 6304 4712 6316
rect 4293 6276 4712 6304
rect 4293 6273 4305 6276
rect 4247 6267 4305 6273
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5644 6304 5672 6400
rect 5583 6276 5672 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6328 6276 6377 6304
rect 6328 6264 6334 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6512 6276 6561 6304
rect 6512 6264 6518 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7374 6264 7380 6316
rect 7432 6313 7438 6316
rect 7432 6307 7460 6313
rect 7448 6273 7460 6307
rect 7432 6267 7460 6273
rect 7432 6264 7438 6267
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 8864 6313 8892 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 9088 6412 10701 6440
rect 9088 6400 9094 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 12526 6440 12532 6452
rect 10689 6403 10747 6409
rect 11716 6412 12532 6440
rect 9950 6313 9956 6316
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8251 6276 8493 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 9907 6307 9956 6313
rect 9907 6273 9919 6307
rect 9953 6273 9956 6307
rect 9907 6267 9956 6273
rect 9950 6264 9956 6267
rect 10008 6264 10014 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11606 6304 11612 6316
rect 11563 6276 11612 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3970 6236 3976 6248
rect 3660 6208 3976 6236
rect 3660 6196 3666 6208
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 8110 6236 8116 6248
rect 7331 6208 8116 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 9398 6236 9404 6248
rect 9079 6208 9404 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9398 6196 9404 6208
rect 9456 6196 9462 6248
rect 9766 6196 9772 6248
rect 9824 6196 9830 6248
rect 10045 6239 10103 6245
rect 10045 6205 10057 6239
rect 10091 6236 10103 6239
rect 10226 6236 10232 6248
rect 10091 6208 10232 6236
rect 10091 6205 10103 6208
rect 10045 6199 10103 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 11716 6245 11744 6412
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 13320 6412 13860 6440
rect 13320 6400 13326 6412
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 10520 6208 11713 6236
rect 3786 6168 3792 6180
rect 1360 6140 2774 6168
rect 3252 6140 3792 6168
rect 1360 6128 1366 6140
rect 1762 6060 1768 6112
rect 1820 6060 1826 6112
rect 2746 6100 2774 6140
rect 3786 6128 3792 6140
rect 3844 6128 3850 6180
rect 7009 6171 7067 6177
rect 7009 6137 7021 6171
rect 7055 6137 7067 6171
rect 7009 6131 7067 6137
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2746 6072 2881 6100
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 2869 6063 2927 6069
rect 5350 6060 5356 6112
rect 5408 6060 5414 6112
rect 7024 6100 7052 6131
rect 7374 6100 7380 6112
rect 7024 6072 7380 6100
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 8128 6100 8156 6196
rect 10520 6180 10548 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 12434 6207 12440 6259
rect 12492 6207 12498 6259
rect 12575 6239 12633 6245
rect 11701 6199 11759 6205
rect 12437 6205 12449 6207
rect 12483 6205 12495 6207
rect 12437 6199 12495 6205
rect 12575 6205 12587 6239
rect 12621 6236 12633 6239
rect 13280 6236 13308 6400
rect 13832 6372 13860 6412
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 13964 6412 14473 6440
rect 13964 6400 13970 6412
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 15470 6400 15476 6452
rect 15528 6440 15534 6452
rect 16758 6440 16764 6452
rect 15528 6412 16764 6440
rect 15528 6400 15534 6412
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 17678 6440 17684 6452
rect 16868 6412 17684 6440
rect 16868 6372 16896 6412
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 17920 6412 17969 6440
rect 17920 6400 17926 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 19058 6440 19064 6452
rect 18288 6412 19064 6440
rect 18288 6400 18294 6412
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6440 19855 6443
rect 21082 6440 21088 6452
rect 19843 6412 21088 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 21082 6400 21088 6412
rect 21140 6440 21146 6452
rect 21140 6412 21312 6440
rect 21140 6400 21146 6412
rect 13832 6344 16896 6372
rect 13707 6337 13765 6343
rect 13707 6303 13719 6337
rect 13753 6334 13765 6337
rect 13753 6316 13768 6334
rect 17494 6332 17500 6384
rect 17552 6372 17558 6384
rect 19886 6372 19892 6384
rect 17552 6344 19892 6372
rect 17552 6332 17558 6344
rect 19886 6332 19892 6344
rect 19944 6332 19950 6384
rect 20622 6372 20628 6384
rect 19996 6344 20628 6372
rect 13707 6297 13728 6303
rect 13722 6264 13728 6297
rect 13780 6264 13786 6316
rect 14921 6307 14979 6313
rect 14921 6273 14933 6307
rect 14967 6304 14979 6307
rect 15102 6304 15108 6316
rect 14967 6276 15108 6304
rect 14967 6273 14979 6276
rect 14921 6267 14979 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15194 6264 15200 6316
rect 15252 6304 15258 6316
rect 16390 6304 16396 6316
rect 15252 6276 16396 6304
rect 15252 6264 15258 6276
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 18230 6304 18236 6316
rect 17727 6276 18236 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 19996 6313 20024 6344
rect 20622 6332 20628 6344
rect 20680 6332 20686 6384
rect 21284 6372 21312 6412
rect 22048 6400 22054 6452
rect 22106 6400 22112 6452
rect 22738 6400 22744 6452
rect 22796 6440 22802 6452
rect 23293 6443 23351 6449
rect 23293 6440 23305 6443
rect 22796 6412 23305 6440
rect 22796 6400 22802 6412
rect 23293 6409 23305 6412
rect 23339 6409 23351 6443
rect 23293 6403 23351 6409
rect 23937 6443 23995 6449
rect 23937 6409 23949 6443
rect 23983 6409 23995 6443
rect 23937 6403 23995 6409
rect 22066 6372 22094 6400
rect 23952 6372 23980 6403
rect 24210 6400 24216 6452
rect 24268 6440 24274 6452
rect 24305 6443 24363 6449
rect 24305 6440 24317 6443
rect 24268 6412 24317 6440
rect 24268 6400 24274 6412
rect 24305 6409 24317 6412
rect 24351 6409 24363 6443
rect 24305 6403 24363 6409
rect 21284 6344 21680 6372
rect 22066 6344 23980 6372
rect 19981 6307 20039 6313
rect 19981 6273 19993 6307
rect 20027 6273 20039 6307
rect 19981 6267 20039 6273
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6304 20407 6307
rect 20530 6304 20536 6316
rect 20395 6276 20536 6304
rect 20395 6273 20407 6276
rect 20349 6267 20407 6273
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 21652 6313 21680 6344
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20732 6276 20821 6304
rect 12621 6208 13308 6236
rect 13449 6239 13507 6245
rect 12621 6205 12633 6208
rect 12575 6199 12633 6205
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6236 18015 6239
rect 18414 6236 18420 6248
rect 18003 6208 18420 6236
rect 18003 6205 18015 6208
rect 17957 6199 18015 6205
rect 9490 6128 9496 6180
rect 9548 6128 9554 6180
rect 10502 6128 10508 6180
rect 10560 6128 10566 6180
rect 12158 6128 12164 6180
rect 12216 6128 12222 6180
rect 13354 6128 13360 6180
rect 13412 6128 13418 6180
rect 11054 6100 11060 6112
rect 8128 6072 11060 6100
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 13464 6100 13492 6199
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 20732 6180 20760 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21177 6308 21235 6313
rect 21177 6307 21312 6308
rect 20947 6276 21131 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21103 6236 21131 6276
rect 21177 6273 21189 6307
rect 21223 6304 21312 6307
rect 21637 6307 21695 6313
rect 21223 6280 21496 6304
rect 21223 6273 21235 6280
rect 21284 6276 21496 6280
rect 21177 6267 21235 6273
rect 21266 6236 21272 6248
rect 21103 6208 21272 6236
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 17773 6171 17831 6177
rect 17773 6137 17785 6171
rect 17819 6168 17831 6171
rect 18138 6168 18144 6180
rect 17819 6140 18144 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 20162 6128 20168 6180
rect 20220 6168 20226 6180
rect 20533 6171 20591 6177
rect 20533 6168 20545 6171
rect 20220 6140 20545 6168
rect 20220 6128 20226 6140
rect 20533 6137 20545 6140
rect 20579 6137 20591 6171
rect 20533 6131 20591 6137
rect 20622 6128 20628 6180
rect 20680 6128 20686 6180
rect 20714 6128 20720 6180
rect 20772 6128 20778 6180
rect 21174 6128 21180 6180
rect 21232 6128 21238 6180
rect 21468 6177 21496 6276
rect 21637 6273 21649 6307
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 21818 6264 21824 6316
rect 21876 6264 21882 6316
rect 22063 6307 22121 6313
rect 22063 6273 22075 6307
rect 22109 6304 22121 6307
rect 22646 6304 22652 6316
rect 22109 6302 22140 6304
rect 22296 6302 22652 6304
rect 22109 6276 22652 6302
rect 22109 6274 22324 6276
rect 22109 6273 22121 6274
rect 22063 6267 22121 6273
rect 22646 6264 22652 6276
rect 22704 6264 22710 6316
rect 23201 6307 23259 6313
rect 23201 6273 23213 6307
rect 23247 6304 23259 6307
rect 23290 6304 23296 6316
rect 23247 6276 23296 6304
rect 23247 6273 23259 6276
rect 23201 6267 23259 6273
rect 21453 6171 21511 6177
rect 21453 6137 21465 6171
rect 21499 6137 21511 6171
rect 21453 6131 21511 6137
rect 22833 6171 22891 6177
rect 22833 6137 22845 6171
rect 22879 6168 22891 6171
rect 23216 6168 23244 6267
rect 23290 6264 23296 6276
rect 23348 6264 23354 6316
rect 23385 6307 23443 6313
rect 23385 6273 23397 6307
rect 23431 6273 23443 6307
rect 23385 6267 23443 6273
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6273 23719 6307
rect 23661 6267 23719 6273
rect 22879 6140 23244 6168
rect 22879 6137 22891 6140
rect 22833 6131 22891 6137
rect 11756 6072 13492 6100
rect 15933 6103 15991 6109
rect 11756 6060 11762 6072
rect 15933 6069 15945 6103
rect 15979 6100 15991 6103
rect 16298 6100 16304 6112
rect 15979 6072 16304 6100
rect 15979 6069 15991 6072
rect 15933 6063 15991 6069
rect 16298 6060 16304 6072
rect 16356 6060 16362 6112
rect 20070 6060 20076 6112
rect 20128 6060 20134 6112
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 21085 6103 21143 6109
rect 21085 6100 21097 6103
rect 20956 6072 21097 6100
rect 20956 6060 20962 6072
rect 21085 6069 21097 6072
rect 21131 6069 21143 6103
rect 21192 6100 21220 6128
rect 21269 6103 21327 6109
rect 21269 6100 21281 6103
rect 21192 6072 21281 6100
rect 21085 6063 21143 6069
rect 21269 6069 21281 6072
rect 21315 6069 21327 6103
rect 21269 6063 21327 6069
rect 21542 6060 21548 6112
rect 21600 6100 21606 6112
rect 23400 6100 23428 6267
rect 23676 6236 23704 6267
rect 23750 6264 23756 6316
rect 23808 6264 23814 6316
rect 24026 6264 24032 6316
rect 24084 6264 24090 6316
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 24210 6236 24216 6248
rect 23676 6208 24216 6236
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 21600 6072 23428 6100
rect 21600 6060 21606 6072
rect 23474 6060 23480 6112
rect 23532 6060 23538 6112
rect 24118 6060 24124 6112
rect 24176 6060 24182 6112
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1452 5868 1593 5896
rect 1452 5856 1458 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 2130 5856 2136 5908
rect 2188 5856 2194 5908
rect 3237 5899 3295 5905
rect 3237 5896 3249 5899
rect 2746 5868 3249 5896
rect 1026 5788 1032 5840
rect 1084 5828 1090 5840
rect 2746 5828 2774 5868
rect 3237 5865 3249 5868
rect 3283 5865 3295 5899
rect 3237 5859 3295 5865
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 5350 5896 5356 5908
rect 3936 5868 5356 5896
rect 3936 5856 3942 5868
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 5500 5868 5641 5896
rect 5500 5856 5506 5868
rect 5629 5865 5641 5868
rect 5675 5865 5687 5899
rect 5629 5859 5687 5865
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 7101 5899 7159 5905
rect 6144 5868 6774 5896
rect 6144 5856 6150 5868
rect 1084 5800 2774 5828
rect 4724 5800 6132 5828
rect 1084 5788 1090 5800
rect 4724 5772 4752 5800
rect 3050 5720 3056 5772
rect 3108 5760 3114 5772
rect 3970 5760 3976 5772
rect 3108 5732 3976 5760
rect 3108 5720 3114 5732
rect 3970 5720 3976 5732
rect 4028 5720 4034 5772
rect 4706 5720 4712 5772
rect 4764 5720 4770 5772
rect 5902 5760 5908 5772
rect 5552 5732 5908 5760
rect 2593 5695 2651 5701
rect 1504 5664 2176 5692
rect 1504 5633 1532 5664
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5593 1547 5627
rect 1489 5587 1547 5593
rect 2038 5584 2044 5636
rect 2096 5584 2102 5636
rect 2148 5624 2176 5664
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3145 5695 3203 5701
rect 2639 5664 3096 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3068 5624 3096 5664
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3878 5692 3884 5704
rect 3191 5664 3884 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 4247 5695 4305 5701
rect 4247 5661 4259 5695
rect 4293 5692 4305 5695
rect 5258 5692 5264 5704
rect 4293 5664 5264 5692
rect 4293 5661 4305 5664
rect 4247 5655 4305 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5552 5701 5580 5732
rect 5902 5720 5908 5732
rect 5960 5720 5966 5772
rect 6104 5769 6132 5800
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5729 6147 5763
rect 6746 5760 6774 5868
rect 7101 5865 7113 5899
rect 7147 5896 7159 5899
rect 7558 5896 7564 5908
rect 7147 5868 7564 5896
rect 7147 5865 7159 5868
rect 7101 5859 7159 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 9490 5896 9496 5908
rect 8527 5868 9496 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 10594 5896 10600 5908
rect 9600 5868 10600 5896
rect 7469 5763 7527 5769
rect 7469 5760 7481 5763
rect 6746 5732 7481 5760
rect 6089 5723 6147 5729
rect 7469 5729 7481 5732
rect 7515 5729 7527 5763
rect 7469 5723 7527 5729
rect 5537 5695 5595 5701
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 2148 5596 3004 5624
rect 3068 5596 5396 5624
rect 2866 5516 2872 5568
rect 2924 5516 2930 5568
rect 2976 5556 3004 5596
rect 4338 5556 4344 5568
rect 2976 5528 4344 5556
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4982 5516 4988 5568
rect 5040 5516 5046 5568
rect 5368 5565 5396 5596
rect 5353 5559 5411 5565
rect 5353 5525 5365 5559
rect 5399 5525 5411 5559
rect 6104 5556 6132 5723
rect 6347 5665 6405 5671
rect 6347 5631 6359 5665
rect 6393 5662 6405 5665
rect 6393 5631 6406 5662
rect 6347 5625 6406 5631
rect 6378 5624 6406 5625
rect 6638 5624 6644 5636
rect 6378 5596 6644 5624
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 7484 5624 7512 5723
rect 7743 5695 7801 5701
rect 7743 5661 7755 5695
rect 7789 5692 7801 5695
rect 9600 5692 9628 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 12158 5896 12164 5908
rect 10919 5868 12164 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 14458 5896 14464 5908
rect 12492 5868 14464 5896
rect 12492 5856 12498 5868
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 14918 5896 14924 5908
rect 14792 5868 14924 5896
rect 14792 5856 14798 5868
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15378 5856 15384 5908
rect 15436 5856 15442 5908
rect 16298 5896 16304 5908
rect 15948 5868 16304 5896
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 12084 5800 12265 5828
rect 9674 5720 9680 5772
rect 9732 5760 9738 5772
rect 9732 5732 9904 5760
rect 9732 5720 9738 5732
rect 9876 5701 9904 5732
rect 7789 5664 9628 5692
rect 9861 5695 9919 5701
rect 7789 5661 7801 5664
rect 7743 5655 7801 5661
rect 9861 5661 9873 5695
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 7558 5624 7564 5636
rect 7484 5596 7564 5624
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 9876 5624 9904 5655
rect 10134 5652 10140 5704
rect 10192 5692 10198 5704
rect 10192 5664 10235 5692
rect 10192 5652 10198 5664
rect 11146 5652 11152 5704
rect 11204 5692 11210 5704
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 11204 5664 11253 5692
rect 11204 5652 11210 5664
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11515 5695 11573 5701
rect 11515 5692 11527 5695
rect 11241 5655 11299 5661
rect 11440 5664 11527 5692
rect 11440 5636 11468 5664
rect 11515 5661 11527 5664
rect 11561 5661 11573 5695
rect 12084 5692 12112 5800
rect 12253 5797 12265 5800
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 12710 5788 12716 5840
rect 12768 5788 12774 5840
rect 15396 5828 15424 5856
rect 15948 5837 15976 5868
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 16390 5856 16396 5908
rect 16448 5896 16454 5908
rect 16448 5868 17908 5896
rect 16448 5856 16454 5868
rect 15304 5800 15424 5828
rect 15933 5831 15991 5837
rect 12158 5720 12164 5772
rect 12216 5760 12222 5772
rect 12434 5760 12440 5772
rect 12216 5732 12440 5760
rect 12216 5720 12222 5732
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 12728 5692 12756 5788
rect 15304 5772 15332 5800
rect 15933 5797 15945 5831
rect 15979 5797 15991 5831
rect 15933 5791 15991 5797
rect 15286 5720 15292 5772
rect 15344 5720 15350 5772
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 16209 5763 16267 5769
rect 16209 5760 16221 5763
rect 15436 5732 16221 5760
rect 15436 5720 15442 5732
rect 16209 5729 16221 5732
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 16298 5720 16304 5772
rect 16356 5769 16362 5772
rect 16356 5763 16384 5769
rect 16372 5729 16384 5763
rect 16356 5723 16384 5729
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 17126 5760 17132 5772
rect 16531 5732 17132 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16356 5720 16362 5723
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 12084 5664 12756 5692
rect 11515 5655 11573 5661
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 15470 5692 15476 5704
rect 14976 5664 15476 5692
rect 14976 5652 14982 5664
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5661 17279 5695
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17221 5655 17279 5661
rect 9950 5624 9956 5636
rect 9876 5596 9956 5624
rect 9950 5584 9956 5596
rect 10008 5584 10014 5636
rect 11422 5584 11428 5636
rect 11480 5584 11486 5636
rect 15378 5624 15384 5636
rect 15120 5596 15384 5624
rect 6362 5556 6368 5568
rect 6104 5528 6368 5556
rect 5353 5519 5411 5525
rect 6362 5516 6368 5528
rect 6420 5556 6426 5568
rect 8018 5556 8024 5568
rect 6420 5528 8024 5556
rect 6420 5516 6426 5528
rect 8018 5516 8024 5528
rect 8076 5516 8082 5568
rect 9674 5516 9680 5568
rect 9732 5556 9738 5568
rect 10134 5556 10140 5568
rect 9732 5528 10140 5556
rect 9732 5516 9738 5528
rect 10134 5516 10140 5528
rect 10192 5556 10198 5568
rect 10962 5556 10968 5568
rect 10192 5528 10968 5556
rect 10192 5516 10198 5528
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 15120 5556 15148 5596
rect 15378 5584 15384 5596
rect 15436 5584 15442 5636
rect 11112 5528 15148 5556
rect 11112 5516 11118 5528
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 17129 5559 17187 5565
rect 17129 5556 17141 5559
rect 15252 5528 17141 5556
rect 15252 5516 15258 5528
rect 17129 5525 17141 5528
rect 17175 5525 17187 5559
rect 17236 5556 17264 5655
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17880 5624 17908 5868
rect 18230 5856 18236 5908
rect 18288 5856 18294 5908
rect 19150 5856 19156 5908
rect 19208 5896 19214 5908
rect 19208 5868 19923 5896
rect 19208 5856 19214 5868
rect 19895 5828 19923 5868
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 22925 5899 22983 5905
rect 22925 5896 22937 5899
rect 20772 5868 22937 5896
rect 20772 5856 20778 5868
rect 22925 5865 22937 5868
rect 22971 5865 22983 5899
rect 22925 5859 22983 5865
rect 23290 5856 23296 5908
rect 23348 5896 23354 5908
rect 23566 5896 23572 5908
rect 23348 5868 23572 5896
rect 23348 5856 23354 5868
rect 23566 5856 23572 5868
rect 23624 5856 23630 5908
rect 24118 5856 24124 5908
rect 24176 5856 24182 5908
rect 20901 5831 20959 5837
rect 20901 5828 20913 5831
rect 19895 5800 20913 5828
rect 20901 5797 20913 5800
rect 20947 5797 20959 5831
rect 20901 5791 20959 5797
rect 21174 5788 21180 5840
rect 21232 5828 21238 5840
rect 21453 5831 21511 5837
rect 21453 5828 21465 5831
rect 21232 5800 21465 5828
rect 21232 5788 21238 5800
rect 21453 5797 21465 5800
rect 21499 5797 21511 5831
rect 21453 5791 21511 5797
rect 23198 5788 23204 5840
rect 23256 5828 23262 5840
rect 23937 5831 23995 5837
rect 23937 5828 23949 5831
rect 23256 5800 23949 5828
rect 23256 5788 23262 5800
rect 23937 5797 23949 5800
rect 23983 5797 23995 5831
rect 23937 5791 23995 5797
rect 19058 5720 19064 5772
rect 19116 5760 19122 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 19116 5732 19257 5760
rect 19116 5720 19122 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 24136 5760 24164 5856
rect 19245 5723 19303 5729
rect 21100 5732 21680 5760
rect 21100 5704 21128 5732
rect 19487 5695 19545 5701
rect 19487 5692 19499 5695
rect 19352 5664 19499 5692
rect 19352 5624 19380 5664
rect 19487 5661 19499 5664
rect 19533 5661 19545 5695
rect 19487 5655 19545 5661
rect 20714 5652 20720 5704
rect 20772 5652 20778 5704
rect 20990 5652 20996 5704
rect 21048 5652 21054 5704
rect 21082 5652 21088 5704
rect 21140 5652 21146 5704
rect 21269 5671 21327 5677
rect 21269 5637 21281 5671
rect 21315 5668 21327 5671
rect 21315 5640 21404 5668
rect 21542 5652 21548 5704
rect 21600 5652 21606 5704
rect 21315 5637 21327 5640
rect 21269 5631 21327 5637
rect 17880 5596 19380 5624
rect 21376 5624 21404 5640
rect 21652 5624 21680 5732
rect 23676 5732 24164 5760
rect 23293 5695 23351 5701
rect 23293 5661 23305 5695
rect 23339 5692 23351 5695
rect 23566 5692 23572 5704
rect 23339 5664 23572 5692
rect 23339 5661 23351 5664
rect 23293 5655 23351 5661
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 23676 5701 23704 5732
rect 23661 5695 23719 5701
rect 23661 5661 23673 5695
rect 23707 5661 23719 5695
rect 23661 5655 23719 5661
rect 23934 5652 23940 5704
rect 23992 5652 23998 5704
rect 21790 5627 21848 5633
rect 21790 5624 21802 5627
rect 21376 5596 21588 5624
rect 21652 5596 21802 5624
rect 19058 5556 19064 5568
rect 17236 5528 19064 5556
rect 17129 5519 17187 5525
rect 19058 5516 19064 5528
rect 19116 5556 19122 5568
rect 19242 5556 19248 5568
rect 19116 5528 19248 5556
rect 19116 5516 19122 5528
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 19576 5528 20269 5556
rect 19576 5516 19582 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 21177 5559 21235 5565
rect 21177 5525 21189 5559
rect 21223 5556 21235 5559
rect 21450 5556 21456 5568
rect 21223 5528 21456 5556
rect 21223 5525 21235 5528
rect 21177 5519 21235 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 21560 5556 21588 5596
rect 21790 5593 21802 5596
rect 21836 5593 21848 5627
rect 21790 5587 21848 5593
rect 23198 5556 23204 5568
rect 21560 5528 23204 5556
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 2958 5352 2964 5364
rect 1688 5324 2964 5352
rect 1688 5255 1716 5324
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3326 5352 3332 5364
rect 3108 5324 3332 5352
rect 3108 5312 3114 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 4706 5352 4712 5364
rect 4028 5324 4712 5352
rect 4028 5312 4034 5324
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5868 5324 6193 5352
rect 5868 5312 5874 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 6181 5315 6239 5321
rect 9506 5324 9718 5352
rect 3602 5284 3608 5296
rect 1655 5249 1716 5255
rect 1118 5176 1124 5228
rect 1176 5216 1182 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1176 5188 1409 5216
rect 1176 5176 1182 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1655 5215 1667 5249
rect 1701 5218 1716 5249
rect 2792 5256 3608 5284
rect 1701 5215 1713 5218
rect 1655 5209 1713 5215
rect 1397 5179 1455 5185
rect 1412 5012 1440 5179
rect 2792 5157 2820 5256
rect 3602 5244 3608 5256
rect 3660 5244 3666 5296
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 9214 5284 9220 5296
rect 6512 5256 9220 5284
rect 6512 5244 6518 5256
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 9506 5235 9534 5324
rect 9690 5284 9718 5324
rect 10226 5312 10232 5364
rect 10284 5312 10290 5364
rect 14366 5352 14372 5364
rect 12912 5324 14372 5352
rect 10870 5284 10876 5296
rect 9690 5256 10876 5284
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 9491 5229 9549 5235
rect 3051 5219 3109 5225
rect 3051 5185 3063 5219
rect 3097 5216 3109 5219
rect 3510 5216 3516 5228
rect 3097 5188 3516 5216
rect 3097 5185 3109 5188
rect 3051 5179 3109 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4430 5216 4436 5228
rect 4387 5188 4436 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4430 5176 4436 5188
rect 4488 5216 4494 5228
rect 4488 5188 4752 5216
rect 4488 5176 4494 5188
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 2332 5120 2789 5148
rect 1670 5012 1676 5024
rect 1412 4984 1676 5012
rect 1670 4972 1676 4984
rect 1728 5012 1734 5024
rect 2332 5012 2360 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 2777 5111 2835 5117
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4614 5148 4620 5160
rect 4571 5120 4620 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 4724 5148 4752 5188
rect 5350 5176 5356 5228
rect 5408 5225 5414 5228
rect 5408 5219 5436 5225
rect 5424 5185 5436 5219
rect 5408 5179 5436 5185
rect 5408 5176 5414 5179
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6639 5219 6697 5225
rect 6639 5185 6651 5219
rect 6685 5216 6697 5219
rect 7466 5216 7472 5228
rect 6685 5188 7472 5216
rect 6685 5185 6697 5188
rect 6639 5179 6697 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 7616 5188 9260 5216
rect 9491 5195 9503 5229
rect 9537 5195 9549 5229
rect 9491 5189 9549 5195
rect 7616 5176 7622 5188
rect 9232 5160 9260 5188
rect 12618 5176 12624 5228
rect 12676 5216 12682 5228
rect 12713 5219 12771 5225
rect 12713 5216 12725 5219
rect 12676 5188 12725 5216
rect 12676 5176 12682 5188
rect 12713 5185 12725 5188
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 4890 5148 4896 5160
rect 4724 5120 4896 5148
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 4982 5108 4988 5160
rect 5040 5108 5046 5160
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 5132 5120 5273 5148
rect 5132 5108 5138 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5534 5108 5540 5160
rect 5592 5108 5598 5160
rect 9214 5108 9220 5160
rect 9272 5108 9278 5160
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 12912 5157 12940 5324
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 15286 5352 15292 5364
rect 14660 5324 15292 5352
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5185 13691 5219
rect 13633 5179 13691 5185
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 10284 5120 12909 5148
rect 10284 5108 10290 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13078 5108 13084 5160
rect 13136 5148 13142 5160
rect 13648 5148 13676 5179
rect 13906 5176 13912 5228
rect 13964 5176 13970 5228
rect 14660 5225 14688 5324
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 16298 5352 16304 5364
rect 15804 5324 16304 5352
rect 15804 5312 15810 5324
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17681 5355 17739 5361
rect 17681 5352 17693 5355
rect 17184 5324 17693 5352
rect 17184 5312 17190 5324
rect 17681 5321 17693 5324
rect 17727 5321 17739 5355
rect 17681 5315 17739 5321
rect 18138 5312 18144 5364
rect 18196 5312 18202 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 18288 5324 18368 5352
rect 18288 5312 18294 5324
rect 17586 5284 17592 5296
rect 16958 5256 17592 5284
rect 15746 5225 15752 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 15703 5219 15752 5225
rect 15703 5185 15715 5219
rect 15749 5185 15752 5219
rect 15703 5179 15752 5185
rect 15746 5176 15752 5179
rect 15804 5176 15810 5228
rect 16958 5225 16986 5256
rect 17586 5244 17592 5256
rect 17644 5244 17650 5296
rect 16943 5219 17001 5225
rect 16943 5185 16955 5219
rect 16989 5185 17001 5219
rect 16943 5179 17001 5185
rect 13814 5157 13820 5160
rect 13136 5120 13676 5148
rect 13771 5151 13820 5157
rect 13136 5108 13142 5120
rect 13771 5117 13783 5151
rect 13817 5117 13820 5151
rect 13771 5111 13820 5117
rect 13814 5108 13820 5111
rect 13872 5108 13878 5160
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 14918 5148 14924 5160
rect 14875 5120 14924 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15436 5120 15577 5148
rect 15436 5108 15442 5120
rect 15565 5117 15577 5120
rect 15611 5117 15623 5151
rect 15565 5111 15623 5117
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16390 5148 16396 5160
rect 15887 5120 16396 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5117 16727 5151
rect 17604 5148 17632 5244
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18340 5225 18368 5324
rect 18414 5312 18420 5364
rect 18472 5312 18478 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 18524 5324 18613 5352
rect 18524 5225 18552 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 18601 5315 18659 5321
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 19886 5352 19892 5364
rect 18748 5324 19892 5352
rect 18748 5312 18754 5324
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 20070 5312 20076 5364
rect 20128 5352 20134 5364
rect 20128 5324 23336 5352
rect 20128 5312 20134 5324
rect 19518 5244 19524 5296
rect 19576 5244 19582 5296
rect 20162 5244 20168 5296
rect 20220 5284 20226 5296
rect 20220 5256 21496 5284
rect 20220 5244 20226 5256
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 18012 5188 18061 5216
rect 18012 5176 18018 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18049 5179 18107 5185
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 18782 5176 18788 5228
rect 18840 5176 18846 5228
rect 18966 5176 18972 5228
rect 19024 5216 19030 5228
rect 19153 5219 19211 5225
rect 19153 5216 19165 5219
rect 19024 5188 19165 5216
rect 19024 5176 19030 5188
rect 19153 5185 19165 5188
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 19337 5219 19395 5225
rect 19337 5185 19349 5219
rect 19383 5216 19395 5219
rect 19426 5216 19432 5228
rect 19383 5188 19432 5216
rect 19383 5185 19395 5188
rect 19337 5179 19395 5185
rect 19426 5176 19432 5188
rect 19484 5176 19490 5228
rect 19855 5219 19913 5225
rect 19855 5216 19867 5219
rect 19536 5188 19867 5216
rect 19536 5148 19564 5188
rect 19855 5185 19867 5188
rect 19901 5185 19913 5219
rect 19855 5179 19913 5185
rect 17604 5120 19564 5148
rect 19613 5151 19671 5157
rect 16669 5111 16727 5117
rect 19613 5117 19625 5151
rect 19659 5117 19671 5151
rect 20806 5148 20812 5160
rect 19613 5111 19671 5117
rect 20640 5120 20812 5148
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8294 5080 8300 5092
rect 7616 5052 8300 5080
rect 7616 5040 7622 5052
rect 8294 5040 8300 5052
rect 8352 5040 8358 5092
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 11146 5080 11152 5092
rect 10008 5052 11152 5080
rect 10008 5040 10014 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 13354 5040 13360 5092
rect 13412 5040 13418 5092
rect 14476 5052 14688 5080
rect 1728 4984 2360 5012
rect 2409 5015 2467 5021
rect 1728 4972 1734 4984
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 2498 5012 2504 5024
rect 2455 4984 2504 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 3602 4972 3608 5024
rect 3660 5012 3666 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3660 4984 3801 5012
rect 3660 4972 3666 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3789 4975 3847 4981
rect 7374 4972 7380 5024
rect 7432 4972 7438 5024
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 14476 5012 14504 5052
rect 8720 4984 14504 5012
rect 8720 4972 8726 4984
rect 14550 4972 14556 5024
rect 14608 4972 14614 5024
rect 14660 5012 14688 5052
rect 15286 5040 15292 5092
rect 15344 5040 15350 5092
rect 16298 5040 16304 5092
rect 16356 5080 16362 5092
rect 16684 5080 16712 5111
rect 16356 5052 16712 5080
rect 19153 5083 19211 5089
rect 16356 5040 16362 5052
rect 19153 5049 19165 5083
rect 19199 5049 19211 5083
rect 19153 5043 19211 5049
rect 16485 5015 16543 5021
rect 16485 5012 16497 5015
rect 14660 4984 16497 5012
rect 16485 4981 16497 4984
rect 16531 4981 16543 5015
rect 16485 4975 16543 4981
rect 17770 4972 17776 5024
rect 17828 5012 17834 5024
rect 19168 5012 19196 5043
rect 19242 5040 19248 5092
rect 19300 5080 19306 5092
rect 19628 5080 19656 5111
rect 20640 5089 20668 5120
rect 20806 5108 20812 5120
rect 20864 5148 20870 5160
rect 20916 5157 21036 5182
rect 21174 5176 21180 5228
rect 21232 5176 21238 5228
rect 21468 5225 21496 5256
rect 21453 5219 21511 5225
rect 21453 5185 21465 5219
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 21542 5176 21548 5228
rect 21600 5176 21606 5228
rect 22189 5219 22247 5225
rect 22189 5185 22201 5219
rect 22235 5216 22247 5219
rect 22278 5216 22284 5228
rect 22235 5188 22284 5216
rect 22235 5185 22247 5188
rect 22189 5179 22247 5185
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 23308 5216 23336 5324
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 24489 5355 24547 5361
rect 24489 5352 24501 5355
rect 24268 5324 24501 5352
rect 24268 5312 24274 5324
rect 24489 5321 24501 5324
rect 24535 5321 24547 5355
rect 24489 5315 24547 5321
rect 23376 5219 23434 5225
rect 23376 5216 23388 5219
rect 23308 5188 23388 5216
rect 23376 5185 23388 5188
rect 23422 5216 23434 5219
rect 24302 5216 24308 5228
rect 23422 5188 24308 5216
rect 23422 5185 23434 5188
rect 23376 5179 23434 5185
rect 24302 5176 24308 5188
rect 24360 5176 24366 5228
rect 20916 5154 21051 5157
rect 20916 5148 20944 5154
rect 20864 5120 20944 5148
rect 20993 5151 21051 5154
rect 20864 5108 20870 5120
rect 20993 5117 21005 5151
rect 21039 5117 21051 5151
rect 20993 5111 21051 5117
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 22152 5120 22385 5148
rect 22152 5108 22158 5120
rect 22373 5117 22385 5120
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 23109 5151 23167 5157
rect 23109 5117 23121 5151
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 19300 5052 19656 5080
rect 19300 5040 19306 5052
rect 17828 4984 19196 5012
rect 19628 5012 19656 5052
rect 20625 5083 20683 5089
rect 20625 5049 20637 5083
rect 20671 5049 20683 5083
rect 20625 5043 20683 5049
rect 20898 5040 20904 5092
rect 20956 5080 20962 5092
rect 21174 5080 21180 5092
rect 20956 5052 21180 5080
rect 20956 5040 20962 5052
rect 21174 5040 21180 5052
rect 21232 5040 21238 5092
rect 21450 5040 21456 5092
rect 21508 5080 21514 5092
rect 22830 5080 22836 5092
rect 21508 5052 22836 5080
rect 21508 5040 21514 5052
rect 22830 5040 22836 5052
rect 22888 5080 22894 5092
rect 23124 5080 23152 5111
rect 22888 5052 23152 5080
rect 22888 5040 22894 5052
rect 24210 5040 24216 5092
rect 24268 5080 24274 5092
rect 24578 5080 24584 5092
rect 24268 5052 24584 5080
rect 24268 5040 24274 5052
rect 24578 5040 24584 5052
rect 24636 5040 24642 5092
rect 20530 5012 20536 5024
rect 19628 4984 20536 5012
rect 17828 4972 17834 4984
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 20990 4972 20996 5024
rect 21048 5012 21054 5024
rect 25498 5012 25504 5024
rect 21048 4984 25504 5012
rect 21048 4972 21054 4984
rect 25498 4972 25504 4984
rect 25556 4972 25562 5024
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 1486 4768 1492 4820
rect 1544 4768 1550 4820
rect 2406 4768 2412 4820
rect 2464 4768 2470 4820
rect 3326 4808 3332 4820
rect 2516 4780 3332 4808
rect 2424 4740 2452 4768
rect 1964 4712 2452 4740
rect 1964 4681 1992 4712
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4641 2007 4675
rect 2314 4672 2320 4684
rect 1949 4635 2007 4641
rect 2148 4644 2320 4672
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 2148 4604 2176 4644
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 2406 4632 2412 4684
rect 2464 4632 2470 4684
rect 2516 4672 2544 4780
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3786 4768 3792 4820
rect 3844 4768 3850 4820
rect 5258 4808 5264 4820
rect 4356 4780 5264 4808
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 2516 4644 2697 4672
rect 2685 4641 2697 4644
rect 2731 4641 2743 4675
rect 2685 4635 2743 4641
rect 2823 4675 2881 4681
rect 2823 4641 2835 4675
rect 2869 4672 2881 4675
rect 3510 4672 3516 4684
rect 2869 4644 3516 4672
rect 2869 4641 2881 4644
rect 2823 4635 2881 4641
rect 3510 4632 3516 4644
rect 3568 4672 3574 4684
rect 4356 4672 4384 4780
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 12342 4808 12348 4820
rect 8904 4780 12348 4808
rect 8904 4768 8910 4780
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12636 4780 13308 4808
rect 5350 4700 5356 4752
rect 5408 4740 5414 4752
rect 10226 4740 10232 4752
rect 5408 4712 10232 4740
rect 5408 4700 5414 4712
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 11146 4700 11152 4752
rect 11204 4740 11210 4752
rect 12636 4740 12664 4780
rect 11204 4712 12664 4740
rect 13280 4740 13308 4780
rect 13354 4768 13360 4820
rect 13412 4808 13418 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13412 4780 13645 4808
rect 13412 4768 13418 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14458 4808 14464 4820
rect 14148 4780 14464 4808
rect 14148 4768 14154 4780
rect 14458 4768 14464 4780
rect 14516 4768 14522 4820
rect 16298 4808 16304 4820
rect 15396 4780 16304 4808
rect 13280 4712 14136 4740
rect 11204 4700 11210 4712
rect 3568 4644 4384 4672
rect 3568 4632 3574 4644
rect 7834 4632 7840 4684
rect 7892 4632 7898 4684
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 12158 4672 12164 4684
rect 9916 4644 12164 4672
rect 9916 4632 9922 4644
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 12636 4681 12664 4712
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 1811 4576 2176 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 1688 4468 1716 4567
rect 2958 4564 2964 4616
rect 3016 4564 3022 4616
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4604 4583 4607
rect 4706 4604 4712 4616
rect 4571 4576 4712 4604
rect 4571 4573 4583 4576
rect 4525 4567 4583 4573
rect 4262 4566 4292 4567
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 1688 4440 3617 4468
rect 3605 4437 3617 4440
rect 3651 4437 3663 4471
rect 3605 4431 3663 4437
rect 4062 4428 4068 4480
rect 4120 4428 4126 4480
rect 4262 4468 4290 4566
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 7852 4604 7880 4632
rect 14108 4616 14136 4712
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 15102 4672 15108 4684
rect 14424 4644 15108 4672
rect 14424 4632 14430 4644
rect 15102 4632 15108 4644
rect 15160 4672 15166 4684
rect 15396 4681 15424 4780
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 19242 4808 19248 4820
rect 17420 4780 19248 4808
rect 17420 4681 17448 4780
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 19613 4811 19671 4817
rect 19613 4808 19625 4811
rect 19576 4780 19625 4808
rect 19576 4768 19582 4780
rect 19613 4777 19625 4780
rect 19659 4777 19671 4811
rect 19613 4771 19671 4777
rect 21082 4768 21088 4820
rect 21140 4768 21146 4820
rect 21174 4768 21180 4820
rect 21232 4768 21238 4820
rect 21269 4811 21327 4817
rect 21269 4777 21281 4811
rect 21315 4808 21327 4811
rect 21542 4808 21548 4820
rect 21315 4780 21548 4808
rect 21315 4777 21327 4780
rect 21269 4771 21327 4777
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 23290 4808 23296 4820
rect 22112 4780 23296 4808
rect 18782 4700 18788 4752
rect 18840 4700 18846 4752
rect 18877 4743 18935 4749
rect 18877 4709 18889 4743
rect 18923 4709 18935 4743
rect 18877 4703 18935 4709
rect 15381 4675 15439 4681
rect 15381 4672 15393 4675
rect 15160 4644 15393 4672
rect 15160 4632 15166 4644
rect 15381 4641 15393 4644
rect 15427 4641 15439 4675
rect 15381 4635 15439 4641
rect 17405 4675 17463 4681
rect 17405 4641 17417 4675
rect 17451 4641 17463 4675
rect 18892 4672 18920 4703
rect 18966 4700 18972 4752
rect 19024 4740 19030 4752
rect 19337 4743 19395 4749
rect 19337 4740 19349 4743
rect 19024 4712 19349 4740
rect 19024 4700 19030 4712
rect 19337 4709 19349 4712
rect 19383 4709 19395 4743
rect 19337 4703 19395 4709
rect 19797 4743 19855 4749
rect 19797 4709 19809 4743
rect 19843 4740 19855 4743
rect 20898 4740 20904 4752
rect 19843 4712 20904 4740
rect 19843 4709 19855 4712
rect 19797 4703 19855 4709
rect 20898 4700 20904 4712
rect 20956 4700 20962 4752
rect 20993 4743 21051 4749
rect 20993 4709 21005 4743
rect 21039 4740 21051 4743
rect 21100 4740 21128 4768
rect 21039 4712 21128 4740
rect 21192 4740 21220 4768
rect 22005 4743 22063 4749
rect 22005 4740 22017 4743
rect 21192 4712 22017 4740
rect 21039 4709 21051 4712
rect 20993 4703 21051 4709
rect 22005 4709 22017 4712
rect 22051 4709 22063 4743
rect 22005 4703 22063 4709
rect 20714 4672 20720 4684
rect 18892 4644 20720 4672
rect 17405 4635 17463 4641
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 21082 4632 21088 4684
rect 21140 4672 21146 4684
rect 21140 4644 21312 4672
rect 21140 4632 21146 4644
rect 4948 4576 7880 4604
rect 4948 4564 4954 4576
rect 10318 4564 10324 4616
rect 10376 4604 10382 4616
rect 10870 4604 10876 4616
rect 10376 4576 10876 4604
rect 10376 4564 10382 4576
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 12895 4607 12953 4613
rect 12895 4604 12907 4607
rect 12860 4576 12907 4604
rect 12860 4564 12866 4576
rect 12895 4573 12907 4576
rect 12941 4573 12953 4607
rect 12895 4567 12953 4573
rect 14090 4564 14096 4616
rect 14148 4564 14154 4616
rect 14918 4564 14924 4616
rect 14976 4604 14982 4616
rect 16114 4604 16120 4616
rect 14976 4577 16120 4604
rect 14976 4576 15651 4577
rect 14976 4564 14982 4576
rect 8018 4496 8024 4548
rect 8076 4536 8082 4548
rect 14550 4536 14556 4548
rect 8076 4508 14556 4536
rect 8076 4496 8082 4508
rect 14550 4496 14556 4508
rect 14608 4496 14614 4548
rect 15639 4543 15651 4576
rect 15685 4576 16120 4577
rect 15685 4546 15698 4576
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 18598 4564 18604 4616
rect 18656 4604 18662 4616
rect 19061 4607 19119 4613
rect 19061 4604 19073 4607
rect 18656 4576 19073 4604
rect 18656 4564 18662 4576
rect 19061 4573 19073 4576
rect 19107 4573 19119 4607
rect 19061 4567 19119 4573
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19484 4576 19533 4604
rect 19484 4564 19490 4576
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 15685 4543 15697 4546
rect 15639 4537 15697 4543
rect 17672 4539 17730 4545
rect 17672 4505 17684 4539
rect 17718 4536 17730 4539
rect 17862 4536 17868 4548
rect 17718 4508 17868 4536
rect 17718 4505 17730 4508
rect 17672 4499 17730 4505
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 19720 4536 19748 4567
rect 19978 4564 19984 4616
rect 20036 4564 20042 4616
rect 20070 4564 20076 4616
rect 20128 4564 20134 4616
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4604 20315 4607
rect 20346 4604 20352 4616
rect 20303 4576 20352 4604
rect 20303 4573 20315 4576
rect 20257 4567 20315 4573
rect 20346 4564 20352 4576
rect 20404 4564 20410 4616
rect 20530 4564 20536 4616
rect 20588 4564 20594 4616
rect 20806 4564 20812 4616
rect 20864 4564 20870 4616
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21177 4607 21235 4613
rect 20947 4576 21036 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21008 4574 21036 4576
rect 21008 4546 21131 4574
rect 21177 4573 21189 4607
rect 21223 4604 21235 4607
rect 21284 4604 21312 4644
rect 21450 4632 21456 4684
rect 21508 4672 21514 4684
rect 22112 4672 22140 4780
rect 23290 4768 23296 4780
rect 23348 4768 23354 4820
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 25774 4808 25780 4820
rect 24075 4780 25780 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 21508 4644 22140 4672
rect 21508 4632 21514 4644
rect 22186 4632 22192 4684
rect 22244 4672 22250 4684
rect 22244 4644 22508 4672
rect 22244 4632 22250 4644
rect 22480 4616 22508 4644
rect 21223 4576 21312 4604
rect 21361 4607 21419 4613
rect 21223 4573 21235 4576
rect 21177 4567 21235 4573
rect 21361 4573 21373 4607
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21103 4536 21131 4546
rect 19720 4508 20668 4536
rect 21103 4508 21220 4536
rect 7742 4468 7748 4480
rect 4262 4440 7748 4468
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 20162 4468 20168 4480
rect 7892 4440 20168 4468
rect 7892 4428 7898 4440
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 20254 4428 20260 4480
rect 20312 4428 20318 4480
rect 20346 4428 20352 4480
rect 20404 4428 20410 4480
rect 20640 4477 20668 4508
rect 21192 4480 21220 4508
rect 20625 4471 20683 4477
rect 20625 4437 20637 4471
rect 20671 4437 20683 4471
rect 20625 4431 20683 4437
rect 21174 4428 21180 4480
rect 21232 4428 21238 4480
rect 21376 4468 21404 4567
rect 21634 4564 21640 4616
rect 21692 4564 21698 4616
rect 21818 4564 21824 4616
rect 21876 4564 21882 4616
rect 22281 4607 22339 4613
rect 22281 4573 22293 4607
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 22296 4536 22324 4567
rect 22462 4564 22468 4616
rect 22520 4564 22526 4616
rect 22739 4607 22797 4613
rect 22739 4573 22751 4607
rect 22785 4604 22797 4607
rect 23106 4604 23112 4616
rect 22785 4576 23112 4604
rect 22785 4573 22797 4576
rect 22739 4567 22797 4573
rect 23106 4564 23112 4576
rect 23164 4564 23170 4616
rect 23198 4536 23204 4548
rect 22296 4508 23204 4536
rect 23198 4496 23204 4508
rect 23256 4496 23262 4548
rect 23842 4496 23848 4548
rect 23900 4536 23906 4548
rect 23937 4539 23995 4545
rect 23937 4536 23949 4539
rect 23900 4508 23949 4536
rect 23900 4496 23906 4508
rect 23937 4505 23949 4508
rect 23983 4505 23995 4539
rect 23937 4499 23995 4505
rect 21453 4471 21511 4477
rect 21453 4468 21465 4471
rect 21376 4440 21465 4468
rect 21453 4437 21465 4440
rect 21499 4437 21511 4471
rect 21453 4431 21511 4437
rect 22094 4428 22100 4480
rect 22152 4428 22158 4480
rect 23477 4471 23535 4477
rect 23477 4437 23489 4471
rect 23523 4468 23535 4471
rect 23566 4468 23572 4480
rect 23523 4440 23572 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 4062 4264 4068 4276
rect 1688 4236 4068 4264
rect 1688 4205 1716 4236
rect 4062 4224 4068 4236
rect 4120 4224 4126 4276
rect 9122 4264 9128 4276
rect 8128 4236 9128 4264
rect 1673 4199 1731 4205
rect 1673 4165 1685 4199
rect 1719 4165 1731 4199
rect 5074 4196 5080 4208
rect 1673 4159 1731 4165
rect 4172 4168 5080 4196
rect 658 4088 664 4140
rect 716 4128 722 4140
rect 1854 4128 1860 4140
rect 716 4100 1860 4128
rect 716 4088 722 4100
rect 1854 4088 1860 4100
rect 1912 4088 1918 4140
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 1946 4020 1952 4072
rect 2004 4020 2010 4072
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 2096 3896 2145 3924
rect 2096 3884 2102 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2332 3924 2360 4091
rect 2590 4088 2596 4140
rect 2648 4088 2654 4140
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 3510 4137 3516 4140
rect 3467 4131 3516 4137
rect 3467 4097 3479 4131
rect 3513 4097 3516 4131
rect 3467 4091 3516 4097
rect 3510 4088 3516 4091
rect 3568 4088 3574 4140
rect 3602 4088 3608 4140
rect 3660 4088 3666 4140
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 3142 4060 3148 4072
rect 2455 4032 3148 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3344 4060 3372 4088
rect 4172 4060 4200 4168
rect 5074 4156 5080 4168
rect 5132 4156 5138 4208
rect 7374 4196 7380 4208
rect 6748 4168 7380 4196
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4295 4100 4537 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 6748 4137 6776 4168
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6144 4100 6745 4128
rect 6144 4088 6150 4100
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7007 4131 7065 4137
rect 7007 4097 7019 4131
rect 7053 4128 7065 4131
rect 7558 4128 7564 4140
rect 7053 4100 7564 4128
rect 7053 4097 7065 4100
rect 7007 4091 7065 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 3344 4032 4200 4060
rect 4338 4020 4344 4072
rect 4396 4020 4402 4072
rect 8128 4069 8156 4236
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10100 4236 11560 4264
rect 10100 4224 10106 4236
rect 10226 4196 10232 4208
rect 10152 4168 10232 4196
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 10152 4128 10180 4168
rect 10226 4156 10232 4168
rect 10284 4196 10290 4208
rect 10284 4168 10456 4196
rect 10284 4156 10290 4168
rect 10428 4140 10456 4168
rect 10318 4128 10324 4140
rect 9876 4100 10180 4128
rect 10279 4100 10324 4128
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8662 4060 8668 4072
rect 8343 4032 8668 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9033 4063 9091 4069
rect 9033 4060 9045 4063
rect 8864 4032 9045 4060
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 3053 3995 3111 4001
rect 3053 3992 3065 3995
rect 2556 3964 3065 3992
rect 2556 3952 2562 3964
rect 3053 3961 3065 3964
rect 3099 3961 3111 3995
rect 3053 3955 3111 3961
rect 4154 3924 4160 3936
rect 2332 3896 4160 3924
rect 2133 3887 2191 3893
rect 4154 3884 4160 3896
rect 4212 3884 4218 3936
rect 4356 3933 4384 4020
rect 8757 3995 8815 4001
rect 8757 3961 8769 3995
rect 8803 3961 8815 3995
rect 8757 3955 8815 3961
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3924 7803 3927
rect 8772 3924 8800 3955
rect 7791 3896 8800 3924
rect 8864 3924 8892 4032
rect 9033 4029 9045 4032
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9171 4063 9229 4069
rect 9171 4029 9183 4063
rect 9217 4060 9229 4063
rect 9876 4060 9904 4100
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10410 4088 10416 4140
rect 10468 4088 10474 4140
rect 11532 4137 11560 4236
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 13170 4264 13176 4276
rect 12400 4236 13176 4264
rect 12400 4224 12406 4236
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 14734 4224 14740 4276
rect 14792 4224 14798 4276
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 15344 4236 15577 4264
rect 15344 4224 15350 4236
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 16298 4224 16304 4276
rect 16356 4264 16362 4276
rect 19886 4264 19892 4276
rect 16356 4236 19892 4264
rect 16356 4224 16362 4236
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 20070 4224 20076 4276
rect 20128 4224 20134 4276
rect 20622 4224 20628 4276
rect 20680 4264 20686 4276
rect 20990 4264 20996 4276
rect 20680 4236 20996 4264
rect 20680 4224 20686 4236
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 21453 4267 21511 4273
rect 21453 4233 21465 4267
rect 21499 4264 21511 4267
rect 21634 4264 21640 4276
rect 21499 4236 21640 4264
rect 21499 4233 21511 4236
rect 21453 4227 21511 4233
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 12710 4196 12716 4208
rect 11900 4168 12716 4196
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4128 11575 4131
rect 11698 4128 11704 4140
rect 11563 4100 11704 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11791 4131 11849 4137
rect 11791 4097 11803 4131
rect 11837 4128 11849 4131
rect 11900 4128 11928 4168
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 11837 4100 11928 4128
rect 11837 4097 11849 4100
rect 11791 4091 11849 4097
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14424 4100 14565 4128
rect 14424 4088 14430 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14752 4128 14780 4224
rect 16758 4156 16764 4208
rect 16816 4196 16822 4208
rect 19245 4199 19303 4205
rect 19245 4196 19257 4199
rect 16816 4168 19257 4196
rect 16816 4156 16822 4168
rect 19245 4165 19257 4168
rect 19291 4165 19303 4199
rect 20088 4196 20116 4224
rect 23750 4196 23756 4208
rect 20088 4168 23756 4196
rect 19245 4159 19303 4165
rect 23750 4156 23756 4168
rect 23808 4156 23814 4208
rect 24305 4199 24363 4205
rect 24305 4165 24317 4199
rect 24351 4196 24363 4199
rect 24578 4196 24584 4208
rect 24351 4168 24584 4196
rect 24351 4165 24363 4168
rect 24305 4159 24363 4165
rect 24578 4156 24584 4168
rect 24636 4156 24642 4208
rect 14827 4131 14885 4137
rect 14827 4128 14839 4131
rect 14752 4100 14839 4128
rect 14553 4091 14611 4097
rect 14827 4097 14839 4100
rect 14873 4097 14885 4131
rect 14827 4091 14885 4097
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 17920 4100 18184 4128
rect 17920 4088 17926 4100
rect 9217 4032 9904 4060
rect 9217 4029 9229 4032
rect 9171 4023 9229 4029
rect 10042 4020 10048 4072
rect 10100 4020 10106 4072
rect 15562 4020 15568 4072
rect 15620 4060 15626 4072
rect 16206 4060 16212 4072
rect 15620 4032 16212 4060
rect 15620 4020 15626 4032
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 17954 4020 17960 4072
rect 18012 4020 18018 4072
rect 18156 4060 18184 4100
rect 18506 4088 18512 4140
rect 18564 4088 18570 4140
rect 18782 4088 18788 4140
rect 18840 4088 18846 4140
rect 19058 4088 19064 4140
rect 19116 4088 19122 4140
rect 19886 4088 19892 4140
rect 19944 4088 19950 4140
rect 20346 4137 20352 4140
rect 20340 4091 20352 4137
rect 20404 4128 20410 4140
rect 20622 4128 20628 4140
rect 20404 4100 20628 4128
rect 20346 4088 20352 4091
rect 20404 4088 20410 4100
rect 20622 4088 20628 4100
rect 20680 4088 20686 4140
rect 22370 4088 22376 4140
rect 22428 4088 22434 4140
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4097 22707 4131
rect 22649 4091 22707 4097
rect 18156 4032 18644 4060
rect 17681 3995 17739 4001
rect 17681 3961 17693 3995
rect 17727 3992 17739 3995
rect 17972 3992 18000 4020
rect 18616 4001 18644 4032
rect 19426 4020 19432 4072
rect 19484 4060 19490 4072
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 19484 4032 20085 4060
rect 19484 4020 19490 4032
rect 20073 4029 20085 4032
rect 20119 4029 20131 4063
rect 20073 4023 20131 4029
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22462 4060 22468 4072
rect 22051 4032 22468 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 22664 4060 22692 4091
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 22796 4100 23029 4128
rect 22796 4088 22802 4100
rect 23017 4097 23029 4100
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 24486 4088 24492 4140
rect 24544 4088 24550 4140
rect 23845 4063 23903 4069
rect 22664 4032 23796 4060
rect 17727 3964 18000 3992
rect 18601 3995 18659 4001
rect 17727 3961 17739 3964
rect 17681 3955 17739 3961
rect 18601 3961 18613 3995
rect 18647 3961 18659 3995
rect 18601 3955 18659 3961
rect 19242 3952 19248 4004
rect 19300 3992 19306 4004
rect 19705 3995 19763 4001
rect 19705 3992 19717 3995
rect 19300 3964 19717 3992
rect 19300 3952 19306 3964
rect 19705 3961 19717 3964
rect 19751 3961 19763 3995
rect 19705 3955 19763 3961
rect 21082 3952 21088 4004
rect 21140 3992 21146 4004
rect 22649 3995 22707 4001
rect 22649 3992 22661 3995
rect 21140 3964 22661 3992
rect 21140 3952 21146 3964
rect 22649 3961 22661 3964
rect 22695 3961 22707 3995
rect 23768 3992 23796 4032
rect 23845 4029 23857 4063
rect 23891 4060 23903 4063
rect 24210 4060 24216 4072
rect 23891 4032 24216 4060
rect 23891 4029 23903 4032
rect 23845 4023 23903 4029
rect 24210 4020 24216 4032
rect 24268 4020 24274 4072
rect 24118 3992 24124 4004
rect 23768 3964 24124 3992
rect 22649 3955 22707 3961
rect 24118 3952 24124 3964
rect 24176 3952 24182 4004
rect 9398 3924 9404 3936
rect 8864 3896 9404 3924
rect 7791 3893 7803 3896
rect 7745 3887 7803 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 9953 3927 10011 3933
rect 9953 3924 9965 3927
rect 9732 3896 9965 3924
rect 9732 3884 9738 3896
rect 9953 3893 9965 3896
rect 9999 3893 10011 3927
rect 9953 3887 10011 3893
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10376 3896 11069 3924
rect 10376 3884 10382 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 18322 3884 18328 3936
rect 18380 3884 18386 3936
rect 18690 3884 18696 3936
rect 18748 3924 18754 3936
rect 18877 3927 18935 3933
rect 18877 3924 18889 3927
rect 18748 3896 18889 3924
rect 18748 3884 18754 3896
rect 18877 3893 18889 3896
rect 18923 3893 18935 3927
rect 18877 3887 18935 3893
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19337 3927 19395 3933
rect 19337 3924 19349 3927
rect 19208 3896 19349 3924
rect 19208 3884 19214 3896
rect 19337 3893 19349 3896
rect 19383 3893 19395 3927
rect 19337 3887 19395 3893
rect 19610 3884 19616 3936
rect 19668 3924 19674 3936
rect 25130 3924 25136 3936
rect 19668 3896 25136 3924
rect 19668 3884 19674 3896
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 1578 3680 1584 3732
rect 1636 3680 1642 3732
rect 2130 3680 2136 3732
rect 2188 3680 2194 3732
rect 2682 3680 2688 3732
rect 2740 3680 2746 3732
rect 4890 3680 4896 3732
rect 4948 3680 4954 3732
rect 6362 3720 6368 3732
rect 5000 3692 6368 3720
rect 3694 3584 3700 3596
rect 1504 3556 3700 3584
rect 1504 3525 1532 3556
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 2501 3519 2559 3525
rect 2501 3485 2513 3519
rect 2547 3516 2559 3519
rect 5000 3516 5028 3692
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 9122 3720 9128 3732
rect 7208 3692 9128 3720
rect 7208 3661 7236 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9398 3680 9404 3732
rect 9456 3720 9462 3732
rect 11054 3720 11060 3732
rect 9456 3692 11060 3720
rect 9456 3680 9462 3692
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3621 7251 3655
rect 7193 3615 7251 3621
rect 7282 3612 7288 3664
rect 7340 3612 7346 3664
rect 7374 3612 7380 3664
rect 7432 3652 7438 3664
rect 8481 3655 8539 3661
rect 7432 3624 7512 3652
rect 7432 3612 7438 3624
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7300 3584 7328 3612
rect 7484 3593 7512 3624
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 9585 3655 9643 3661
rect 9585 3652 9597 3655
rect 8527 3624 9597 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 9585 3621 9597 3624
rect 9631 3621 9643 3655
rect 9585 3615 9643 3621
rect 7469 3587 7527 3593
rect 6963 3556 7420 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 2547 3488 5028 3516
rect 2547 3485 2559 3488
rect 2501 3479 2559 3485
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5351 3519 5409 3525
rect 5351 3485 5363 3519
rect 5397 3516 5409 3519
rect 5442 3516 5448 3528
rect 5397 3488 5448 3516
rect 5397 3485 5409 3488
rect 5351 3479 5409 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 7392 3525 7420 3556
rect 7469 3553 7481 3587
rect 7515 3553 7527 3587
rect 7469 3547 7527 3553
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9030 3584 9036 3596
rect 8987 3556 9036 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9490 3584 9496 3596
rect 9140 3556 9496 3584
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7743 3519 7801 3525
rect 7743 3485 7755 3519
rect 7789 3516 7801 3519
rect 8846 3516 8852 3528
rect 7789 3488 8852 3516
rect 7789 3485 7801 3488
rect 7743 3479 7801 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9140 3525 9168 3556
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9692 3584 9720 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11146 3680 11152 3732
rect 11204 3720 11210 3732
rect 12066 3720 12072 3732
rect 11204 3692 12072 3720
rect 11204 3680 11210 3692
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 13964 3692 15117 3720
rect 13964 3680 13970 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 15105 3683 15163 3689
rect 18233 3723 18291 3729
rect 18233 3689 18245 3723
rect 18279 3720 18291 3723
rect 18414 3720 18420 3732
rect 18279 3692 18420 3720
rect 18279 3689 18291 3692
rect 18233 3683 18291 3689
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 20625 3723 20683 3729
rect 18524 3692 20576 3720
rect 18524 3661 18552 3692
rect 13541 3655 13599 3661
rect 13541 3621 13553 3655
rect 13587 3621 13599 3655
rect 13541 3615 13599 3621
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3621 18567 3655
rect 20548 3652 20576 3692
rect 20625 3689 20637 3723
rect 20671 3720 20683 3723
rect 20806 3720 20812 3732
rect 20671 3692 20812 3720
rect 20671 3689 20683 3692
rect 20625 3683 20683 3689
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21284 3692 22692 3720
rect 20548 3624 20944 3652
rect 18509 3615 18567 3621
rect 10042 3593 10048 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9692 3556 9873 3584
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 9999 3587 10048 3593
rect 9999 3553 10011 3587
rect 10045 3553 10048 3587
rect 9999 3547 10048 3553
rect 10042 3544 10048 3547
rect 10100 3544 10106 3596
rect 10502 3584 10508 3596
rect 10152 3556 10508 3584
rect 10152 3525 10180 3556
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 12526 3544 12532 3596
rect 12584 3544 12590 3596
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 13556 3584 13584 3615
rect 13228 3556 13584 3584
rect 18064 3556 19380 3584
rect 13228 3544 13234 3556
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 2038 3408 2044 3460
rect 2096 3408 2102 3460
rect 2332 3420 2774 3448
rect 2332 3392 2360 3420
rect 2314 3340 2320 3392
rect 2372 3340 2378 3392
rect 2746 3380 2774 3420
rect 3786 3408 3792 3460
rect 3844 3448 3850 3460
rect 4801 3451 4859 3457
rect 4801 3448 4813 3451
rect 3844 3420 4813 3448
rect 3844 3408 3850 3420
rect 4801 3417 4813 3420
rect 4847 3448 4859 3451
rect 8294 3448 8300 3460
rect 4847 3420 8300 3448
rect 4847 3417 4859 3420
rect 4801 3411 4859 3417
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 9140 3448 9168 3479
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 11790 3476 11796 3528
rect 11848 3476 11854 3528
rect 13630 3516 13636 3528
rect 12084 3488 13636 3516
rect 8720 3420 9168 3448
rect 8720 3408 8726 3420
rect 10686 3408 10692 3460
rect 10744 3448 10750 3460
rect 12084 3457 12112 3488
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13688 3488 13737 3516
rect 13688 3476 13694 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 14090 3476 14096 3528
rect 14148 3476 14154 3528
rect 14274 3476 14280 3528
rect 14332 3516 14338 3528
rect 14367 3519 14425 3525
rect 14367 3516 14379 3519
rect 14332 3488 14379 3516
rect 14332 3476 14338 3488
rect 14367 3485 14379 3488
rect 14413 3516 14425 3519
rect 14826 3516 14832 3528
rect 14413 3488 14832 3516
rect 14413 3485 14425 3488
rect 14367 3479 14425 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 16298 3476 16304 3528
rect 16356 3476 16362 3528
rect 17218 3476 17224 3528
rect 17276 3476 17282 3528
rect 17310 3476 17316 3528
rect 17368 3476 17374 3528
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 18064 3525 18092 3556
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18371 3488 18552 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 12069 3451 12127 3457
rect 10744 3420 11744 3448
rect 10744 3408 10750 3420
rect 5166 3380 5172 3392
rect 2746 3352 5172 3380
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 6086 3340 6092 3392
rect 6144 3340 6150 3392
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 10781 3383 10839 3389
rect 10781 3380 10793 3383
rect 6512 3352 10793 3380
rect 6512 3340 6518 3352
rect 10781 3349 10793 3352
rect 10827 3349 10839 3383
rect 10781 3343 10839 3349
rect 11330 3340 11336 3392
rect 11388 3340 11394 3392
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 11716 3380 11744 3420
rect 12069 3417 12081 3451
rect 12115 3417 12127 3451
rect 12069 3411 12127 3417
rect 12342 3408 12348 3460
rect 12400 3408 12406 3460
rect 12434 3408 12440 3460
rect 12492 3408 12498 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 12584 3420 12817 3448
rect 12584 3408 12590 3420
rect 12805 3417 12817 3420
rect 12851 3417 12863 3451
rect 12805 3411 12863 3417
rect 12894 3408 12900 3460
rect 12952 3448 12958 3460
rect 14108 3448 14136 3476
rect 16316 3448 16344 3476
rect 17328 3448 17356 3476
rect 18524 3460 18552 3488
rect 18708 3488 19196 3516
rect 12952 3420 13400 3448
rect 14108 3420 16344 3448
rect 16408 3420 17356 3448
rect 18156 3420 18368 3448
rect 12952 3408 12958 3420
rect 13372 3389 13400 3420
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 11716 3352 13185 3380
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3380 13415 3383
rect 16408 3380 16436 3420
rect 13403 3352 16436 3380
rect 17037 3383 17095 3389
rect 13403 3349 13415 3352
rect 13357 3343 13415 3349
rect 17037 3349 17049 3383
rect 17083 3380 17095 3383
rect 17402 3380 17408 3392
rect 17083 3352 17408 3380
rect 17083 3349 17095 3352
rect 17037 3343 17095 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17770 3340 17776 3392
rect 17828 3340 17834 3392
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 18156 3380 18184 3420
rect 18104 3352 18184 3380
rect 18340 3380 18368 3420
rect 18506 3408 18512 3460
rect 18564 3408 18570 3460
rect 18708 3457 18736 3488
rect 18693 3451 18751 3457
rect 18693 3417 18705 3451
rect 18739 3417 18751 3451
rect 18693 3411 18751 3417
rect 19061 3451 19119 3457
rect 19061 3417 19073 3451
rect 19107 3417 19119 3451
rect 19168 3448 19196 3488
rect 19242 3476 19248 3528
rect 19300 3476 19306 3528
rect 19352 3516 19380 3556
rect 19512 3519 19570 3525
rect 19352 3488 19472 3516
rect 19444 3448 19472 3488
rect 19512 3485 19524 3519
rect 19558 3516 19570 3519
rect 19886 3516 19892 3528
rect 19558 3488 19892 3516
rect 19558 3485 19570 3488
rect 19512 3479 19570 3485
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20772 3488 20821 3516
rect 20772 3476 20778 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20916 3516 20944 3624
rect 20990 3544 20996 3596
rect 21048 3584 21054 3596
rect 21284 3593 21312 3692
rect 22664 3593 22692 3692
rect 23661 3655 23719 3661
rect 23661 3621 23673 3655
rect 23707 3652 23719 3655
rect 23750 3652 23756 3664
rect 23707 3624 23756 3652
rect 23707 3621 23719 3624
rect 23661 3615 23719 3621
rect 23750 3612 23756 3624
rect 23808 3652 23814 3664
rect 24210 3652 24216 3664
rect 23808 3624 24216 3652
rect 23808 3612 23814 3624
rect 24210 3612 24216 3624
rect 24268 3612 24274 3664
rect 21269 3587 21327 3593
rect 21269 3584 21281 3587
rect 21048 3556 21281 3584
rect 21048 3544 21054 3556
rect 21269 3553 21281 3556
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 22649 3587 22707 3593
rect 22649 3553 22661 3587
rect 22695 3553 22707 3587
rect 22649 3547 22707 3553
rect 21450 3516 21456 3528
rect 20916 3488 21456 3516
rect 20809 3479 20867 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 21543 3519 21601 3525
rect 21543 3485 21555 3519
rect 21589 3516 21601 3519
rect 21634 3516 21640 3528
rect 21589 3488 21640 3516
rect 21589 3485 21601 3488
rect 21543 3479 21601 3485
rect 21634 3476 21640 3488
rect 21692 3476 21698 3528
rect 22922 3476 22928 3528
rect 22980 3476 22986 3528
rect 24213 3519 24271 3525
rect 24213 3485 24225 3519
rect 24259 3485 24271 3519
rect 24213 3479 24271 3485
rect 19978 3448 19984 3460
rect 19168 3420 19380 3448
rect 19444 3420 19984 3448
rect 19061 3411 19119 3417
rect 18782 3380 18788 3392
rect 18340 3352 18788 3380
rect 18104 3340 18110 3352
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 19076 3380 19104 3411
rect 19352 3392 19380 3420
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 24228 3448 24256 3479
rect 20680 3420 24256 3448
rect 20680 3408 20686 3420
rect 19242 3380 19248 3392
rect 19076 3352 19248 3380
rect 19242 3340 19248 3352
rect 19300 3340 19306 3392
rect 19334 3340 19340 3392
rect 19392 3340 19398 3392
rect 19702 3340 19708 3392
rect 19760 3380 19766 3392
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 19760 3352 20913 3380
rect 19760 3340 19766 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 22281 3383 22339 3389
rect 22281 3349 22293 3383
rect 22327 3380 22339 3383
rect 22462 3380 22468 3392
rect 22327 3352 22468 3380
rect 22327 3349 22339 3352
rect 22281 3343 22339 3349
rect 22462 3340 22468 3352
rect 22520 3380 22526 3392
rect 22922 3380 22928 3392
rect 22520 3352 22928 3380
rect 22520 3340 22526 3352
rect 22922 3340 22928 3352
rect 22980 3340 22986 3392
rect 23750 3340 23756 3392
rect 23808 3380 23814 3392
rect 24029 3383 24087 3389
rect 24029 3380 24041 3383
rect 23808 3352 24041 3380
rect 23808 3340 23814 3352
rect 24029 3349 24041 3352
rect 24075 3349 24087 3383
rect 24029 3343 24087 3349
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 2038 3176 2044 3188
rect 1811 3148 2044 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3326 3136 3332 3188
rect 3384 3136 3390 3188
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 4430 3176 4436 3188
rect 3743 3148 4436 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 4522 3136 4528 3188
rect 4580 3136 4586 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6328 3148 6561 3176
rect 6328 3136 6334 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 6696 3148 8033 3176
rect 6696 3136 6702 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 9674 3176 9680 3188
rect 8352 3148 9680 3176
rect 8352 3136 8358 3148
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9876 3148 10180 3176
rect 9876 3120 9904 3148
rect 2314 3108 2320 3120
rect 1964 3080 2320 3108
rect 1026 3000 1032 3052
rect 1084 3040 1090 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 1084 3012 1501 3040
rect 1084 3000 1090 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 1489 3003 1547 3009
rect 1762 3000 1768 3052
rect 1820 3000 1826 3052
rect 1964 3049 1992 3080
rect 2314 3068 2320 3080
rect 2372 3068 2378 3120
rect 6454 3108 6460 3120
rect 2746 3080 6460 3108
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2746 3040 2774 3080
rect 6454 3068 6460 3080
rect 6512 3068 6518 3120
rect 7653 3111 7711 3117
rect 7653 3108 7665 3111
rect 6656 3080 7665 3108
rect 2271 3012 2774 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 3200 3012 3249 3040
rect 3200 3000 3206 3012
rect 3237 3009 3249 3012
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 1780 2972 1808 3000
rect 1596 2944 1808 2972
rect 1596 2836 1624 2944
rect 2682 2932 2688 2984
rect 2740 2972 2746 2984
rect 3528 2972 3556 3003
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 6656 3040 6684 3080
rect 7653 3077 7665 3080
rect 7699 3077 7711 3111
rect 7653 3071 7711 3077
rect 9401 3111 9459 3117
rect 9401 3077 9413 3111
rect 9447 3108 9459 3111
rect 9858 3108 9864 3120
rect 9447 3080 9864 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 9858 3068 9864 3080
rect 9916 3068 9922 3120
rect 9953 3111 10011 3117
rect 9953 3077 9965 3111
rect 9999 3077 10011 3111
rect 10152 3108 10180 3148
rect 10410 3136 10416 3188
rect 10468 3176 10474 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 10468 3148 11253 3176
rect 10468 3136 10474 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 11241 3139 11299 3145
rect 11974 3136 11980 3188
rect 12032 3136 12038 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 12492 3148 13185 3176
rect 12492 3136 12498 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 14274 3136 14280 3188
rect 14332 3136 14338 3188
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 19153 3179 19211 3185
rect 18564 3148 19104 3176
rect 18564 3136 18570 3148
rect 10208 3111 10266 3117
rect 10208 3108 10220 3111
rect 10152 3080 10220 3108
rect 9953 3071 10011 3077
rect 10208 3077 10220 3080
rect 10254 3077 10266 3111
rect 10208 3071 10266 3077
rect 4488 3012 6684 3040
rect 4488 3000 4494 3012
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 7282 3000 7288 3052
rect 7340 3000 7346 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8205 3043 8263 3049
rect 8205 3040 8217 3043
rect 7800 3012 8217 3040
rect 7800 3000 7806 3012
rect 8205 3009 8217 3012
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 2740 2944 3556 2972
rect 2740 2932 2746 2944
rect 6086 2932 6092 2984
rect 6144 2972 6150 2984
rect 8496 2972 8524 3003
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 9968 3040 9996 3071
rect 10318 3068 10324 3120
rect 10376 3068 10382 3120
rect 10428 3080 11008 3108
rect 10428 3040 10456 3080
rect 9968 3012 10456 3040
rect 10686 3000 10692 3052
rect 10744 3000 10750 3052
rect 10980 3040 11008 3080
rect 11054 3068 11060 3120
rect 11112 3068 11118 3120
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 10980 3012 11713 3040
rect 11701 3009 11713 3012
rect 11747 3040 11759 3043
rect 11992 3040 12020 3136
rect 12618 3108 12624 3120
rect 12452 3080 12624 3108
rect 12452 3079 12480 3080
rect 12419 3073 12480 3079
rect 11747 3012 12020 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 12066 3000 12072 3052
rect 12124 3000 12130 3052
rect 12419 3039 12431 3073
rect 12465 3042 12480 3073
rect 12618 3068 12624 3080
rect 12676 3108 12682 3120
rect 14292 3108 14320 3136
rect 18230 3108 18236 3120
rect 12676 3080 14320 3108
rect 17972 3080 18236 3108
rect 12676 3068 12682 3080
rect 12465 3039 12477 3042
rect 12419 3033 12477 3039
rect 15654 3000 15660 3052
rect 15712 3000 15718 3052
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 16991 3012 17417 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17405 3009 17417 3012
rect 17451 3040 17463 3043
rect 17586 3040 17592 3052
rect 17451 3012 17592 3040
rect 17451 3009 17463 3012
rect 17405 3003 17463 3009
rect 17586 3000 17592 3012
rect 17644 3000 17650 3052
rect 17678 3000 17684 3052
rect 17736 3000 17742 3052
rect 17972 3049 18000 3080
rect 18230 3068 18236 3080
rect 18288 3068 18294 3120
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 18693 3111 18751 3117
rect 18693 3108 18705 3111
rect 18656 3080 18705 3108
rect 18656 3068 18662 3080
rect 18693 3077 18705 3080
rect 18739 3077 18751 3111
rect 19076 3108 19104 3148
rect 19153 3145 19165 3179
rect 19199 3176 19211 3179
rect 19886 3176 19892 3188
rect 19199 3148 19892 3176
rect 19199 3145 19211 3148
rect 19153 3139 19211 3145
rect 19886 3136 19892 3148
rect 19944 3136 19950 3188
rect 19996 3148 22876 3176
rect 19996 3108 20024 3148
rect 19076 3080 20024 3108
rect 18693 3071 18751 3077
rect 20898 3068 20904 3120
rect 20956 3108 20962 3120
rect 21913 3111 21971 3117
rect 21913 3108 21925 3111
rect 20956 3080 21925 3108
rect 20956 3068 20962 3080
rect 21913 3077 21925 3080
rect 21959 3077 21971 3111
rect 22848 3108 22876 3148
rect 24026 3136 24032 3188
rect 24084 3176 24090 3188
rect 24305 3179 24363 3185
rect 24305 3176 24317 3179
rect 24084 3148 24317 3176
rect 24084 3136 24090 3148
rect 24305 3145 24317 3148
rect 24351 3145 24363 3179
rect 24305 3139 24363 3145
rect 23078 3111 23136 3117
rect 23078 3108 23090 3111
rect 21913 3071 21971 3077
rect 22112 3080 22598 3108
rect 22848 3080 23090 3108
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3009 18015 3043
rect 17957 3003 18015 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3040 18383 3043
rect 19058 3040 19064 3052
rect 18371 3012 19064 3040
rect 18371 3009 18383 3012
rect 18325 3003 18383 3009
rect 9582 2972 9588 2984
rect 6144 2944 6394 2972
rect 8496 2944 9588 2972
rect 6144 2932 6150 2944
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 10778 2932 10784 2984
rect 10836 2932 10842 2984
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 11974 2972 11980 2984
rect 11848 2944 11980 2972
rect 11848 2932 11854 2944
rect 11974 2932 11980 2944
rect 12032 2972 12038 2984
rect 12161 2975 12219 2981
rect 12161 2972 12173 2975
rect 12032 2944 12173 2972
rect 12032 2932 12038 2944
rect 12161 2941 12173 2944
rect 12207 2941 12219 2975
rect 18064 2972 18092 3003
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3040 19395 3043
rect 20714 3040 20720 3052
rect 19383 3012 20720 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21266 3040 21272 3052
rect 20855 3012 21272 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 22112 2984 22140 3080
rect 22465 3043 22523 3049
rect 22465 3009 22477 3043
rect 22511 3009 22523 3043
rect 22570 3040 22598 3080
rect 23078 3077 23090 3080
rect 23124 3077 23136 3111
rect 23078 3071 23136 3077
rect 23382 3068 23388 3120
rect 23440 3068 23446 3120
rect 22833 3043 22891 3049
rect 22833 3040 22845 3043
rect 22570 3012 22845 3040
rect 22465 3003 22523 3009
rect 22833 3009 22845 3012
rect 22879 3009 22891 3043
rect 23400 3040 23428 3068
rect 23400 3012 23888 3040
rect 22833 3003 22891 3009
rect 19521 2975 19579 2981
rect 18064 2944 19472 2972
rect 12161 2935 12219 2941
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 5350 2904 5356 2916
rect 1719 2876 5356 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 6178 2864 6184 2916
rect 6236 2904 6242 2916
rect 6454 2904 6460 2916
rect 6236 2876 6460 2904
rect 6236 2864 6242 2876
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 7837 2907 7895 2913
rect 7837 2873 7849 2907
rect 7883 2904 7895 2907
rect 8110 2904 8116 2916
rect 7883 2876 8116 2904
rect 7883 2873 7895 2876
rect 7837 2867 7895 2873
rect 8110 2864 8116 2876
rect 8168 2864 8174 2916
rect 18966 2904 18972 2916
rect 11532 2876 12018 2904
rect 2041 2839 2099 2845
rect 2041 2836 2053 2839
rect 1596 2808 2053 2836
rect 2041 2805 2053 2808
rect 2087 2805 2099 2839
rect 2041 2799 2099 2805
rect 8294 2796 8300 2848
rect 8352 2796 8358 2848
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 11532 2845 11560 2876
rect 8941 2839 8999 2845
rect 8941 2836 8953 2839
rect 8628 2808 8953 2836
rect 8628 2796 8634 2808
rect 8941 2805 8953 2808
rect 8987 2805 8999 2839
rect 8941 2799 8999 2805
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2805 11575 2839
rect 11517 2799 11575 2805
rect 11882 2796 11888 2848
rect 11940 2796 11946 2848
rect 11990 2836 12018 2876
rect 18248 2876 18972 2904
rect 13446 2836 13452 2848
rect 11990 2808 13452 2836
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 15470 2796 15476 2848
rect 15528 2796 15534 2848
rect 17218 2796 17224 2848
rect 17276 2796 17282 2848
rect 17494 2796 17500 2848
rect 17552 2796 17558 2848
rect 17770 2796 17776 2848
rect 17828 2796 17834 2848
rect 18248 2845 18276 2876
rect 18966 2864 18972 2876
rect 19024 2864 19030 2916
rect 19444 2904 19472 2944
rect 19521 2941 19533 2975
rect 19567 2972 19579 2975
rect 19610 2972 19616 2984
rect 19567 2944 19616 2972
rect 19567 2941 19579 2944
rect 19521 2935 19579 2941
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 19794 2932 19800 2984
rect 19852 2932 19858 2984
rect 20438 2932 20444 2984
rect 20496 2972 20502 2984
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20496 2944 21005 2972
rect 20496 2932 20502 2944
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 22094 2932 22100 2984
rect 22152 2932 22158 2984
rect 20622 2904 20628 2916
rect 19444 2876 20628 2904
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 22480 2904 22508 3003
rect 22830 2904 22836 2916
rect 22480 2876 22836 2904
rect 22830 2864 22836 2876
rect 22888 2864 22894 2916
rect 23860 2904 23888 3012
rect 24302 3000 24308 3052
rect 24360 3040 24366 3052
rect 24489 3043 24547 3049
rect 24489 3040 24501 3043
rect 24360 3012 24501 3040
rect 24360 3000 24366 3012
rect 24489 3009 24501 3012
rect 24535 3009 24547 3043
rect 24489 3003 24547 3009
rect 25406 2932 25412 2984
rect 25464 2932 25470 2984
rect 24213 2907 24271 2913
rect 24213 2904 24225 2907
rect 23860 2876 24225 2904
rect 24213 2873 24225 2876
rect 24259 2873 24271 2907
rect 25424 2904 25452 2932
rect 24213 2867 24271 2873
rect 24320 2876 25452 2904
rect 18233 2839 18291 2845
rect 18233 2805 18245 2839
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 18782 2796 18788 2848
rect 18840 2796 18846 2848
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 20036 2808 22017 2836
rect 20036 2796 20042 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 24320 2836 24348 2876
rect 22603 2808 24348 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 382 2592 388 2644
rect 440 2632 446 2644
rect 1949 2635 2007 2641
rect 1949 2632 1961 2635
rect 440 2604 1961 2632
rect 440 2592 446 2604
rect 1949 2601 1961 2604
rect 1995 2601 2007 2635
rect 1949 2595 2007 2601
rect 2332 2604 2912 2632
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 2332 2564 2360 2604
rect 1719 2536 2360 2564
rect 2884 2564 2912 2604
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 3016 2604 3249 2632
rect 3016 2592 3022 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 3694 2592 3700 2644
rect 3752 2592 3758 2644
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 3973 2635 4031 2641
rect 3973 2632 3985 2635
rect 3844 2604 3985 2632
rect 3844 2592 3850 2604
rect 3973 2601 3985 2604
rect 4019 2601 4031 2635
rect 3973 2595 4031 2601
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 5626 2632 5632 2644
rect 4755 2604 5632 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6825 2635 6883 2641
rect 5920 2604 6776 2632
rect 3712 2564 3740 2592
rect 2884 2536 3740 2564
rect 5537 2567 5595 2573
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 5537 2533 5549 2567
rect 5583 2564 5595 2567
rect 5920 2564 5948 2604
rect 5583 2536 5948 2564
rect 6748 2564 6776 2604
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 6914 2632 6920 2644
rect 6871 2604 6920 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 8294 2632 8300 2644
rect 7432 2604 8300 2632
rect 7432 2592 7438 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8444 2604 9628 2632
rect 8444 2592 8450 2604
rect 9600 2564 9628 2604
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 9732 2604 10548 2632
rect 9732 2592 9738 2604
rect 9766 2564 9772 2576
rect 6748 2536 9536 2564
rect 9600 2536 9772 2564
rect 5583 2533 5595 2536
rect 5537 2527 5595 2533
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 5316 2468 5825 2496
rect 5316 2456 5322 2468
rect 5813 2465 5825 2468
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 474 2388 480 2440
rect 532 2428 538 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 532 2400 1777 2428
rect 532 2388 538 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2499 2431 2557 2437
rect 2499 2397 2511 2431
rect 2545 2428 2557 2431
rect 3050 2428 3056 2440
rect 2545 2400 3056 2428
rect 2545 2397 2557 2400
rect 2499 2391 2557 2397
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 256 2332 1501 2360
rect 256 2320 262 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 1670 2320 1676 2372
rect 1728 2360 1734 2372
rect 2240 2360 2268 2391
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3292 2400 3801 2428
rect 3292 2388 3298 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 4982 2388 4988 2440
rect 5040 2388 5046 2440
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 5736 2360 5764 2391
rect 1728 2332 2268 2360
rect 2332 2332 5396 2360
rect 1728 2320 1734 2332
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 2332 2292 2360 2332
rect 5368 2304 5396 2332
rect 5460 2332 5764 2360
rect 5828 2360 5856 2459
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7742 2496 7748 2508
rect 7524 2468 7748 2496
rect 7524 2456 7530 2468
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8386 2496 8392 2508
rect 8036 2468 8392 2496
rect 6087 2431 6145 2437
rect 6087 2397 6099 2431
rect 6133 2428 6145 2431
rect 6454 2428 6460 2440
rect 6133 2400 6460 2428
rect 6133 2397 6145 2400
rect 6087 2391 6145 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 7561 2431 7619 2437
rect 7561 2397 7573 2431
rect 7607 2428 7619 2431
rect 7650 2428 7656 2440
rect 7607 2400 7656 2428
rect 7607 2397 7619 2400
rect 7561 2391 7619 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8036 2360 8064 2468
rect 8386 2456 8392 2468
rect 8444 2456 8450 2508
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 9508 2496 9536 2536
rect 9766 2524 9772 2536
rect 9824 2564 9830 2576
rect 10520 2564 10548 2604
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10836 2604 10885 2632
rect 10836 2592 10842 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 13262 2592 13268 2644
rect 13320 2632 13326 2644
rect 13538 2632 13544 2644
rect 13320 2604 13544 2632
rect 13320 2592 13326 2604
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 14921 2635 14979 2641
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15378 2632 15384 2644
rect 14967 2604 15384 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 15378 2592 15384 2604
rect 15436 2632 15442 2644
rect 16114 2632 16120 2644
rect 15436 2604 16120 2632
rect 15436 2592 15442 2604
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 16666 2592 16672 2644
rect 16724 2592 16730 2644
rect 16758 2592 16764 2644
rect 16816 2592 16822 2644
rect 19426 2632 19432 2644
rect 16868 2604 19432 2632
rect 11256 2564 11284 2592
rect 9824 2536 9904 2564
rect 10520 2536 11284 2564
rect 11609 2567 11667 2573
rect 9824 2524 9830 2536
rect 9876 2505 9904 2536
rect 11609 2533 11621 2567
rect 11655 2564 11667 2567
rect 12158 2564 12164 2576
rect 11655 2536 12164 2564
rect 11655 2533 11667 2536
rect 11609 2527 11667 2533
rect 12158 2524 12164 2536
rect 12216 2524 12222 2576
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 13906 2564 13912 2576
rect 13403 2536 13912 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 16868 2564 16896 2604
rect 19426 2592 19432 2604
rect 19484 2592 19490 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 20070 2632 20076 2644
rect 19576 2604 20076 2632
rect 19576 2592 19582 2604
rect 20070 2592 20076 2604
rect 20128 2632 20134 2644
rect 22094 2632 22100 2644
rect 20128 2604 22100 2632
rect 20128 2592 20134 2604
rect 14016 2536 16896 2564
rect 9861 2499 9919 2505
rect 8536 2468 9352 2496
rect 9508 2468 9812 2496
rect 8536 2456 8542 2468
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2428 8355 2431
rect 8570 2428 8576 2440
rect 8343 2400 8576 2428
rect 8343 2397 8355 2400
rect 8297 2391 8355 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 5828 2332 8064 2360
rect 5460 2304 5488 2332
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 8260 2332 8432 2360
rect 8260 2320 8266 2332
rect 992 2264 2360 2292
rect 4801 2295 4859 2301
rect 992 2252 998 2264
rect 4801 2261 4813 2295
rect 4847 2292 4859 2295
rect 5074 2292 5080 2304
rect 4847 2264 5080 2292
rect 4847 2261 4859 2264
rect 4801 2255 4859 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5258 2252 5264 2304
rect 5316 2252 5322 2304
rect 5350 2252 5356 2304
rect 5408 2252 5414 2304
rect 5442 2252 5448 2304
rect 5500 2252 5506 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 6512 2264 7389 2292
rect 6512 2252 6518 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7377 2255 7435 2261
rect 7466 2252 7472 2304
rect 7524 2292 7530 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7524 2264 7665 2292
rect 7524 2252 7530 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8404 2301 8432 2332
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 8772 2360 8800 2391
rect 8938 2388 8944 2440
rect 8996 2428 9002 2440
rect 9324 2437 9352 2468
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8996 2400 9137 2428
rect 8996 2388 9002 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9674 2428 9680 2440
rect 9309 2391 9367 2397
rect 9646 2388 9680 2428
rect 9732 2388 9738 2440
rect 9646 2360 9674 2388
rect 8536 2332 8800 2360
rect 9600 2332 9674 2360
rect 9784 2360 9812 2468
rect 9861 2465 9873 2499
rect 9907 2465 9919 2499
rect 9861 2459 9919 2465
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 14016 2496 14044 2536
rect 19058 2524 19064 2576
rect 19116 2564 19122 2576
rect 19610 2564 19616 2576
rect 19116 2536 19616 2564
rect 19116 2524 19122 2536
rect 19610 2524 19616 2536
rect 19668 2524 19674 2576
rect 21008 2536 21496 2564
rect 12032 2468 14044 2496
rect 12032 2456 12038 2468
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 16393 2499 16451 2505
rect 14516 2468 15700 2496
rect 14516 2456 14522 2468
rect 10135 2431 10193 2437
rect 10135 2397 10147 2431
rect 10181 2428 10193 2431
rect 10594 2428 10600 2440
rect 10181 2400 10600 2428
rect 10181 2397 10193 2400
rect 10135 2391 10193 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 11514 2388 11520 2440
rect 11572 2388 11578 2440
rect 11790 2388 11796 2440
rect 11848 2388 11854 2440
rect 12066 2388 12072 2440
rect 12124 2388 12130 2440
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12483 2400 12909 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12897 2397 12909 2400
rect 12943 2428 12955 2431
rect 13262 2428 13268 2440
rect 12943 2400 13268 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13538 2388 13544 2440
rect 13596 2388 13602 2440
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14366 2428 14372 2440
rect 14056 2400 14372 2428
rect 14056 2388 14062 2400
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 15378 2388 15384 2440
rect 15436 2388 15442 2440
rect 15672 2437 15700 2468
rect 16393 2465 16405 2499
rect 16439 2496 16451 2499
rect 17034 2496 17040 2508
rect 16439 2468 17040 2496
rect 16439 2465 16451 2468
rect 16393 2459 16451 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 18966 2496 18972 2508
rect 17144 2468 18972 2496
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2428 15991 2431
rect 16206 2428 16212 2440
rect 15979 2400 16212 2428
rect 15979 2397 15991 2400
rect 15933 2391 15991 2397
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 17052 2428 17080 2456
rect 16991 2400 17080 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 12526 2360 12532 2372
rect 9784 2332 12532 2360
rect 8536 2320 8542 2332
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2261 8447 2295
rect 8389 2255 8447 2261
rect 8570 2252 8576 2304
rect 8628 2252 8634 2304
rect 8938 2252 8944 2304
rect 8996 2252 9002 2304
rect 9493 2295 9551 2301
rect 9493 2261 9505 2295
rect 9539 2292 9551 2295
rect 9600 2292 9628 2332
rect 12526 2320 12532 2332
rect 12584 2320 12590 2372
rect 15102 2320 15108 2372
rect 15160 2360 15166 2372
rect 16500 2360 16528 2391
rect 17144 2360 17172 2468
rect 18966 2456 18972 2468
rect 19024 2496 19030 2508
rect 21008 2496 21036 2536
rect 19024 2468 21036 2496
rect 19024 2456 19030 2468
rect 21082 2456 21088 2508
rect 21140 2456 21146 2508
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 17678 2428 17684 2440
rect 17267 2400 17684 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 17920 2400 18705 2428
rect 17920 2388 17926 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 19334 2388 19340 2440
rect 19392 2388 19398 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 20625 2431 20683 2437
rect 19475 2400 19564 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 15160 2332 15792 2360
rect 16500 2332 17172 2360
rect 15160 2320 15166 2332
rect 9539 2264 9628 2292
rect 9539 2261 9551 2264
rect 9493 2255 9551 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 11333 2295 11391 2301
rect 11333 2292 11345 2295
rect 9732 2264 11345 2292
rect 9732 2252 9738 2264
rect 11333 2261 11345 2264
rect 11379 2261 11391 2295
rect 11333 2255 11391 2261
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 12713 2295 12771 2301
rect 12713 2292 12725 2295
rect 12492 2264 12725 2292
rect 12492 2252 12498 2264
rect 12713 2261 12725 2264
rect 12759 2261 12771 2295
rect 12713 2255 12771 2261
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13228 2264 13645 2292
rect 13228 2252 13234 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 13998 2252 14004 2304
rect 14056 2292 14062 2304
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 14056 2264 15209 2292
rect 14056 2252 14062 2264
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15197 2255 15255 2261
rect 15470 2252 15476 2304
rect 15528 2252 15534 2304
rect 15764 2301 15792 2332
rect 17586 2320 17592 2372
rect 17644 2320 17650 2372
rect 18141 2363 18199 2369
rect 18141 2329 18153 2363
rect 18187 2360 18199 2363
rect 18506 2360 18512 2372
rect 18187 2332 18512 2360
rect 18187 2329 18199 2332
rect 18141 2323 18199 2329
rect 18506 2320 18512 2332
rect 18564 2320 18570 2372
rect 15749 2295 15807 2301
rect 15749 2261 15761 2295
rect 15795 2261 15807 2295
rect 15749 2255 15807 2261
rect 17034 2252 17040 2304
rect 17092 2252 17098 2304
rect 17126 2252 17132 2304
rect 17184 2292 17190 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17184 2264 17693 2292
rect 17184 2252 17190 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 18230 2252 18236 2304
rect 18288 2252 18294 2304
rect 18414 2252 18420 2304
rect 18472 2292 18478 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18472 2264 18797 2292
rect 18472 2252 18478 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 19352 2292 19380 2388
rect 19536 2372 19564 2400
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 21174 2428 21180 2440
rect 20671 2400 21180 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 21468 2428 21496 2536
rect 21836 2505 21864 2604
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 23198 2592 23204 2644
rect 23256 2592 23262 2644
rect 23308 2604 23888 2632
rect 21821 2499 21879 2505
rect 21821 2465 21833 2499
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 21468 2400 21680 2428
rect 19518 2320 19524 2372
rect 19576 2320 19582 2372
rect 20162 2320 20168 2372
rect 20220 2320 20226 2372
rect 21652 2360 21680 2400
rect 21726 2388 21732 2440
rect 21784 2388 21790 2440
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 23308 2428 23336 2604
rect 23566 2564 23572 2576
rect 23400 2536 23572 2564
rect 23400 2437 23428 2536
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 23860 2573 23888 2604
rect 23934 2592 23940 2644
rect 23992 2592 23998 2644
rect 23845 2567 23903 2573
rect 23845 2533 23857 2567
rect 23891 2533 23903 2567
rect 23845 2527 23903 2533
rect 23477 2499 23535 2505
rect 23477 2465 23489 2499
rect 23523 2496 23535 2499
rect 23952 2496 23980 2592
rect 23523 2468 23980 2496
rect 24029 2499 24087 2505
rect 23523 2465 23535 2468
rect 23477 2459 23535 2465
rect 24029 2465 24041 2499
rect 24075 2496 24087 2499
rect 24210 2496 24216 2508
rect 24075 2468 24216 2496
rect 24075 2465 24087 2468
rect 24029 2459 24087 2465
rect 24210 2456 24216 2468
rect 24268 2456 24274 2508
rect 21968 2400 23336 2428
rect 23385 2431 23443 2437
rect 21968 2388 21974 2400
rect 23385 2397 23397 2431
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 23566 2388 23572 2440
rect 23624 2388 23630 2440
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 23845 2431 23903 2437
rect 23845 2428 23857 2431
rect 23808 2400 23857 2428
rect 23808 2388 23814 2400
rect 23845 2397 23857 2400
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 22066 2363 22124 2369
rect 22066 2360 22078 2363
rect 21652 2332 22078 2360
rect 22066 2329 22078 2332
rect 22112 2329 22124 2363
rect 24213 2363 24271 2369
rect 22066 2323 22124 2329
rect 23124 2332 23612 2360
rect 21545 2295 21603 2301
rect 21545 2292 21557 2295
rect 19352 2264 21557 2292
rect 18785 2255 18843 2261
rect 21545 2261 21557 2264
rect 21591 2261 21603 2295
rect 21545 2255 21603 2261
rect 21634 2252 21640 2304
rect 21692 2292 21698 2304
rect 23124 2292 23152 2332
rect 21692 2264 23152 2292
rect 23584 2292 23612 2332
rect 24213 2329 24225 2363
rect 24259 2329 24271 2363
rect 24213 2323 24271 2329
rect 24228 2292 24256 2323
rect 23584 2264 24256 2292
rect 21692 2252 21698 2264
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 1581 2091 1639 2097
rect 1581 2057 1593 2091
rect 1627 2088 1639 2091
rect 1627 2060 2360 2088
rect 1627 2057 1639 2060
rect 1581 2051 1639 2057
rect 1946 1991 1952 2032
rect 1931 1985 1952 1991
rect 1394 1912 1400 1964
rect 1452 1912 1458 1964
rect 1670 1912 1676 1964
rect 1728 1912 1734 1964
rect 1931 1951 1943 1985
rect 2004 1980 2010 2032
rect 2332 2020 2360 2060
rect 2406 2048 2412 2100
rect 2464 2088 2470 2100
rect 2685 2091 2743 2097
rect 2685 2088 2697 2091
rect 2464 2060 2697 2088
rect 2464 2048 2470 2060
rect 2685 2057 2697 2060
rect 2731 2057 2743 2091
rect 2685 2051 2743 2057
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 4249 2091 4307 2097
rect 4249 2088 4261 2091
rect 4028 2060 4261 2088
rect 4028 2048 4034 2060
rect 4249 2057 4261 2060
rect 4295 2057 4307 2091
rect 4249 2051 4307 2057
rect 4982 2048 4988 2100
rect 5040 2048 5046 2100
rect 5258 2048 5264 2100
rect 5316 2048 5322 2100
rect 5350 2048 5356 2100
rect 5408 2048 5414 2100
rect 6454 2088 6460 2100
rect 5644 2060 6460 2088
rect 3326 2020 3332 2032
rect 2332 1992 3332 2020
rect 3326 1980 3332 1992
rect 3384 1980 3390 2032
rect 4614 2020 4620 2032
rect 3712 1992 4620 2020
rect 1977 1954 1992 1980
rect 1977 1951 1989 1954
rect 1931 1945 1989 1951
rect 3418 1912 3424 1964
rect 3476 1912 3482 1964
rect 3712 1961 3740 1992
rect 4614 1980 4620 1992
rect 4672 1980 4678 2032
rect 5276 2020 5304 2048
rect 5644 2029 5672 2060
rect 6454 2048 6460 2060
rect 6512 2048 6518 2100
rect 6638 2088 6644 2100
rect 6564 2060 6644 2088
rect 4816 1992 5304 2020
rect 5629 2023 5687 2029
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 3786 1912 3792 1964
rect 3844 1912 3850 1964
rect 4154 1912 4160 1964
rect 4212 1912 4218 1964
rect 4816 1961 4844 1992
rect 5629 1989 5641 2023
rect 5675 1989 5687 2023
rect 5629 1983 5687 1989
rect 5810 1980 5816 2032
rect 5868 1980 5874 2032
rect 5997 2023 6055 2029
rect 5997 1989 6009 2023
rect 6043 2020 6055 2023
rect 6564 2020 6592 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 6730 2048 6736 2100
rect 6788 2088 6794 2100
rect 6825 2091 6883 2097
rect 6825 2088 6837 2091
rect 6788 2060 6837 2088
rect 6788 2048 6794 2060
rect 6825 2057 6837 2060
rect 6871 2057 6883 2091
rect 7466 2088 7472 2100
rect 6825 2051 6883 2057
rect 7024 2060 7472 2088
rect 6043 1992 6592 2020
rect 6043 1989 6055 1992
rect 5997 1983 6055 1989
rect 4433 1955 4491 1961
rect 4433 1921 4445 1955
rect 4479 1952 4491 1955
rect 4801 1955 4859 1961
rect 4479 1924 4752 1952
rect 4479 1921 4491 1924
rect 4433 1915 4491 1921
rect 3510 1844 3516 1896
rect 3568 1884 3574 1896
rect 4724 1884 4752 1924
rect 4801 1921 4813 1955
rect 4847 1921 4859 1955
rect 4801 1915 4859 1921
rect 5074 1912 5080 1964
rect 5132 1952 5138 1964
rect 5261 1955 5319 1961
rect 5261 1952 5273 1955
rect 5132 1924 5273 1952
rect 5132 1912 5138 1924
rect 5261 1921 5273 1924
rect 5307 1921 5319 1955
rect 5261 1915 5319 1921
rect 6178 1912 6184 1964
rect 6236 1912 6242 1964
rect 6546 1912 6552 1964
rect 6604 1912 6610 1964
rect 6641 1955 6699 1961
rect 6641 1921 6653 1955
rect 6687 1952 6699 1955
rect 7024 1952 7052 2060
rect 7466 2048 7472 2060
rect 7524 2048 7530 2100
rect 7558 2048 7564 2100
rect 7616 2048 7622 2100
rect 8570 2088 8576 2100
rect 7668 2060 8576 2088
rect 7668 2020 7696 2060
rect 8570 2048 8576 2060
rect 8628 2048 8634 2100
rect 8938 2048 8944 2100
rect 8996 2048 9002 2100
rect 9125 2091 9183 2097
rect 9125 2057 9137 2091
rect 9171 2088 9183 2091
rect 9306 2088 9312 2100
rect 9171 2060 9312 2088
rect 9171 2057 9183 2060
rect 9125 2051 9183 2057
rect 9306 2048 9312 2060
rect 9364 2048 9370 2100
rect 10502 2048 10508 2100
rect 10560 2048 10566 2100
rect 11882 2048 11888 2100
rect 11940 2048 11946 2100
rect 13630 2048 13636 2100
rect 13688 2048 13694 2100
rect 13998 2048 14004 2100
rect 14056 2048 14062 2100
rect 15102 2048 15108 2100
rect 15160 2048 15166 2100
rect 15197 2091 15255 2097
rect 15197 2057 15209 2091
rect 15243 2057 15255 2091
rect 17770 2088 17776 2100
rect 15197 2051 15255 2057
rect 17328 2060 17776 2088
rect 8956 2020 8984 2048
rect 7116 1992 7696 2020
rect 7760 1992 8984 2020
rect 9692 1992 11100 2020
rect 7116 1961 7144 1992
rect 7484 1961 7604 1962
rect 6687 1924 7052 1952
rect 7101 1955 7159 1961
rect 6687 1921 6699 1924
rect 6641 1915 6699 1921
rect 7101 1921 7113 1955
rect 7147 1921 7159 1955
rect 7101 1915 7159 1921
rect 7469 1955 7604 1961
rect 7469 1921 7481 1955
rect 7515 1952 7604 1955
rect 7760 1952 7788 1992
rect 7515 1934 7788 1952
rect 7515 1921 7527 1934
rect 7576 1924 7788 1934
rect 7837 1955 7895 1961
rect 7469 1915 7527 1921
rect 7837 1921 7849 1955
rect 7883 1921 7895 1955
rect 7837 1915 7895 1921
rect 5902 1884 5908 1896
rect 3568 1856 4016 1884
rect 4724 1856 5908 1884
rect 3568 1844 3574 1856
rect 3988 1825 4016 1856
rect 5902 1844 5908 1856
rect 5960 1844 5966 1896
rect 7852 1884 7880 1915
rect 7926 1912 7932 1964
rect 7984 1952 7990 1964
rect 8021 1955 8079 1961
rect 8021 1952 8033 1955
rect 7984 1924 8033 1952
rect 7984 1912 7990 1924
rect 8021 1921 8033 1924
rect 8067 1921 8079 1955
rect 8021 1915 8079 1921
rect 8113 1955 8171 1961
rect 8113 1921 8125 1955
rect 8159 1952 8171 1955
rect 8294 1952 8300 1964
rect 8159 1924 8300 1952
rect 8159 1921 8171 1924
rect 8113 1915 8171 1921
rect 6380 1856 7880 1884
rect 6380 1825 6408 1856
rect 3973 1819 4031 1825
rect 3973 1785 3985 1819
rect 4019 1785 4031 1819
rect 6365 1819 6423 1825
rect 3973 1779 4031 1785
rect 4448 1788 5396 1816
rect 3237 1751 3295 1757
rect 3237 1717 3249 1751
rect 3283 1748 3295 1751
rect 3326 1748 3332 1760
rect 3283 1720 3332 1748
rect 3283 1717 3295 1720
rect 3237 1711 3295 1717
rect 3326 1708 3332 1720
rect 3384 1708 3390 1760
rect 3513 1751 3571 1757
rect 3513 1717 3525 1751
rect 3559 1748 3571 1751
rect 4448 1748 4476 1788
rect 3559 1720 4476 1748
rect 4617 1751 4675 1757
rect 3559 1717 3571 1720
rect 3513 1711 3571 1717
rect 4617 1717 4629 1751
rect 4663 1748 4675 1751
rect 5074 1748 5080 1760
rect 4663 1720 5080 1748
rect 4663 1717 4675 1720
rect 4617 1711 4675 1717
rect 5074 1708 5080 1720
rect 5132 1708 5138 1760
rect 5368 1748 5396 1788
rect 6365 1785 6377 1819
rect 6411 1785 6423 1819
rect 6365 1779 6423 1785
rect 7190 1776 7196 1828
rect 7248 1776 7254 1828
rect 7285 1819 7343 1825
rect 7285 1785 7297 1819
rect 7331 1816 7343 1819
rect 8018 1816 8024 1828
rect 7331 1788 8024 1816
rect 7331 1785 7343 1788
rect 7285 1779 7343 1785
rect 8018 1776 8024 1788
rect 8076 1776 8082 1828
rect 7208 1748 7236 1776
rect 5368 1720 7236 1748
rect 8128 1748 8156 1915
rect 8294 1912 8300 1924
rect 8352 1912 8358 1964
rect 8387 1955 8445 1961
rect 8387 1921 8399 1955
rect 8433 1952 8445 1955
rect 9692 1952 9720 1992
rect 8433 1924 9720 1952
rect 9767 1955 9825 1961
rect 8433 1921 8445 1924
rect 8387 1915 8445 1921
rect 9767 1921 9779 1955
rect 9813 1952 9825 1955
rect 10318 1952 10324 1964
rect 9813 1924 10324 1952
rect 9813 1921 9825 1924
rect 9767 1915 9825 1921
rect 10318 1912 10324 1924
rect 10376 1912 10382 1964
rect 10965 1955 11023 1961
rect 10965 1921 10977 1955
rect 11011 1921 11023 1955
rect 11072 1952 11100 1992
rect 11606 1980 11612 2032
rect 11664 2020 11670 2032
rect 11793 2023 11851 2029
rect 11793 2020 11805 2023
rect 11664 1992 11805 2020
rect 11664 1980 11670 1992
rect 11793 1989 11805 1992
rect 11839 1989 11851 2023
rect 11900 2020 11928 2048
rect 12345 2023 12403 2029
rect 12345 2020 12357 2023
rect 11900 1992 12357 2020
rect 11793 1983 11851 1989
rect 12345 1989 12357 1992
rect 12391 1989 12403 2023
rect 12345 1983 12403 1989
rect 12618 1952 12624 1964
rect 11072 1924 12624 1952
rect 10965 1915 11023 1921
rect 9493 1887 9551 1893
rect 9493 1853 9505 1887
rect 9539 1853 9551 1887
rect 10980 1884 11008 1915
rect 12618 1912 12624 1924
rect 12676 1912 12682 1964
rect 13081 1955 13139 1961
rect 13081 1921 13093 1955
rect 13127 1952 13139 1955
rect 13541 1955 13599 1961
rect 13541 1952 13553 1955
rect 13127 1924 13553 1952
rect 13127 1921 13139 1924
rect 13081 1915 13139 1921
rect 13541 1921 13553 1924
rect 13587 1952 13599 1955
rect 13648 1952 13676 2048
rect 13587 1924 13676 1952
rect 13587 1921 13599 1924
rect 13541 1915 13599 1921
rect 13814 1912 13820 1964
rect 13872 1912 13878 1964
rect 14016 1884 14044 2048
rect 15120 2020 15148 2048
rect 14476 1992 15148 2020
rect 14274 1912 14280 1964
rect 14332 1912 14338 1964
rect 14476 1961 14504 1992
rect 14461 1955 14519 1961
rect 14461 1921 14473 1955
rect 14507 1921 14519 1955
rect 14461 1915 14519 1921
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1952 14887 1955
rect 15212 1952 15240 2051
rect 15562 1980 15568 2032
rect 15620 2020 15626 2032
rect 17328 2029 17356 2060
rect 17770 2048 17776 2060
rect 17828 2048 17834 2100
rect 18325 2091 18383 2097
rect 18325 2057 18337 2091
rect 18371 2057 18383 2091
rect 18325 2051 18383 2057
rect 17313 2023 17371 2029
rect 15620 1992 16160 2020
rect 15620 1980 15626 1992
rect 16132 1961 16160 1992
rect 17313 1989 17325 2023
rect 17359 1989 17371 2023
rect 17313 1983 17371 1989
rect 17494 1980 17500 2032
rect 17552 2020 17558 2032
rect 17865 2023 17923 2029
rect 17865 2020 17877 2023
rect 17552 1992 17877 2020
rect 17552 1980 17558 1992
rect 17865 1989 17877 1992
rect 17911 1989 17923 2023
rect 17865 1983 17923 1989
rect 14875 1924 15240 1952
rect 15381 1955 15439 1961
rect 14875 1921 14887 1924
rect 14829 1915 14887 1921
rect 15381 1921 15393 1955
rect 15427 1921 15439 1955
rect 15381 1915 15439 1921
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1921 15715 1955
rect 15657 1915 15715 1921
rect 16117 1955 16175 1961
rect 16117 1921 16129 1955
rect 16163 1921 16175 1955
rect 16117 1915 16175 1921
rect 16761 1955 16819 1961
rect 16761 1921 16773 1955
rect 16807 1952 16819 1955
rect 18340 1952 18368 2051
rect 19426 2048 19432 2100
rect 19484 2048 19490 2100
rect 19610 2048 19616 2100
rect 19668 2088 19674 2100
rect 22002 2088 22008 2100
rect 19668 2060 22008 2088
rect 19668 2048 19674 2060
rect 22002 2048 22008 2060
rect 22060 2048 22066 2100
rect 22373 2091 22431 2097
rect 22373 2057 22385 2091
rect 22419 2088 22431 2091
rect 22462 2088 22468 2100
rect 22419 2060 22468 2088
rect 22419 2057 22431 2060
rect 22373 2051 22431 2057
rect 22462 2048 22468 2060
rect 22520 2048 22526 2100
rect 22922 2048 22928 2100
rect 22980 2088 22986 2100
rect 23934 2088 23940 2100
rect 22980 2060 23940 2088
rect 22980 2048 22986 2060
rect 23934 2048 23940 2060
rect 23992 2048 23998 2100
rect 16807 1924 18368 1952
rect 18509 1955 18567 1961
rect 16807 1921 16819 1924
rect 16761 1915 16819 1921
rect 18509 1921 18521 1955
rect 18555 1921 18567 1955
rect 18509 1915 18567 1921
rect 10980 1856 14044 1884
rect 9493 1847 9551 1853
rect 9508 1748 9536 1847
rect 15010 1844 15016 1896
rect 15068 1884 15074 1896
rect 15396 1884 15424 1915
rect 15068 1856 15424 1884
rect 15672 1884 15700 1915
rect 16298 1884 16304 1896
rect 15672 1856 16304 1884
rect 15068 1844 15074 1856
rect 16298 1844 16304 1856
rect 16356 1844 16362 1896
rect 16574 1844 16580 1896
rect 16632 1884 16638 1896
rect 18524 1884 18552 1915
rect 16632 1856 18552 1884
rect 18601 1887 18659 1893
rect 16632 1844 16638 1856
rect 18601 1853 18613 1887
rect 18647 1884 18659 1887
rect 18782 1884 18788 1896
rect 18647 1856 18788 1884
rect 18647 1853 18659 1856
rect 18601 1847 18659 1853
rect 18782 1844 18788 1856
rect 18840 1844 18846 1896
rect 18877 1887 18935 1893
rect 18877 1853 18889 1887
rect 18923 1853 18935 1887
rect 19444 1884 19472 2048
rect 21450 1980 21456 2032
rect 21508 1980 21514 2032
rect 22741 2023 22799 2029
rect 22741 2020 22753 2023
rect 21652 1992 22753 2020
rect 19705 1955 19763 1961
rect 19705 1921 19717 1955
rect 19751 1952 19763 1955
rect 20162 1952 20168 1964
rect 19751 1924 20168 1952
rect 19751 1921 19763 1924
rect 19705 1915 19763 1921
rect 20162 1912 20168 1924
rect 20220 1912 20226 1964
rect 20806 1912 20812 1964
rect 20864 1912 20870 1964
rect 21082 1912 21088 1964
rect 21140 1952 21146 1964
rect 21652 1952 21680 1992
rect 22741 1989 22753 1992
rect 22787 1989 22799 2023
rect 22741 1983 22799 1989
rect 24302 1980 24308 2032
rect 24360 1980 24366 2032
rect 21140 1924 21680 1952
rect 21913 1955 21971 1961
rect 21140 1912 21146 1924
rect 21913 1921 21925 1955
rect 21959 1952 21971 1955
rect 22189 1955 22247 1961
rect 21959 1924 22094 1952
rect 21959 1921 21971 1924
rect 21913 1915 21971 1921
rect 19889 1887 19947 1893
rect 19889 1884 19901 1887
rect 19444 1856 19901 1884
rect 18877 1847 18935 1853
rect 19889 1853 19901 1856
rect 19935 1853 19947 1887
rect 19889 1847 19947 1853
rect 13357 1819 13415 1825
rect 13357 1785 13369 1819
rect 13403 1816 13415 1819
rect 13998 1816 14004 1828
rect 13403 1788 14004 1816
rect 13403 1785 13415 1788
rect 13357 1779 13415 1785
rect 13998 1776 14004 1788
rect 14056 1776 14062 1828
rect 14093 1819 14151 1825
rect 14093 1785 14105 1819
rect 14139 1816 14151 1819
rect 15194 1816 15200 1828
rect 14139 1788 15200 1816
rect 14139 1785 14151 1788
rect 14093 1779 14151 1785
rect 15194 1776 15200 1788
rect 15252 1776 15258 1828
rect 15378 1776 15384 1828
rect 15436 1816 15442 1828
rect 15436 1788 16344 1816
rect 15436 1776 15442 1788
rect 8128 1720 9536 1748
rect 11054 1708 11060 1760
rect 11112 1708 11118 1760
rect 11882 1708 11888 1760
rect 11940 1708 11946 1760
rect 12618 1708 12624 1760
rect 12676 1708 12682 1760
rect 13630 1708 13636 1760
rect 13688 1708 13694 1760
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14645 1751 14703 1757
rect 14645 1748 14657 1751
rect 14332 1720 14657 1748
rect 14332 1708 14338 1720
rect 14645 1717 14657 1720
rect 14691 1717 14703 1751
rect 14645 1711 14703 1717
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14792 1720 15025 1748
rect 14792 1708 14798 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15654 1708 15660 1760
rect 15712 1748 15718 1760
rect 16316 1757 16344 1788
rect 18138 1776 18144 1828
rect 18196 1816 18202 1828
rect 18892 1816 18920 1847
rect 20254 1844 20260 1896
rect 20312 1884 20318 1896
rect 21634 1884 21640 1896
rect 20312 1856 21640 1884
rect 20312 1844 20318 1856
rect 21634 1844 21640 1856
rect 21692 1844 21698 1896
rect 22066 1884 22094 1924
rect 22189 1921 22201 1955
rect 22235 1952 22247 1955
rect 23106 1952 23112 1964
rect 22235 1924 23112 1952
rect 22235 1921 22247 1924
rect 22189 1915 22247 1921
rect 23106 1912 23112 1924
rect 23164 1912 23170 1964
rect 23658 1884 23664 1896
rect 22066 1856 23664 1884
rect 23658 1844 23664 1856
rect 23716 1844 23722 1896
rect 18196 1788 18920 1816
rect 18196 1776 18202 1788
rect 22830 1776 22836 1828
rect 22888 1816 22894 1828
rect 24486 1816 24492 1828
rect 22888 1788 24492 1816
rect 22888 1776 22894 1788
rect 24486 1776 24492 1788
rect 24544 1776 24550 1828
rect 15749 1751 15807 1757
rect 15749 1748 15761 1751
rect 15712 1720 15761 1748
rect 15712 1708 15718 1720
rect 15749 1717 15761 1720
rect 15795 1717 15807 1751
rect 15749 1711 15807 1717
rect 16301 1751 16359 1757
rect 16301 1717 16313 1751
rect 16347 1717 16359 1751
rect 16301 1711 16359 1717
rect 16850 1708 16856 1760
rect 16908 1708 16914 1760
rect 17402 1708 17408 1760
rect 17460 1708 17466 1760
rect 17586 1708 17592 1760
rect 17644 1748 17650 1760
rect 17957 1751 18015 1757
rect 17957 1748 17969 1751
rect 17644 1720 17969 1748
rect 17644 1708 17650 1720
rect 17957 1717 17969 1720
rect 18003 1717 18015 1751
rect 17957 1711 18015 1717
rect 19518 1708 19524 1760
rect 19576 1748 19582 1760
rect 21634 1748 21640 1760
rect 19576 1720 21640 1748
rect 19576 1708 19582 1720
rect 21634 1708 21640 1720
rect 21692 1708 21698 1760
rect 22005 1751 22063 1757
rect 22005 1717 22017 1751
rect 22051 1748 22063 1751
rect 25314 1748 25320 1760
rect 22051 1720 25320 1748
rect 22051 1717 22063 1720
rect 22005 1711 22063 1717
rect 25314 1708 25320 1720
rect 25372 1708 25378 1760
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 2774 1504 2780 1556
rect 2832 1504 2838 1556
rect 4157 1547 4215 1553
rect 4157 1513 4169 1547
rect 4203 1544 4215 1547
rect 4890 1544 4896 1556
rect 4203 1516 4896 1544
rect 4203 1513 4215 1516
rect 4157 1507 4215 1513
rect 4890 1504 4896 1516
rect 4948 1504 4954 1556
rect 6546 1504 6552 1556
rect 6604 1544 6610 1556
rect 9306 1544 9312 1556
rect 6604 1516 9312 1544
rect 6604 1504 6610 1516
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 10686 1504 10692 1556
rect 10744 1504 10750 1556
rect 13170 1544 13176 1556
rect 11808 1516 13176 1544
rect 3326 1436 3332 1488
rect 3384 1476 3390 1488
rect 8846 1476 8852 1488
rect 3384 1448 8852 1476
rect 3384 1436 3390 1448
rect 8846 1436 8852 1448
rect 8904 1436 8910 1488
rect 8941 1479 8999 1485
rect 8941 1445 8953 1479
rect 8987 1445 8999 1479
rect 8941 1439 8999 1445
rect 566 1368 572 1420
rect 624 1408 630 1420
rect 624 1380 1992 1408
rect 624 1368 630 1380
rect 1394 1300 1400 1352
rect 1452 1300 1458 1352
rect 1670 1300 1676 1352
rect 1728 1300 1734 1352
rect 1578 1164 1584 1216
rect 1636 1164 1642 1216
rect 1854 1164 1860 1216
rect 1912 1164 1918 1216
rect 1964 1204 1992 1380
rect 3786 1368 3792 1420
rect 3844 1408 3850 1420
rect 4706 1408 4712 1420
rect 3844 1380 4712 1408
rect 3844 1368 3850 1380
rect 4706 1368 4712 1380
rect 4764 1368 4770 1420
rect 2038 1300 2044 1352
rect 2096 1340 2102 1352
rect 4893 1343 4951 1349
rect 2096 1312 2728 1340
rect 2096 1300 2102 1312
rect 2314 1232 2320 1284
rect 2372 1232 2378 1284
rect 2498 1232 2504 1284
rect 2556 1232 2562 1284
rect 2700 1281 2728 1312
rect 2976 1312 3648 1340
rect 2685 1275 2743 1281
rect 2685 1241 2697 1275
rect 2731 1241 2743 1275
rect 2685 1235 2743 1241
rect 2976 1204 3004 1312
rect 3050 1232 3056 1284
rect 3108 1232 3114 1284
rect 3620 1281 3648 1312
rect 4893 1309 4905 1343
rect 4939 1340 4951 1343
rect 4939 1312 5212 1340
rect 4939 1309 4951 1312
rect 4893 1303 4951 1309
rect 3421 1275 3479 1281
rect 3421 1241 3433 1275
rect 3467 1241 3479 1275
rect 3421 1235 3479 1241
rect 3605 1275 3663 1281
rect 3605 1241 3617 1275
rect 3651 1241 3663 1275
rect 3605 1235 3663 1241
rect 1964 1176 3004 1204
rect 3142 1164 3148 1216
rect 3200 1164 3206 1216
rect 3436 1204 3464 1235
rect 3878 1232 3884 1284
rect 3936 1232 3942 1284
rect 4430 1232 4436 1284
rect 4488 1272 4494 1284
rect 4617 1275 4675 1281
rect 4617 1272 4629 1275
rect 4488 1244 4629 1272
rect 4488 1232 4494 1244
rect 4617 1241 4629 1244
rect 4663 1241 4675 1275
rect 4617 1235 4675 1241
rect 3786 1204 3792 1216
rect 3436 1176 3792 1204
rect 3786 1164 3792 1176
rect 3844 1164 3850 1216
rect 4709 1207 4767 1213
rect 4709 1173 4721 1207
rect 4755 1204 4767 1207
rect 4982 1204 4988 1216
rect 4755 1176 4988 1204
rect 4755 1173 4767 1176
rect 4709 1167 4767 1173
rect 4982 1164 4988 1176
rect 5040 1164 5046 1216
rect 5074 1164 5080 1216
rect 5132 1164 5138 1216
rect 5184 1204 5212 1312
rect 5258 1300 5264 1352
rect 5316 1300 5322 1352
rect 5534 1300 5540 1352
rect 5592 1300 5598 1352
rect 6362 1300 6368 1352
rect 6420 1340 6426 1352
rect 6549 1343 6607 1349
rect 6549 1340 6561 1343
rect 6420 1312 6561 1340
rect 6420 1300 6426 1312
rect 6549 1309 6561 1312
rect 6595 1309 6607 1343
rect 7377 1343 7435 1349
rect 7377 1340 7389 1343
rect 6549 1303 6607 1309
rect 6656 1312 7389 1340
rect 6656 1272 6684 1312
rect 7377 1309 7389 1312
rect 7423 1309 7435 1343
rect 7377 1303 7435 1309
rect 7745 1343 7803 1349
rect 7745 1309 7757 1343
rect 7791 1340 7803 1343
rect 8018 1340 8024 1352
rect 7791 1312 8024 1340
rect 7791 1309 7803 1312
rect 7745 1303 7803 1309
rect 8018 1300 8024 1312
rect 8076 1300 8082 1352
rect 8113 1343 8171 1349
rect 8113 1309 8125 1343
rect 8159 1309 8171 1343
rect 8113 1303 8171 1309
rect 8481 1343 8539 1349
rect 8481 1309 8493 1343
rect 8527 1340 8539 1343
rect 8956 1340 8984 1439
rect 9030 1436 9036 1488
rect 9088 1476 9094 1488
rect 10704 1476 10732 1504
rect 9088 1448 10732 1476
rect 9088 1436 9094 1448
rect 9950 1368 9956 1420
rect 10008 1368 10014 1420
rect 11238 1368 11244 1420
rect 11296 1368 11302 1420
rect 8527 1312 8984 1340
rect 8527 1309 8539 1312
rect 8481 1303 8539 1309
rect 6380 1244 6684 1272
rect 6270 1204 6276 1216
rect 5184 1176 6276 1204
rect 6270 1164 6276 1176
rect 6328 1164 6334 1216
rect 6380 1213 6408 1244
rect 6730 1232 6736 1284
rect 6788 1232 6794 1284
rect 6917 1275 6975 1281
rect 6917 1241 6929 1275
rect 6963 1272 6975 1275
rect 7006 1272 7012 1284
rect 6963 1244 7012 1272
rect 6963 1241 6975 1244
rect 6917 1235 6975 1241
rect 7006 1232 7012 1244
rect 7064 1232 7070 1284
rect 7101 1275 7159 1281
rect 7101 1241 7113 1275
rect 7147 1272 7159 1275
rect 8128 1272 8156 1303
rect 9030 1300 9036 1352
rect 9088 1340 9094 1352
rect 9125 1343 9183 1349
rect 9125 1340 9137 1343
rect 9088 1312 9137 1340
rect 9088 1300 9094 1312
rect 9125 1309 9137 1312
rect 9171 1340 9183 1343
rect 9401 1343 9459 1349
rect 9401 1340 9413 1343
rect 9171 1312 9413 1340
rect 9171 1309 9183 1312
rect 9125 1303 9183 1309
rect 9401 1309 9413 1312
rect 9447 1309 9459 1343
rect 9401 1303 9459 1309
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 10413 1343 10471 1349
rect 10413 1340 10425 1343
rect 9876 1312 10425 1340
rect 7147 1244 7788 1272
rect 8128 1244 9168 1272
rect 7147 1241 7159 1244
rect 7101 1235 7159 1241
rect 7760 1216 7788 1244
rect 6365 1207 6423 1213
rect 6365 1173 6377 1207
rect 6411 1173 6423 1207
rect 6365 1167 6423 1173
rect 6454 1164 6460 1216
rect 6512 1204 6518 1216
rect 7193 1207 7251 1213
rect 7193 1204 7205 1207
rect 6512 1176 7205 1204
rect 6512 1164 6518 1176
rect 7193 1173 7205 1176
rect 7239 1173 7251 1207
rect 7193 1167 7251 1173
rect 7558 1164 7564 1216
rect 7616 1164 7622 1216
rect 7742 1164 7748 1216
rect 7800 1164 7806 1216
rect 7926 1164 7932 1216
rect 7984 1164 7990 1216
rect 8294 1164 8300 1216
rect 8352 1164 8358 1216
rect 8662 1164 8668 1216
rect 8720 1164 8726 1216
rect 9140 1204 9168 1244
rect 9214 1232 9220 1284
rect 9272 1272 9278 1284
rect 9876 1272 9904 1312
rect 10413 1309 10425 1312
rect 10459 1309 10471 1343
rect 10413 1303 10471 1309
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1340 11023 1343
rect 11011 1312 11652 1340
rect 11011 1309 11023 1312
rect 10965 1303 11023 1309
rect 11330 1272 11336 1284
rect 9272 1244 9904 1272
rect 10428 1244 11336 1272
rect 9272 1232 9278 1244
rect 10428 1204 10456 1244
rect 11330 1232 11336 1244
rect 11388 1232 11394 1284
rect 11624 1272 11652 1312
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11808 1349 11836 1516
rect 13170 1504 13176 1516
rect 13228 1504 13234 1556
rect 13814 1504 13820 1556
rect 13872 1544 13878 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13872 1516 14289 1544
rect 13872 1504 13878 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 14918 1504 14924 1556
rect 14976 1544 14982 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 14976 1516 15393 1544
rect 14976 1504 14982 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 13633 1479 13691 1485
rect 13633 1476 13645 1479
rect 12268 1448 13645 1476
rect 12268 1408 12296 1448
rect 13633 1445 13645 1448
rect 13679 1445 13691 1479
rect 13633 1439 13691 1445
rect 15102 1436 15108 1488
rect 15160 1476 15166 1488
rect 15948 1476 15976 1507
rect 16298 1504 16304 1556
rect 16356 1504 16362 1556
rect 16390 1504 16396 1556
rect 16448 1544 16454 1556
rect 16853 1547 16911 1553
rect 16853 1544 16865 1547
rect 16448 1516 16865 1544
rect 16448 1504 16454 1516
rect 16853 1513 16865 1516
rect 16899 1513 16911 1547
rect 16853 1507 16911 1513
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1513 17463 1547
rect 17405 1507 17463 1513
rect 15160 1448 15976 1476
rect 15160 1436 15166 1448
rect 16574 1436 16580 1488
rect 16632 1476 16638 1488
rect 17420 1476 17448 1507
rect 17954 1504 17960 1556
rect 18012 1544 18018 1556
rect 18509 1547 18567 1553
rect 18509 1544 18521 1547
rect 18012 1516 18521 1544
rect 18012 1504 18018 1516
rect 18509 1513 18521 1516
rect 18555 1513 18567 1547
rect 18509 1507 18567 1513
rect 18782 1504 18788 1556
rect 18840 1544 18846 1556
rect 18840 1516 22094 1544
rect 18840 1504 18846 1516
rect 16632 1448 17448 1476
rect 18049 1479 18107 1485
rect 16632 1436 16638 1448
rect 18049 1445 18061 1479
rect 18095 1445 18107 1479
rect 18877 1479 18935 1485
rect 18877 1476 18889 1479
rect 18049 1439 18107 1445
rect 18524 1448 18889 1476
rect 11900 1380 12296 1408
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1309 11851 1343
rect 11793 1303 11851 1309
rect 11900 1272 11928 1380
rect 12342 1368 12348 1420
rect 12400 1408 12406 1420
rect 12529 1411 12587 1417
rect 12529 1408 12541 1411
rect 12400 1380 12541 1408
rect 12400 1368 12406 1380
rect 12529 1377 12541 1380
rect 12575 1377 12587 1411
rect 12529 1371 12587 1377
rect 13538 1368 13544 1420
rect 13596 1408 13602 1420
rect 13596 1380 13768 1408
rect 13596 1368 13602 1380
rect 12710 1340 12716 1352
rect 11624 1244 11928 1272
rect 11992 1312 12716 1340
rect 9140 1176 10456 1204
rect 10502 1164 10508 1216
rect 10560 1164 10566 1216
rect 11517 1207 11575 1213
rect 11517 1173 11529 1207
rect 11563 1204 11575 1207
rect 11882 1204 11888 1216
rect 11563 1176 11888 1204
rect 11563 1173 11575 1176
rect 11517 1167 11575 1173
rect 11882 1164 11888 1176
rect 11940 1164 11946 1216
rect 11992 1213 12020 1312
rect 12710 1300 12716 1312
rect 12768 1300 12774 1352
rect 12897 1343 12955 1349
rect 12897 1309 12909 1343
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 13265 1343 13323 1349
rect 13265 1309 13277 1343
rect 13311 1340 13323 1343
rect 13630 1340 13636 1352
rect 13311 1312 13636 1340
rect 13311 1309 13323 1312
rect 13265 1303 13323 1309
rect 12158 1232 12164 1284
rect 12216 1272 12222 1284
rect 12253 1275 12311 1281
rect 12253 1272 12265 1275
rect 12216 1244 12265 1272
rect 12216 1232 12222 1244
rect 12253 1241 12265 1244
rect 12299 1241 12311 1275
rect 12253 1235 12311 1241
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1173 12035 1207
rect 11977 1167 12035 1173
rect 12066 1164 12072 1216
rect 12124 1204 12130 1216
rect 12912 1204 12940 1303
rect 13630 1300 13636 1312
rect 13688 1300 13694 1352
rect 13740 1340 13768 1380
rect 16666 1368 16672 1420
rect 16724 1408 16730 1420
rect 18064 1408 18092 1439
rect 18524 1420 18552 1448
rect 18877 1445 18889 1448
rect 18923 1445 18935 1479
rect 18877 1439 18935 1445
rect 20530 1436 20536 1488
rect 20588 1436 20594 1488
rect 22066 1476 22094 1516
rect 22554 1504 22560 1556
rect 22612 1544 22618 1556
rect 23109 1547 23167 1553
rect 23109 1544 23121 1547
rect 22612 1516 23121 1544
rect 22612 1504 22618 1516
rect 23109 1513 23121 1516
rect 23155 1513 23167 1547
rect 23109 1507 23167 1513
rect 23842 1504 23848 1556
rect 23900 1504 23906 1556
rect 25314 1476 25320 1488
rect 22066 1448 25320 1476
rect 25314 1436 25320 1448
rect 25372 1436 25378 1488
rect 16724 1380 18092 1408
rect 16724 1368 16730 1380
rect 18506 1368 18512 1420
rect 18564 1368 18570 1420
rect 21174 1368 21180 1420
rect 21232 1408 21238 1420
rect 22830 1408 22836 1420
rect 21232 1380 22836 1408
rect 21232 1368 21238 1380
rect 22830 1368 22836 1380
rect 22888 1368 22894 1420
rect 23768 1380 24072 1408
rect 13817 1343 13875 1349
rect 13817 1340 13829 1343
rect 13740 1312 13829 1340
rect 13817 1309 13829 1312
rect 13863 1309 13875 1343
rect 13817 1303 13875 1309
rect 13906 1300 13912 1352
rect 13964 1300 13970 1352
rect 13998 1300 14004 1352
rect 14056 1340 14062 1352
rect 14645 1343 14703 1349
rect 14645 1340 14657 1343
rect 14056 1312 14657 1340
rect 14056 1300 14062 1312
rect 14645 1309 14657 1312
rect 14691 1309 14703 1343
rect 14645 1303 14703 1309
rect 15194 1300 15200 1352
rect 15252 1340 15258 1352
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 15252 1312 15301 1340
rect 15252 1300 15258 1312
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 15470 1300 15476 1352
rect 15528 1340 15534 1352
rect 15841 1343 15899 1349
rect 15841 1340 15853 1343
rect 15528 1312 15853 1340
rect 15528 1300 15534 1312
rect 15841 1309 15853 1312
rect 15887 1309 15899 1343
rect 15841 1303 15899 1309
rect 16482 1300 16488 1352
rect 16540 1300 16546 1352
rect 16761 1343 16819 1349
rect 16761 1309 16773 1343
rect 16807 1340 16819 1343
rect 17034 1340 17040 1352
rect 16807 1312 17040 1340
rect 16807 1309 16819 1312
rect 16761 1303 16819 1309
rect 17034 1300 17040 1312
rect 17092 1300 17098 1352
rect 17218 1300 17224 1352
rect 17276 1340 17282 1352
rect 17313 1343 17371 1349
rect 17313 1340 17325 1343
rect 17276 1312 17325 1340
rect 17276 1300 17282 1312
rect 17313 1309 17325 1312
rect 17359 1309 17371 1343
rect 17313 1303 17371 1309
rect 17494 1300 17500 1352
rect 17552 1340 17558 1352
rect 17865 1343 17923 1349
rect 17865 1340 17877 1343
rect 17552 1312 17877 1340
rect 17552 1300 17558 1312
rect 17865 1309 17877 1312
rect 17911 1309 17923 1343
rect 17865 1303 17923 1309
rect 18322 1300 18328 1352
rect 18380 1340 18386 1352
rect 18417 1343 18475 1349
rect 18417 1340 18429 1343
rect 18380 1312 18429 1340
rect 18380 1300 18386 1312
rect 18417 1309 18429 1312
rect 18463 1309 18475 1343
rect 18417 1303 18475 1309
rect 19058 1300 19064 1352
rect 19116 1300 19122 1352
rect 20622 1300 20628 1352
rect 20680 1340 20686 1352
rect 20680 1312 21496 1340
rect 20680 1300 20686 1312
rect 13924 1272 13952 1300
rect 14185 1275 14243 1281
rect 14185 1272 14197 1275
rect 13924 1244 14197 1272
rect 14185 1241 14197 1244
rect 14231 1241 14243 1275
rect 14185 1235 14243 1241
rect 17678 1232 17684 1284
rect 17736 1232 17742 1284
rect 19245 1275 19303 1281
rect 19245 1241 19257 1275
rect 19291 1272 19303 1275
rect 21082 1272 21088 1284
rect 19291 1244 21088 1272
rect 19291 1241 19303 1244
rect 19245 1235 19303 1241
rect 21082 1232 21088 1244
rect 21140 1232 21146 1284
rect 21174 1232 21180 1284
rect 21232 1232 21238 1284
rect 21358 1232 21364 1284
rect 21416 1232 21422 1284
rect 21468 1272 21496 1312
rect 21634 1300 21640 1352
rect 21692 1300 21698 1352
rect 23382 1300 23388 1352
rect 23440 1340 23446 1352
rect 23661 1343 23719 1349
rect 23661 1340 23673 1343
rect 23440 1312 23673 1340
rect 23440 1300 23446 1312
rect 23661 1309 23673 1312
rect 23707 1309 23719 1343
rect 23661 1303 23719 1309
rect 21821 1275 21879 1281
rect 21821 1272 21833 1275
rect 21468 1244 21833 1272
rect 21821 1241 21833 1244
rect 21867 1241 21879 1275
rect 21821 1235 21879 1241
rect 22186 1232 22192 1284
rect 22244 1272 22250 1284
rect 23768 1272 23796 1380
rect 23934 1300 23940 1352
rect 23992 1300 23998 1352
rect 24044 1340 24072 1380
rect 24121 1343 24179 1349
rect 24121 1340 24133 1343
rect 24044 1312 24133 1340
rect 24121 1309 24133 1312
rect 24167 1309 24179 1343
rect 24121 1303 24179 1309
rect 22244 1244 23796 1272
rect 22244 1232 22250 1244
rect 12124 1176 12940 1204
rect 12124 1164 12130 1176
rect 13078 1164 13084 1216
rect 13136 1164 13142 1216
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13998 1164 14004 1216
rect 14056 1204 14062 1216
rect 14829 1207 14887 1213
rect 14829 1204 14841 1207
rect 14056 1176 14841 1204
rect 14056 1164 14062 1176
rect 14829 1173 14841 1176
rect 14875 1173 14887 1207
rect 17696 1204 17724 1232
rect 21453 1207 21511 1213
rect 21453 1204 21465 1207
rect 17696 1176 21465 1204
rect 14829 1167 14887 1173
rect 21453 1173 21465 1176
rect 21499 1173 21511 1207
rect 21453 1167 21511 1173
rect 23290 1164 23296 1216
rect 23348 1204 23354 1216
rect 23934 1204 23940 1216
rect 23348 1176 23940 1204
rect 23348 1164 23354 1176
rect 23934 1164 23940 1176
rect 23992 1164 23998 1216
rect 24118 1164 24124 1216
rect 24176 1164 24182 1216
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 934 960 940 1012
rect 992 1000 998 1012
rect 3878 1000 3884 1012
rect 992 972 3884 1000
rect 992 960 998 972
rect 3878 960 3884 972
rect 3936 960 3942 1012
rect 5810 960 5816 1012
rect 5868 1000 5874 1012
rect 6730 1000 6736 1012
rect 5868 972 6736 1000
rect 5868 960 5874 972
rect 6730 960 6736 972
rect 6788 960 6794 1012
rect 7926 960 7932 1012
rect 7984 1000 7990 1012
rect 10686 1000 10692 1012
rect 7984 972 10692 1000
rect 7984 960 7990 972
rect 10686 960 10692 972
rect 10744 960 10750 1012
rect 11698 960 11704 1012
rect 11756 1000 11762 1012
rect 13354 1000 13360 1012
rect 11756 972 13360 1000
rect 11756 960 11762 972
rect 13354 960 13360 972
rect 13412 960 13418 1012
rect 18046 960 18052 1012
rect 18104 1000 18110 1012
rect 20714 1000 20720 1012
rect 18104 972 20720 1000
rect 18104 960 18110 972
rect 20714 960 20720 972
rect 20772 960 20778 1012
rect 21174 960 21180 1012
rect 21232 1000 21238 1012
rect 21232 972 22094 1000
rect 21232 960 21238 972
rect 1578 892 1584 944
rect 1636 932 1642 944
rect 4338 932 4344 944
rect 1636 904 4344 932
rect 1636 892 1642 904
rect 4338 892 4344 904
rect 4396 892 4402 944
rect 5166 892 5172 944
rect 5224 932 5230 944
rect 6914 932 6920 944
rect 5224 904 6920 932
rect 5224 892 5230 904
rect 6914 892 6920 904
rect 6972 892 6978 944
rect 8018 892 8024 944
rect 8076 892 8082 944
rect 8294 892 8300 944
rect 8352 932 8358 944
rect 11514 932 11520 944
rect 8352 904 11520 932
rect 8352 892 8358 904
rect 11514 892 11520 904
rect 11572 892 11578 944
rect 22066 932 22094 972
rect 25590 932 25596 944
rect 22066 904 25596 932
rect 25590 892 25596 904
rect 25648 892 25654 944
rect 3142 824 3148 876
rect 3200 824 3206 876
rect 1394 688 1400 740
rect 1452 728 1458 740
rect 2406 728 2412 740
rect 1452 700 2412 728
rect 1452 688 1458 700
rect 2406 688 2412 700
rect 2464 688 2470 740
rect 3160 728 3188 824
rect 8036 796 8064 892
rect 8662 824 8668 876
rect 8720 864 8726 876
rect 12066 864 12072 876
rect 8720 836 12072 864
rect 8720 824 8726 836
rect 12066 824 12072 836
rect 12124 824 12130 876
rect 12434 796 12440 808
rect 8036 768 12440 796
rect 12434 756 12440 768
rect 12492 756 12498 808
rect 11146 728 11152 740
rect 3160 700 11152 728
rect 11146 688 11152 700
rect 11204 688 11210 740
rect 4430 620 4436 672
rect 4488 660 4494 672
rect 5534 660 5540 672
rect 4488 632 5540 660
rect 4488 620 4494 632
rect 5534 620 5540 632
rect 5592 620 5598 672
rect 6362 620 6368 672
rect 6420 660 6426 672
rect 9858 660 9864 672
rect 6420 632 9864 660
rect 6420 620 6426 632
rect 9858 620 9864 632
rect 9916 620 9922 672
rect 21082 620 21088 672
rect 21140 660 21146 672
rect 22002 660 22008 672
rect 21140 632 22008 660
rect 21140 620 21146 632
rect 22002 620 22008 632
rect 22060 620 22066 672
rect 7282 552 7288 604
rect 7340 592 7346 604
rect 14366 592 14372 604
rect 7340 564 14372 592
rect 7340 552 7346 564
rect 14366 552 14372 564
rect 14424 552 14430 604
rect 4982 484 4988 536
rect 5040 524 5046 536
rect 12250 524 12256 536
rect 5040 496 12256 524
rect 5040 484 5046 496
rect 12250 484 12256 496
rect 12308 484 12314 536
<< via1 >>
rect 18144 43800 18196 43852
rect 21272 43800 21324 43852
rect 21732 43800 21784 43852
rect 22928 43800 22980 43852
rect 20720 43732 20772 43784
rect 22560 43732 22612 43784
rect 5264 43664 5316 43716
rect 16028 43664 16080 43716
rect 18512 43664 18564 43716
rect 20996 43664 21048 43716
rect 3608 43596 3660 43648
rect 10508 43596 10560 43648
rect 17500 43596 17552 43648
rect 22376 43596 22428 43648
rect 6884 43494 6936 43546
rect 6948 43494 7000 43546
rect 7012 43494 7064 43546
rect 7076 43494 7128 43546
rect 7140 43494 7192 43546
rect 12818 43494 12870 43546
rect 12882 43494 12934 43546
rect 12946 43494 12998 43546
rect 13010 43494 13062 43546
rect 13074 43494 13126 43546
rect 18752 43494 18804 43546
rect 18816 43494 18868 43546
rect 18880 43494 18932 43546
rect 18944 43494 18996 43546
rect 19008 43494 19060 43546
rect 24686 43494 24738 43546
rect 24750 43494 24802 43546
rect 24814 43494 24866 43546
rect 24878 43494 24930 43546
rect 24942 43494 24994 43546
rect 1860 43435 1912 43444
rect 1860 43401 1869 43435
rect 1869 43401 1903 43435
rect 1903 43401 1912 43435
rect 1860 43392 1912 43401
rect 2964 43392 3016 43444
rect 388 43324 440 43376
rect 4344 43392 4396 43444
rect 5540 43435 5592 43444
rect 5540 43401 5549 43435
rect 5549 43401 5583 43435
rect 5583 43401 5592 43435
rect 5540 43392 5592 43401
rect 6276 43392 6328 43444
rect 6644 43392 6696 43444
rect 7656 43392 7708 43444
rect 7932 43392 7984 43444
rect 8484 43392 8536 43444
rect 9036 43392 9088 43444
rect 9588 43392 9640 43444
rect 9864 43392 9916 43444
rect 10508 43435 10560 43444
rect 10508 43401 10517 43435
rect 10517 43401 10551 43435
rect 10551 43401 10560 43435
rect 10508 43392 10560 43401
rect 14004 43392 14056 43444
rect 17040 43392 17092 43444
rect 664 43256 716 43308
rect 2504 43299 2556 43308
rect 2504 43265 2513 43299
rect 2513 43265 2547 43299
rect 2547 43265 2556 43299
rect 2504 43256 2556 43265
rect 4344 43256 4396 43308
rect 2964 43188 3016 43240
rect 4252 43188 4304 43240
rect 5448 43256 5500 43308
rect 5540 43256 5592 43308
rect 4712 43120 4764 43172
rect 1768 43052 1820 43104
rect 4436 43052 4488 43104
rect 8944 43324 8996 43376
rect 9404 43324 9456 43376
rect 11152 43324 11204 43376
rect 12440 43367 12492 43376
rect 12440 43333 12449 43367
rect 12449 43333 12483 43367
rect 12483 43333 12492 43367
rect 12440 43324 12492 43333
rect 12808 43367 12860 43376
rect 12808 43333 12817 43367
rect 12817 43333 12851 43367
rect 12851 43333 12860 43367
rect 12808 43324 12860 43333
rect 13360 43324 13412 43376
rect 14740 43367 14792 43376
rect 14740 43333 14749 43367
rect 14749 43333 14783 43367
rect 14783 43333 14792 43367
rect 14740 43324 14792 43333
rect 14832 43324 14884 43376
rect 15936 43324 15988 43376
rect 16396 43324 16448 43376
rect 16856 43324 16908 43376
rect 6276 43256 6328 43308
rect 7288 43256 7340 43308
rect 8116 43188 8168 43240
rect 9496 43299 9548 43308
rect 9496 43265 9505 43299
rect 9505 43265 9539 43299
rect 9539 43265 9548 43299
rect 9496 43256 9548 43265
rect 9956 43299 10008 43308
rect 9956 43265 9965 43299
rect 9965 43265 9999 43299
rect 9999 43265 10008 43299
rect 9956 43256 10008 43265
rect 10324 43299 10376 43308
rect 10324 43265 10333 43299
rect 10333 43265 10367 43299
rect 10367 43265 10376 43299
rect 10324 43256 10376 43265
rect 10692 43299 10744 43308
rect 10692 43265 10701 43299
rect 10701 43265 10735 43299
rect 10735 43265 10744 43299
rect 10692 43256 10744 43265
rect 11060 43299 11112 43308
rect 11060 43265 11069 43299
rect 11069 43265 11103 43299
rect 11103 43265 11112 43299
rect 11060 43256 11112 43265
rect 11244 43256 11296 43308
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 13636 43299 13688 43308
rect 13636 43265 13645 43299
rect 13645 43265 13679 43299
rect 13679 43265 13688 43299
rect 13636 43256 13688 43265
rect 15476 43299 15528 43308
rect 15476 43265 15485 43299
rect 15485 43265 15519 43299
rect 15519 43265 15528 43299
rect 15476 43256 15528 43265
rect 15844 43299 15896 43308
rect 15844 43265 15853 43299
rect 15853 43265 15887 43299
rect 15887 43265 15896 43299
rect 15844 43256 15896 43265
rect 16028 43256 16080 43308
rect 17408 43256 17460 43308
rect 18144 43392 18196 43444
rect 18236 43324 18288 43376
rect 9680 43188 9732 43240
rect 17316 43188 17368 43240
rect 19340 43256 19392 43308
rect 20352 43392 20404 43444
rect 20628 43392 20680 43444
rect 21180 43392 21232 43444
rect 20536 43324 20588 43376
rect 19892 43299 19944 43308
rect 19892 43265 19901 43299
rect 19901 43265 19935 43299
rect 19935 43265 19944 43299
rect 19892 43256 19944 43265
rect 19984 43188 20036 43240
rect 20628 43256 20680 43308
rect 21548 43324 21600 43376
rect 22928 43435 22980 43444
rect 22928 43401 22937 43435
rect 22937 43401 22971 43435
rect 22971 43401 22980 43435
rect 22928 43392 22980 43401
rect 23112 43392 23164 43444
rect 21640 43256 21692 43308
rect 23020 43324 23072 43376
rect 22468 43256 22520 43308
rect 22928 43256 22980 43308
rect 22192 43188 22244 43240
rect 22652 43188 22704 43240
rect 10600 43120 10652 43172
rect 13636 43120 13688 43172
rect 9772 43052 9824 43104
rect 10140 43095 10192 43104
rect 10140 43061 10149 43095
rect 10149 43061 10183 43095
rect 10183 43061 10192 43095
rect 10140 43052 10192 43061
rect 10968 43052 11020 43104
rect 11244 43095 11296 43104
rect 11244 43061 11253 43095
rect 11253 43061 11287 43095
rect 11287 43061 11296 43095
rect 11244 43052 11296 43061
rect 11980 43052 12032 43104
rect 12532 43095 12584 43104
rect 12532 43061 12541 43095
rect 12541 43061 12575 43095
rect 12575 43061 12584 43095
rect 12532 43052 12584 43061
rect 12900 43095 12952 43104
rect 12900 43061 12909 43095
rect 12909 43061 12943 43095
rect 12943 43061 12952 43095
rect 12900 43052 12952 43061
rect 14188 43052 14240 43104
rect 14280 43095 14332 43104
rect 14280 43061 14289 43095
rect 14289 43061 14323 43095
rect 14323 43061 14332 43095
rect 14280 43052 14332 43061
rect 14924 43163 14976 43172
rect 14924 43129 14933 43163
rect 14933 43129 14967 43163
rect 14967 43129 14976 43163
rect 14924 43120 14976 43129
rect 18328 43120 18380 43172
rect 20720 43120 20772 43172
rect 20904 43120 20956 43172
rect 15292 43052 15344 43104
rect 15844 43052 15896 43104
rect 16856 43095 16908 43104
rect 16856 43061 16865 43095
rect 16865 43061 16899 43095
rect 16899 43061 16908 43095
rect 16856 43052 16908 43061
rect 17500 43052 17552 43104
rect 17592 43095 17644 43104
rect 17592 43061 17601 43095
rect 17601 43061 17635 43095
rect 17635 43061 17644 43095
rect 17592 43052 17644 43061
rect 17684 43052 17736 43104
rect 18144 43095 18196 43104
rect 18144 43061 18153 43095
rect 18153 43061 18187 43095
rect 18187 43061 18196 43095
rect 18144 43052 18196 43061
rect 18420 43095 18472 43104
rect 18420 43061 18429 43095
rect 18429 43061 18463 43095
rect 18463 43061 18472 43095
rect 18420 43052 18472 43061
rect 18512 43052 18564 43104
rect 19524 43095 19576 43104
rect 19524 43061 19533 43095
rect 19533 43061 19567 43095
rect 19567 43061 19576 43095
rect 19524 43052 19576 43061
rect 24124 43095 24176 43104
rect 24124 43061 24133 43095
rect 24133 43061 24167 43095
rect 24167 43061 24176 43095
rect 24124 43052 24176 43061
rect 3917 42950 3969 43002
rect 3981 42950 4033 43002
rect 4045 42950 4097 43002
rect 4109 42950 4161 43002
rect 4173 42950 4225 43002
rect 9851 42950 9903 43002
rect 9915 42950 9967 43002
rect 9979 42950 10031 43002
rect 10043 42950 10095 43002
rect 10107 42950 10159 43002
rect 15785 42950 15837 43002
rect 15849 42950 15901 43002
rect 15913 42950 15965 43002
rect 15977 42950 16029 43002
rect 16041 42950 16093 43002
rect 21719 42950 21771 43002
rect 21783 42950 21835 43002
rect 21847 42950 21899 43002
rect 21911 42950 21963 43002
rect 21975 42950 22027 43002
rect 2228 42891 2280 42900
rect 2228 42857 2237 42891
rect 2237 42857 2271 42891
rect 2271 42857 2280 42891
rect 2228 42848 2280 42857
rect 3332 42891 3384 42900
rect 3332 42857 3341 42891
rect 3341 42857 3375 42891
rect 3375 42857 3384 42891
rect 3332 42848 3384 42857
rect 3792 42848 3844 42900
rect 6092 42891 6144 42900
rect 6092 42857 6101 42891
rect 6101 42857 6135 42891
rect 6135 42857 6144 42891
rect 6092 42848 6144 42857
rect 6828 42891 6880 42900
rect 6828 42857 6837 42891
rect 6837 42857 6871 42891
rect 6871 42857 6880 42891
rect 6828 42848 6880 42857
rect 7380 42891 7432 42900
rect 7380 42857 7389 42891
rect 7389 42857 7423 42891
rect 7423 42857 7432 42891
rect 7380 42848 7432 42857
rect 9496 42848 9548 42900
rect 9680 42848 9732 42900
rect 10600 42891 10652 42900
rect 10600 42857 10609 42891
rect 10609 42857 10643 42891
rect 10643 42857 10652 42891
rect 10600 42848 10652 42857
rect 1400 42712 1452 42764
rect 8392 42780 8444 42832
rect 16856 42848 16908 42900
rect 17684 42848 17736 42900
rect 2780 42712 2832 42764
rect 4896 42712 4948 42764
rect 8760 42712 8812 42764
rect 4252 42644 4304 42696
rect 4712 42644 4764 42696
rect 2596 42576 2648 42628
rect 3240 42619 3292 42628
rect 3240 42585 3249 42619
rect 3249 42585 3283 42619
rect 3283 42585 3292 42619
rect 3240 42576 3292 42585
rect 3884 42576 3936 42628
rect 3056 42508 3108 42560
rect 3148 42508 3200 42560
rect 4160 42508 4212 42560
rect 4620 42508 4672 42560
rect 4804 42508 4856 42560
rect 7748 42687 7800 42696
rect 7748 42653 7757 42687
rect 7757 42653 7791 42687
rect 7791 42653 7800 42687
rect 7748 42644 7800 42653
rect 9128 42687 9180 42696
rect 9128 42653 9137 42687
rect 9137 42653 9171 42687
rect 9171 42653 9180 42687
rect 9128 42644 9180 42653
rect 11152 42780 11204 42832
rect 9312 42712 9364 42764
rect 12256 42712 12308 42764
rect 9588 42644 9640 42696
rect 6000 42619 6052 42628
rect 6000 42585 6009 42619
rect 6009 42585 6043 42619
rect 6043 42585 6052 42619
rect 6000 42576 6052 42585
rect 6736 42619 6788 42628
rect 6736 42585 6745 42619
rect 6745 42585 6779 42619
rect 6779 42585 6788 42619
rect 6736 42576 6788 42585
rect 7288 42619 7340 42628
rect 7288 42585 7297 42619
rect 7297 42585 7331 42619
rect 7331 42585 7340 42619
rect 7288 42576 7340 42585
rect 5724 42551 5776 42560
rect 5724 42517 5733 42551
rect 5733 42517 5767 42551
rect 5767 42517 5776 42551
rect 5724 42508 5776 42517
rect 5908 42508 5960 42560
rect 7472 42508 7524 42560
rect 8760 42576 8812 42628
rect 10784 42687 10836 42696
rect 10784 42653 10793 42687
rect 10793 42653 10827 42687
rect 10827 42653 10836 42687
rect 10784 42644 10836 42653
rect 11612 42687 11664 42696
rect 11612 42653 11621 42687
rect 11621 42653 11655 42687
rect 11655 42653 11664 42687
rect 11612 42644 11664 42653
rect 11888 42687 11940 42696
rect 11888 42653 11897 42687
rect 11897 42653 11931 42687
rect 11931 42653 11940 42687
rect 11888 42644 11940 42653
rect 12992 42687 13044 42696
rect 12992 42653 13001 42687
rect 13001 42653 13035 42687
rect 13035 42653 13044 42687
rect 12992 42644 13044 42653
rect 8668 42508 8720 42560
rect 9312 42508 9364 42560
rect 9772 42508 9824 42560
rect 10324 42508 10376 42560
rect 11796 42551 11848 42560
rect 11796 42517 11805 42551
rect 11805 42517 11839 42551
rect 11839 42517 11848 42551
rect 11796 42508 11848 42517
rect 12072 42551 12124 42560
rect 12072 42517 12081 42551
rect 12081 42517 12115 42551
rect 12115 42517 12124 42551
rect 12072 42508 12124 42517
rect 13084 42576 13136 42628
rect 13820 42712 13872 42764
rect 14096 42687 14148 42696
rect 14096 42653 14105 42687
rect 14105 42653 14139 42687
rect 14139 42653 14148 42687
rect 14096 42644 14148 42653
rect 14372 42687 14424 42696
rect 14372 42653 14381 42687
rect 14381 42653 14415 42687
rect 14415 42653 14424 42687
rect 14372 42644 14424 42653
rect 15200 42712 15252 42764
rect 14924 42576 14976 42628
rect 16488 42687 16540 42696
rect 16488 42653 16497 42687
rect 16497 42653 16531 42687
rect 16531 42653 16540 42687
rect 16488 42644 16540 42653
rect 16580 42687 16632 42696
rect 16580 42653 16589 42687
rect 16589 42653 16623 42687
rect 16623 42653 16632 42687
rect 16580 42644 16632 42653
rect 16120 42576 16172 42628
rect 17592 42644 17644 42696
rect 18144 42848 18196 42900
rect 18880 42891 18932 42900
rect 18880 42857 18889 42891
rect 18889 42857 18923 42891
rect 18923 42857 18932 42891
rect 18880 42848 18932 42857
rect 18972 42848 19024 42900
rect 20812 42848 20864 42900
rect 18052 42823 18104 42832
rect 18052 42789 18061 42823
rect 18061 42789 18095 42823
rect 18095 42789 18104 42823
rect 18052 42780 18104 42789
rect 18420 42712 18472 42764
rect 18328 42644 18380 42696
rect 18972 42644 19024 42696
rect 14556 42551 14608 42560
rect 14556 42517 14565 42551
rect 14565 42517 14599 42551
rect 14599 42517 14608 42551
rect 14556 42508 14608 42517
rect 14832 42551 14884 42560
rect 14832 42517 14841 42551
rect 14841 42517 14875 42551
rect 14875 42517 14884 42551
rect 14832 42508 14884 42517
rect 15476 42551 15528 42560
rect 15476 42517 15485 42551
rect 15485 42517 15519 42551
rect 15519 42517 15528 42551
rect 15476 42508 15528 42517
rect 15568 42508 15620 42560
rect 16396 42508 16448 42560
rect 16948 42551 17000 42560
rect 16948 42517 16957 42551
rect 16957 42517 16991 42551
rect 16991 42517 17000 42551
rect 16948 42508 17000 42517
rect 17224 42551 17276 42560
rect 17224 42517 17233 42551
rect 17233 42517 17267 42551
rect 17267 42517 17276 42551
rect 17224 42508 17276 42517
rect 17316 42508 17368 42560
rect 17776 42551 17828 42560
rect 17776 42517 17785 42551
rect 17785 42517 17819 42551
rect 17819 42517 17828 42551
rect 17776 42508 17828 42517
rect 18236 42508 18288 42560
rect 18328 42551 18380 42560
rect 18328 42517 18337 42551
rect 18337 42517 18371 42551
rect 18371 42517 18380 42551
rect 18328 42508 18380 42517
rect 18604 42551 18656 42560
rect 18604 42517 18613 42551
rect 18613 42517 18647 42551
rect 18647 42517 18656 42551
rect 18604 42508 18656 42517
rect 21364 42712 21416 42764
rect 19248 42687 19300 42696
rect 19248 42653 19257 42687
rect 19257 42653 19291 42687
rect 19291 42653 19300 42687
rect 19248 42644 19300 42653
rect 21272 42687 21324 42696
rect 21272 42653 21281 42687
rect 21281 42653 21315 42687
rect 21315 42653 21324 42687
rect 21272 42644 21324 42653
rect 21916 42687 21968 42696
rect 21916 42653 21925 42687
rect 21925 42653 21959 42687
rect 21959 42653 21968 42687
rect 21916 42644 21968 42653
rect 22376 42644 22428 42696
rect 25136 42712 25188 42764
rect 24216 42644 24268 42696
rect 24584 42644 24636 42696
rect 20536 42551 20588 42560
rect 20536 42517 20545 42551
rect 20545 42517 20579 42551
rect 20579 42517 20588 42551
rect 20536 42508 20588 42517
rect 21548 42619 21600 42628
rect 21548 42585 21557 42619
rect 21557 42585 21591 42619
rect 21591 42585 21600 42619
rect 21548 42576 21600 42585
rect 21180 42508 21232 42560
rect 22284 42508 22336 42560
rect 23756 42619 23808 42628
rect 23756 42585 23765 42619
rect 23765 42585 23799 42619
rect 23799 42585 23808 42619
rect 23756 42576 23808 42585
rect 6884 42406 6936 42458
rect 6948 42406 7000 42458
rect 7012 42406 7064 42458
rect 7076 42406 7128 42458
rect 7140 42406 7192 42458
rect 12818 42406 12870 42458
rect 12882 42406 12934 42458
rect 12946 42406 12998 42458
rect 13010 42406 13062 42458
rect 13074 42406 13126 42458
rect 18752 42406 18804 42458
rect 18816 42406 18868 42458
rect 18880 42406 18932 42458
rect 18944 42406 18996 42458
rect 19008 42406 19060 42458
rect 24686 42406 24738 42458
rect 24750 42406 24802 42458
rect 24814 42406 24866 42458
rect 24878 42406 24930 42458
rect 24942 42406 24994 42458
rect 480 42304 532 42356
rect 2320 42304 2372 42356
rect 3148 42304 3200 42356
rect 3240 42304 3292 42356
rect 2044 42279 2096 42288
rect 2044 42245 2053 42279
rect 2053 42245 2087 42279
rect 2087 42245 2096 42279
rect 2044 42236 2096 42245
rect 4896 42304 4948 42356
rect 2136 42168 2188 42220
rect 2780 42211 2832 42220
rect 2780 42177 2789 42211
rect 2789 42177 2823 42211
rect 2823 42177 2832 42211
rect 2780 42168 2832 42177
rect 3332 42168 3384 42220
rect 3700 42168 3752 42220
rect 3976 42211 4028 42220
rect 3976 42177 3985 42211
rect 3985 42177 4019 42211
rect 4019 42177 4028 42211
rect 3976 42168 4028 42177
rect 4068 42168 4120 42220
rect 3516 42100 3568 42152
rect 4712 42211 4764 42220
rect 4712 42177 4721 42211
rect 4721 42177 4755 42211
rect 4755 42177 4764 42211
rect 4712 42168 4764 42177
rect 5172 42168 5224 42220
rect 5908 42304 5960 42356
rect 6276 42304 6328 42356
rect 7196 42304 7248 42356
rect 7380 42304 7432 42356
rect 8208 42304 8260 42356
rect 5448 42236 5500 42288
rect 5816 42236 5868 42288
rect 4988 42100 5040 42152
rect 6276 42100 6328 42152
rect 6920 42100 6972 42152
rect 7472 42211 7524 42220
rect 7472 42177 7481 42211
rect 7481 42177 7515 42211
rect 7515 42177 7524 42211
rect 7472 42168 7524 42177
rect 7656 42168 7708 42220
rect 8208 42211 8260 42220
rect 8208 42177 8217 42211
rect 8217 42177 8251 42211
rect 8251 42177 8260 42211
rect 8208 42168 8260 42177
rect 8576 42236 8628 42288
rect 9128 42236 9180 42288
rect 5816 42032 5868 42084
rect 7564 42032 7616 42084
rect 7840 42100 7892 42152
rect 8852 42168 8904 42220
rect 9036 42211 9088 42220
rect 9036 42177 9045 42211
rect 9045 42177 9079 42211
rect 9079 42177 9088 42211
rect 9036 42168 9088 42177
rect 9496 42168 9548 42220
rect 9772 42236 9824 42288
rect 14740 42236 14792 42288
rect 16396 42236 16448 42288
rect 17224 42304 17276 42356
rect 17316 42304 17368 42356
rect 17776 42304 17828 42356
rect 18328 42304 18380 42356
rect 16948 42236 17000 42288
rect 18052 42236 18104 42288
rect 18420 42236 18472 42288
rect 18604 42279 18656 42288
rect 18604 42245 18613 42279
rect 18613 42245 18647 42279
rect 18647 42245 18656 42279
rect 18604 42236 18656 42245
rect 19524 42236 19576 42288
rect 8760 42100 8812 42152
rect 17040 42168 17092 42220
rect 20628 42304 20680 42356
rect 20812 42347 20864 42356
rect 20812 42313 20821 42347
rect 20821 42313 20855 42347
rect 20855 42313 20864 42347
rect 20812 42304 20864 42313
rect 21640 42304 21692 42356
rect 1308 41964 1360 42016
rect 3332 41964 3384 42016
rect 4436 41964 4488 42016
rect 4528 42007 4580 42016
rect 4528 41973 4537 42007
rect 4537 41973 4571 42007
rect 4571 41973 4580 42007
rect 4528 41964 4580 41973
rect 4896 41964 4948 42016
rect 7104 41964 7156 42016
rect 7380 41964 7432 42016
rect 7932 41964 7984 42016
rect 8024 42007 8076 42016
rect 8024 41973 8033 42007
rect 8033 41973 8067 42007
rect 8067 41973 8076 42007
rect 8024 41964 8076 41973
rect 8852 42007 8904 42016
rect 8852 41973 8861 42007
rect 8861 41973 8895 42007
rect 8895 41973 8904 42007
rect 8852 41964 8904 41973
rect 11704 42100 11756 42152
rect 15384 42032 15436 42084
rect 16488 42032 16540 42084
rect 16948 42075 17000 42084
rect 16948 42041 16957 42075
rect 16957 42041 16991 42075
rect 16991 42041 17000 42075
rect 16948 42032 17000 42041
rect 17316 42075 17368 42084
rect 17316 42041 17325 42075
rect 17325 42041 17359 42075
rect 17359 42041 17368 42075
rect 17316 42032 17368 42041
rect 17684 42075 17736 42084
rect 17684 42041 17693 42075
rect 17693 42041 17727 42075
rect 17727 42041 17736 42075
rect 17684 42032 17736 42041
rect 18052 42075 18104 42084
rect 18052 42041 18061 42075
rect 18061 42041 18095 42075
rect 18095 42041 18104 42075
rect 18052 42032 18104 42041
rect 9772 41964 9824 42016
rect 16304 42007 16356 42016
rect 16304 41973 16313 42007
rect 16313 41973 16347 42007
rect 16347 41973 16356 42007
rect 16304 41964 16356 41973
rect 18328 42007 18380 42016
rect 18328 41973 18337 42007
rect 18337 41973 18371 42007
rect 18371 41973 18380 42007
rect 18328 41964 18380 41973
rect 18512 41964 18564 42016
rect 19524 42075 19576 42084
rect 19524 42041 19533 42075
rect 19533 42041 19567 42075
rect 19567 42041 19576 42075
rect 19524 42032 19576 42041
rect 19892 42032 19944 42084
rect 20260 42100 20312 42152
rect 20996 42211 21048 42220
rect 20996 42177 21005 42211
rect 21005 42177 21039 42211
rect 21039 42177 21048 42211
rect 20996 42168 21048 42177
rect 21272 42211 21324 42220
rect 21272 42177 21281 42211
rect 21281 42177 21315 42211
rect 21315 42177 21324 42211
rect 21272 42168 21324 42177
rect 22744 42236 22796 42288
rect 23204 42304 23256 42356
rect 24492 42304 24544 42356
rect 25596 42304 25648 42356
rect 20904 42100 20956 42152
rect 20996 42032 21048 42084
rect 22836 42211 22888 42220
rect 22836 42177 22845 42211
rect 22845 42177 22879 42211
rect 22879 42177 22888 42211
rect 22836 42168 22888 42177
rect 22376 42100 22428 42152
rect 24032 42211 24084 42220
rect 24032 42177 24041 42211
rect 24041 42177 24075 42211
rect 24075 42177 24084 42211
rect 24032 42168 24084 42177
rect 23572 42032 23624 42084
rect 24584 42100 24636 42152
rect 24216 42032 24268 42084
rect 19708 41964 19760 42016
rect 22284 41964 22336 42016
rect 23480 41964 23532 42016
rect 25136 41964 25188 42016
rect 3917 41862 3969 41914
rect 3981 41862 4033 41914
rect 4045 41862 4097 41914
rect 4109 41862 4161 41914
rect 4173 41862 4225 41914
rect 9851 41862 9903 41914
rect 9915 41862 9967 41914
rect 9979 41862 10031 41914
rect 10043 41862 10095 41914
rect 10107 41862 10159 41914
rect 15785 41862 15837 41914
rect 15849 41862 15901 41914
rect 15913 41862 15965 41914
rect 15977 41862 16029 41914
rect 16041 41862 16093 41914
rect 21719 41862 21771 41914
rect 21783 41862 21835 41914
rect 21847 41862 21899 41914
rect 21911 41862 21963 41914
rect 21975 41862 22027 41914
rect 940 41760 992 41812
rect 1676 41760 1728 41812
rect 2504 41803 2556 41812
rect 2504 41769 2513 41803
rect 2513 41769 2547 41803
rect 2547 41769 2556 41803
rect 2504 41760 2556 41769
rect 2596 41760 2648 41812
rect 2780 41760 2832 41812
rect 3424 41803 3476 41812
rect 3424 41769 3433 41803
rect 3433 41769 3467 41803
rect 3467 41769 3476 41803
rect 3424 41760 3476 41769
rect 3884 41760 3936 41812
rect 4252 41760 4304 41812
rect 4988 41760 5040 41812
rect 1124 41624 1176 41676
rect 2872 41624 2924 41676
rect 4804 41692 4856 41744
rect 5540 41760 5592 41812
rect 6000 41760 6052 41812
rect 6736 41760 6788 41812
rect 7288 41760 7340 41812
rect 7380 41760 7432 41812
rect 7748 41760 7800 41812
rect 7932 41760 7984 41812
rect 8116 41803 8168 41812
rect 8116 41769 8125 41803
rect 8125 41769 8159 41803
rect 8159 41769 8168 41803
rect 8116 41760 8168 41769
rect 8392 41803 8444 41812
rect 8392 41769 8401 41803
rect 8401 41769 8435 41803
rect 8435 41769 8444 41803
rect 8392 41760 8444 41769
rect 8852 41760 8904 41812
rect 8944 41803 8996 41812
rect 8944 41769 8953 41803
rect 8953 41769 8987 41803
rect 8987 41769 8996 41803
rect 8944 41760 8996 41769
rect 9036 41760 9088 41812
rect 12532 41760 12584 41812
rect 17868 41760 17920 41812
rect 1768 41488 1820 41540
rect 3148 41556 3200 41608
rect 3424 41556 3476 41608
rect 4252 41599 4304 41608
rect 4252 41565 4261 41599
rect 4261 41565 4295 41599
rect 4295 41565 4304 41599
rect 4252 41556 4304 41565
rect 4528 41599 4580 41608
rect 4528 41565 4537 41599
rect 4537 41565 4571 41599
rect 4571 41565 4580 41599
rect 4528 41556 4580 41565
rect 4804 41599 4856 41608
rect 4804 41565 4813 41599
rect 4813 41565 4847 41599
rect 4847 41565 4856 41599
rect 4804 41556 4856 41565
rect 572 41420 624 41472
rect 2688 41420 2740 41472
rect 2872 41420 2924 41472
rect 3148 41420 3200 41472
rect 4896 41488 4948 41540
rect 5172 41624 5224 41676
rect 5356 41599 5408 41608
rect 5356 41565 5365 41599
rect 5365 41565 5399 41599
rect 5399 41565 5408 41599
rect 5356 41556 5408 41565
rect 5816 41556 5868 41608
rect 7564 41624 7616 41676
rect 6092 41420 6144 41472
rect 8576 41599 8628 41608
rect 8576 41565 8585 41599
rect 8585 41565 8619 41599
rect 8619 41565 8628 41599
rect 8576 41556 8628 41565
rect 10508 41624 10560 41676
rect 17960 41735 18012 41744
rect 17960 41701 17969 41735
rect 17969 41701 18003 41735
rect 18003 41701 18012 41735
rect 17960 41692 18012 41701
rect 18236 41760 18288 41812
rect 19156 41760 19208 41812
rect 19432 41760 19484 41812
rect 19708 41760 19760 41812
rect 9680 41599 9732 41608
rect 9680 41565 9689 41599
rect 9689 41565 9723 41599
rect 9723 41565 9732 41599
rect 9680 41556 9732 41565
rect 9864 41556 9916 41608
rect 18236 41556 18288 41608
rect 18420 41556 18472 41608
rect 18972 41599 19024 41608
rect 18972 41565 18981 41599
rect 18981 41565 19015 41599
rect 19015 41565 19024 41599
rect 18972 41556 19024 41565
rect 20444 41692 20496 41744
rect 20536 41692 20588 41744
rect 20720 41803 20772 41812
rect 20720 41769 20729 41803
rect 20729 41769 20763 41803
rect 20763 41769 20772 41803
rect 20720 41760 20772 41769
rect 20812 41760 20864 41812
rect 21088 41760 21140 41812
rect 22928 41760 22980 41812
rect 23664 41760 23716 41812
rect 25320 41760 25372 41812
rect 21640 41692 21692 41744
rect 21824 41692 21876 41744
rect 10600 41488 10652 41540
rect 17960 41488 18012 41540
rect 19432 41488 19484 41540
rect 7196 41420 7248 41472
rect 9956 41420 10008 41472
rect 18144 41420 18196 41472
rect 18420 41463 18472 41472
rect 18420 41429 18429 41463
rect 18429 41429 18463 41463
rect 18463 41429 18472 41463
rect 18420 41420 18472 41429
rect 19340 41420 19392 41472
rect 21640 41599 21692 41608
rect 21640 41565 21649 41599
rect 21649 41565 21683 41599
rect 21683 41565 21692 41599
rect 21640 41556 21692 41565
rect 22284 41624 22336 41676
rect 20260 41463 20312 41472
rect 20260 41429 20269 41463
rect 20269 41429 20303 41463
rect 20303 41429 20312 41463
rect 20260 41420 20312 41429
rect 22376 41488 22428 41540
rect 22652 41488 22704 41540
rect 22928 41488 22980 41540
rect 25228 41692 25280 41744
rect 23848 41531 23900 41540
rect 23848 41497 23857 41531
rect 23857 41497 23891 41531
rect 23891 41497 23900 41531
rect 23848 41488 23900 41497
rect 21456 41463 21508 41472
rect 21456 41429 21465 41463
rect 21465 41429 21499 41463
rect 21499 41429 21508 41463
rect 21456 41420 21508 41429
rect 22008 41420 22060 41472
rect 22560 41420 22612 41472
rect 25504 41420 25556 41472
rect 6884 41318 6936 41370
rect 6948 41318 7000 41370
rect 7012 41318 7064 41370
rect 7076 41318 7128 41370
rect 7140 41318 7192 41370
rect 12818 41318 12870 41370
rect 12882 41318 12934 41370
rect 12946 41318 12998 41370
rect 13010 41318 13062 41370
rect 13074 41318 13126 41370
rect 18752 41318 18804 41370
rect 18816 41318 18868 41370
rect 18880 41318 18932 41370
rect 18944 41318 18996 41370
rect 19008 41318 19060 41370
rect 24686 41318 24738 41370
rect 24750 41318 24802 41370
rect 24814 41318 24866 41370
rect 24878 41318 24930 41370
rect 24942 41318 24994 41370
rect 2412 41216 2464 41268
rect 2780 41216 2832 41268
rect 7564 41216 7616 41268
rect 7840 41216 7892 41268
rect 8024 41216 8076 41268
rect 14648 41216 14700 41268
rect 15108 41216 15160 41268
rect 1216 41080 1268 41132
rect 2228 41123 2280 41132
rect 2228 41089 2237 41123
rect 2237 41089 2271 41123
rect 2271 41089 2280 41123
rect 2228 41080 2280 41089
rect 3240 41123 3292 41132
rect 3240 41089 3249 41123
rect 3249 41089 3283 41123
rect 3283 41089 3292 41123
rect 3240 41080 3292 41089
rect 3792 41123 3844 41132
rect 3792 41089 3799 41123
rect 3799 41089 3833 41123
rect 3833 41089 3844 41123
rect 3792 41080 3844 41089
rect 5540 41148 5592 41200
rect 3516 41055 3568 41064
rect 3516 41021 3525 41055
rect 3525 41021 3559 41055
rect 3559 41021 3568 41055
rect 3516 41012 3568 41021
rect 2872 40876 2924 40928
rect 4528 40919 4580 40928
rect 4528 40885 4537 40919
rect 4537 40885 4571 40919
rect 4571 40885 4580 40919
rect 4528 40876 4580 40885
rect 6000 40876 6052 40928
rect 6920 40987 6972 40996
rect 6920 40953 6929 40987
rect 6929 40953 6963 40987
rect 6963 40953 6972 40987
rect 6920 40944 6972 40953
rect 7932 41123 7984 41132
rect 7932 41089 7941 41123
rect 7941 41089 7975 41123
rect 7975 41089 7984 41123
rect 7932 41080 7984 41089
rect 12440 41148 12492 41200
rect 9680 41080 9732 41132
rect 10416 41080 10468 41132
rect 19800 41259 19852 41268
rect 19800 41225 19809 41259
rect 19809 41225 19843 41259
rect 19843 41225 19852 41259
rect 19800 41216 19852 41225
rect 20352 41259 20404 41268
rect 20352 41225 20361 41259
rect 20361 41225 20395 41259
rect 20395 41225 20404 41259
rect 20352 41216 20404 41225
rect 20628 41259 20680 41268
rect 20628 41225 20637 41259
rect 20637 41225 20671 41259
rect 20671 41225 20680 41259
rect 20628 41216 20680 41225
rect 21180 41216 21232 41268
rect 21272 41216 21324 41268
rect 19708 41123 19760 41132
rect 19708 41089 19717 41123
rect 19717 41089 19751 41123
rect 19751 41089 19760 41123
rect 19708 41080 19760 41089
rect 19892 41080 19944 41132
rect 8576 41055 8628 41064
rect 8576 41021 8585 41055
rect 8585 41021 8619 41055
rect 8619 41021 8628 41055
rect 8576 41012 8628 41021
rect 9496 41012 9548 41064
rect 7380 40876 7432 40928
rect 7472 40919 7524 40928
rect 7472 40885 7481 40919
rect 7481 40885 7515 40919
rect 7515 40885 7524 40919
rect 7472 40876 7524 40885
rect 7748 40876 7800 40928
rect 7840 40876 7892 40928
rect 9864 40944 9916 40996
rect 9588 40919 9640 40928
rect 9588 40885 9597 40919
rect 9597 40885 9631 40919
rect 9631 40885 9640 40919
rect 9588 40876 9640 40885
rect 11704 41012 11756 41064
rect 16396 41012 16448 41064
rect 20536 41123 20588 41132
rect 20536 41089 20545 41123
rect 20545 41089 20579 41123
rect 20579 41089 20588 41123
rect 20536 41080 20588 41089
rect 20628 41080 20680 41132
rect 21180 41080 21232 41132
rect 21272 41080 21324 41132
rect 20444 41012 20496 41064
rect 20720 41012 20772 41064
rect 22008 41216 22060 41268
rect 22468 41216 22520 41268
rect 23388 41216 23440 41268
rect 25044 41216 25096 41268
rect 21824 41080 21876 41132
rect 22192 41080 22244 41132
rect 22468 41080 22520 41132
rect 22744 41012 22796 41064
rect 11060 40919 11112 40928
rect 11060 40885 11069 40919
rect 11069 40885 11103 40919
rect 11103 40885 11112 40919
rect 11060 40876 11112 40885
rect 19064 40919 19116 40928
rect 19064 40885 19073 40919
rect 19073 40885 19107 40919
rect 19107 40885 19116 40919
rect 19064 40876 19116 40885
rect 20444 40876 20496 40928
rect 21456 40876 21508 40928
rect 21640 40944 21692 40996
rect 23480 41148 23532 41200
rect 23112 41080 23164 41132
rect 23296 41012 23348 41064
rect 21732 40876 21784 40928
rect 22100 40876 22152 40928
rect 23664 40919 23716 40928
rect 23664 40885 23673 40919
rect 23673 40885 23707 40919
rect 23707 40885 23716 40919
rect 23664 40876 23716 40885
rect 3917 40774 3969 40826
rect 3981 40774 4033 40826
rect 4045 40774 4097 40826
rect 4109 40774 4161 40826
rect 4173 40774 4225 40826
rect 9851 40774 9903 40826
rect 9915 40774 9967 40826
rect 9979 40774 10031 40826
rect 10043 40774 10095 40826
rect 10107 40774 10159 40826
rect 15785 40774 15837 40826
rect 15849 40774 15901 40826
rect 15913 40774 15965 40826
rect 15977 40774 16029 40826
rect 16041 40774 16093 40826
rect 21719 40774 21771 40826
rect 21783 40774 21835 40826
rect 21847 40774 21899 40826
rect 21911 40774 21963 40826
rect 21975 40774 22027 40826
rect 2780 40672 2832 40724
rect 3056 40672 3108 40724
rect 3792 40672 3844 40724
rect 4804 40647 4856 40656
rect 4804 40613 4813 40647
rect 4813 40613 4847 40647
rect 4847 40613 4856 40647
rect 4804 40604 4856 40613
rect 3516 40536 3568 40588
rect 1860 40468 1912 40520
rect 1400 40443 1452 40452
rect 1400 40409 1409 40443
rect 1409 40409 1443 40443
rect 1443 40409 1452 40443
rect 1400 40400 1452 40409
rect 2780 40400 2832 40452
rect 3056 40400 3108 40452
rect 5540 40579 5592 40588
rect 5540 40545 5549 40579
rect 5549 40545 5583 40579
rect 5583 40545 5592 40579
rect 5540 40536 5592 40545
rect 3976 40468 4028 40520
rect 5448 40468 5500 40520
rect 8024 40672 8076 40724
rect 6736 40400 6788 40452
rect 7840 40468 7892 40520
rect 7656 40400 7708 40452
rect 10324 40604 10376 40656
rect 10508 40647 10560 40656
rect 10508 40613 10517 40647
rect 10517 40613 10551 40647
rect 10551 40613 10560 40647
rect 10508 40604 10560 40613
rect 10968 40672 11020 40724
rect 3700 40332 3752 40384
rect 5080 40332 5132 40384
rect 6644 40332 6696 40384
rect 7932 40375 7984 40384
rect 7932 40341 7941 40375
rect 7941 40341 7975 40375
rect 7975 40341 7984 40375
rect 7932 40332 7984 40341
rect 8024 40332 8076 40384
rect 8392 40332 8444 40384
rect 8944 40332 8996 40384
rect 9128 40332 9180 40384
rect 10784 40511 10836 40520
rect 10784 40477 10793 40511
rect 10793 40477 10827 40511
rect 10827 40477 10836 40511
rect 10784 40468 10836 40477
rect 11060 40579 11112 40588
rect 11060 40545 11069 40579
rect 11069 40545 11103 40579
rect 11103 40545 11112 40579
rect 11060 40536 11112 40545
rect 11612 40536 11664 40588
rect 16396 40672 16448 40724
rect 19064 40672 19116 40724
rect 12716 40468 12768 40520
rect 19708 40604 19760 40656
rect 20260 40647 20312 40656
rect 20260 40613 20269 40647
rect 20269 40613 20303 40647
rect 20303 40613 20312 40647
rect 20260 40604 20312 40613
rect 20444 40604 20496 40656
rect 21088 40715 21140 40724
rect 21088 40681 21097 40715
rect 21097 40681 21131 40715
rect 21131 40681 21140 40715
rect 21088 40672 21140 40681
rect 21272 40672 21324 40724
rect 21732 40672 21784 40724
rect 22192 40715 22244 40724
rect 22192 40681 22201 40715
rect 22201 40681 22235 40715
rect 22235 40681 22244 40715
rect 22192 40672 22244 40681
rect 22468 40715 22520 40724
rect 22468 40681 22477 40715
rect 22477 40681 22511 40715
rect 22511 40681 22520 40715
rect 22468 40672 22520 40681
rect 22744 40715 22796 40724
rect 22744 40681 22753 40715
rect 22753 40681 22787 40715
rect 22787 40681 22796 40715
rect 22744 40672 22796 40681
rect 23020 40715 23072 40724
rect 23020 40681 23029 40715
rect 23029 40681 23063 40715
rect 23063 40681 23072 40715
rect 23020 40672 23072 40681
rect 24032 40672 24084 40724
rect 19248 40536 19300 40588
rect 22008 40604 22060 40656
rect 19432 40468 19484 40520
rect 12440 40400 12492 40452
rect 17408 40400 17460 40452
rect 20168 40511 20220 40520
rect 20168 40477 20177 40511
rect 20177 40477 20211 40511
rect 20211 40477 20220 40511
rect 20168 40468 20220 40477
rect 21088 40468 21140 40520
rect 21640 40536 21692 40588
rect 21456 40468 21508 40520
rect 22100 40511 22152 40520
rect 22100 40477 22109 40511
rect 22109 40477 22143 40511
rect 22143 40477 22152 40511
rect 22100 40468 22152 40477
rect 11152 40332 11204 40384
rect 12164 40332 12216 40384
rect 12348 40332 12400 40384
rect 19616 40375 19668 40384
rect 19616 40341 19625 40375
rect 19625 40341 19659 40375
rect 19659 40341 19668 40375
rect 19616 40332 19668 40341
rect 20076 40332 20128 40384
rect 21272 40332 21324 40384
rect 22284 40536 22336 40588
rect 23480 40536 23532 40588
rect 22560 40468 22612 40520
rect 22652 40511 22704 40520
rect 22652 40477 22661 40511
rect 22661 40477 22695 40511
rect 22695 40477 22704 40511
rect 22652 40468 22704 40477
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 23296 40468 23348 40520
rect 23664 40511 23716 40520
rect 23664 40477 23673 40511
rect 23673 40477 23707 40511
rect 23707 40477 23716 40511
rect 23664 40468 23716 40477
rect 23020 40400 23072 40452
rect 25136 40400 25188 40452
rect 22928 40332 22980 40384
rect 23480 40332 23532 40384
rect 25780 40332 25832 40384
rect 6884 40230 6936 40282
rect 6948 40230 7000 40282
rect 7012 40230 7064 40282
rect 7076 40230 7128 40282
rect 7140 40230 7192 40282
rect 12818 40230 12870 40282
rect 12882 40230 12934 40282
rect 12946 40230 12998 40282
rect 13010 40230 13062 40282
rect 13074 40230 13126 40282
rect 18752 40230 18804 40282
rect 18816 40230 18868 40282
rect 18880 40230 18932 40282
rect 18944 40230 18996 40282
rect 19008 40230 19060 40282
rect 24686 40230 24738 40282
rect 24750 40230 24802 40282
rect 24814 40230 24866 40282
rect 24878 40230 24930 40282
rect 24942 40230 24994 40282
rect 2872 40128 2924 40180
rect 2964 40128 3016 40180
rect 2228 40065 2280 40112
rect 1492 39992 1544 40044
rect 2228 40060 2253 40065
rect 2253 40060 2280 40065
rect 5172 40128 5224 40180
rect 5448 40128 5500 40180
rect 2320 39992 2372 40044
rect 3148 39992 3200 40044
rect 1768 39924 1820 39976
rect 3240 39924 3292 39976
rect 4344 40035 4396 40044
rect 4344 40001 4353 40035
rect 4353 40001 4387 40035
rect 4387 40001 4396 40035
rect 4344 39992 4396 40001
rect 5540 40060 5592 40112
rect 7288 40128 7340 40180
rect 7656 40128 7708 40180
rect 8024 40060 8076 40112
rect 8208 40103 8260 40112
rect 8208 40069 8217 40103
rect 8217 40069 8251 40103
rect 8251 40069 8260 40103
rect 8208 40060 8260 40069
rect 6460 39992 6512 40044
rect 9128 40103 9180 40112
rect 9128 40069 9137 40103
rect 9137 40069 9171 40103
rect 9171 40069 9180 40103
rect 9128 40060 9180 40069
rect 9312 40060 9364 40112
rect 9772 40060 9824 40112
rect 19616 40128 19668 40180
rect 7932 39924 7984 39976
rect 2872 39856 2924 39908
rect 3976 39856 4028 39908
rect 9680 39992 9732 40044
rect 10324 40060 10376 40112
rect 21824 40171 21876 40180
rect 21824 40137 21833 40171
rect 21833 40137 21867 40171
rect 21867 40137 21876 40171
rect 21824 40128 21876 40137
rect 21916 40128 21968 40180
rect 22192 40128 22244 40180
rect 10784 39992 10836 40044
rect 12716 40035 12768 40044
rect 12716 40001 12725 40035
rect 12725 40001 12759 40035
rect 12759 40001 12768 40035
rect 12716 39992 12768 40001
rect 19984 40035 20036 40044
rect 19984 40001 19993 40035
rect 19993 40001 20027 40035
rect 20027 40001 20036 40035
rect 19984 39992 20036 40001
rect 22652 40060 22704 40112
rect 20720 39992 20772 40044
rect 20904 39992 20956 40044
rect 21272 39992 21324 40044
rect 21364 40035 21416 40044
rect 21364 40001 21373 40035
rect 21373 40001 21407 40035
rect 21407 40001 21416 40035
rect 21364 39992 21416 40001
rect 21640 40035 21692 40044
rect 21640 40001 21649 40035
rect 21649 40001 21683 40035
rect 21683 40001 21692 40035
rect 21640 39992 21692 40001
rect 22008 40035 22060 40044
rect 22008 40001 22017 40035
rect 22017 40001 22051 40035
rect 22051 40001 22060 40035
rect 22008 39992 22060 40001
rect 22192 39992 22244 40044
rect 9588 39924 9640 39976
rect 11244 39924 11296 39976
rect 2320 39788 2372 39840
rect 3516 39788 3568 39840
rect 4620 39831 4672 39840
rect 4620 39797 4629 39831
rect 4629 39797 4663 39831
rect 4663 39797 4672 39831
rect 4620 39788 4672 39797
rect 5908 39831 5960 39840
rect 5908 39797 5917 39831
rect 5917 39797 5951 39831
rect 5951 39797 5960 39831
rect 5908 39788 5960 39797
rect 10416 39831 10468 39840
rect 10416 39797 10425 39831
rect 10425 39797 10459 39831
rect 10459 39797 10468 39831
rect 10416 39788 10468 39797
rect 11796 39788 11848 39840
rect 12348 39924 12400 39976
rect 12164 39788 12216 39840
rect 13360 39924 13412 39976
rect 22744 39992 22796 40044
rect 23848 40128 23900 40180
rect 19432 39899 19484 39908
rect 19432 39865 19441 39899
rect 19441 39865 19475 39899
rect 19475 39865 19484 39899
rect 19432 39856 19484 39865
rect 19800 39899 19852 39908
rect 19800 39865 19809 39899
rect 19809 39865 19843 39899
rect 19843 39865 19852 39899
rect 19800 39856 19852 39865
rect 20076 39899 20128 39908
rect 20076 39865 20085 39899
rect 20085 39865 20119 39899
rect 20119 39865 20128 39899
rect 20076 39856 20128 39865
rect 21824 39856 21876 39908
rect 20904 39788 20956 39840
rect 21272 39788 21324 39840
rect 21732 39788 21784 39840
rect 22836 39856 22888 39908
rect 23756 39992 23808 40044
rect 24124 40035 24176 40044
rect 24124 40001 24133 40035
rect 24133 40001 24167 40035
rect 24167 40001 24176 40035
rect 24124 39992 24176 40001
rect 22284 39788 22336 39840
rect 22928 39831 22980 39840
rect 22928 39797 22937 39831
rect 22937 39797 22971 39831
rect 22971 39797 22980 39831
rect 22928 39788 22980 39797
rect 23940 39788 23992 39840
rect 24400 39831 24452 39840
rect 24400 39797 24409 39831
rect 24409 39797 24443 39831
rect 24443 39797 24452 39831
rect 24400 39788 24452 39797
rect 3917 39686 3969 39738
rect 3981 39686 4033 39738
rect 4045 39686 4097 39738
rect 4109 39686 4161 39738
rect 4173 39686 4225 39738
rect 9851 39686 9903 39738
rect 9915 39686 9967 39738
rect 9979 39686 10031 39738
rect 10043 39686 10095 39738
rect 10107 39686 10159 39738
rect 15785 39686 15837 39738
rect 15849 39686 15901 39738
rect 15913 39686 15965 39738
rect 15977 39686 16029 39738
rect 16041 39686 16093 39738
rect 21719 39686 21771 39738
rect 21783 39686 21835 39738
rect 21847 39686 21899 39738
rect 21911 39686 21963 39738
rect 21975 39686 22027 39738
rect 3148 39584 3200 39636
rect 3516 39584 3568 39636
rect 5908 39584 5960 39636
rect 6736 39584 6788 39636
rect 2688 39448 2740 39500
rect 4804 39448 4856 39500
rect 5264 39448 5316 39500
rect 7748 39584 7800 39636
rect 8392 39627 8444 39636
rect 8392 39593 8401 39627
rect 8401 39593 8435 39627
rect 8435 39593 8444 39627
rect 8392 39584 8444 39593
rect 9772 39584 9824 39636
rect 13360 39627 13412 39636
rect 13360 39593 13369 39627
rect 13369 39593 13403 39627
rect 13403 39593 13412 39627
rect 13360 39584 13412 39593
rect 19984 39584 20036 39636
rect 20996 39584 21048 39636
rect 21088 39584 21140 39636
rect 22284 39584 22336 39636
rect 22560 39584 22612 39636
rect 3516 39380 3568 39432
rect 4528 39380 4580 39432
rect 1492 39355 1544 39364
rect 1492 39321 1501 39355
rect 1501 39321 1535 39355
rect 1535 39321 1544 39355
rect 1492 39312 1544 39321
rect 1676 39355 1728 39364
rect 1676 39321 1685 39355
rect 1685 39321 1719 39355
rect 1719 39321 1728 39355
rect 1676 39312 1728 39321
rect 2320 39355 2372 39364
rect 2320 39321 2329 39355
rect 2329 39321 2363 39355
rect 2363 39321 2372 39355
rect 2320 39312 2372 39321
rect 2596 39312 2648 39364
rect 1952 39287 2004 39296
rect 1952 39253 1961 39287
rect 1961 39253 1995 39287
rect 1995 39253 2004 39287
rect 1952 39244 2004 39253
rect 2964 39244 3016 39296
rect 3976 39287 4028 39296
rect 3976 39253 3985 39287
rect 3985 39253 4019 39287
rect 4019 39253 4028 39287
rect 3976 39244 4028 39253
rect 4252 39355 4304 39364
rect 4252 39321 4261 39355
rect 4261 39321 4295 39355
rect 4295 39321 4304 39355
rect 4252 39312 4304 39321
rect 4712 39355 4764 39364
rect 4712 39321 4721 39355
rect 4721 39321 4755 39355
rect 4755 39321 4764 39355
rect 6460 39423 6512 39432
rect 6460 39389 6494 39423
rect 6494 39389 6512 39423
rect 6460 39380 6512 39389
rect 6644 39423 6696 39432
rect 6644 39389 6653 39423
rect 6653 39389 6687 39423
rect 6687 39389 6696 39423
rect 6644 39380 6696 39389
rect 11612 39448 11664 39500
rect 7564 39380 7616 39432
rect 8576 39380 8628 39432
rect 9404 39380 9456 39432
rect 9772 39423 9824 39432
rect 9772 39389 9779 39423
rect 9779 39389 9813 39423
rect 9813 39389 9824 39423
rect 9772 39380 9824 39389
rect 20904 39423 20956 39432
rect 20904 39389 20913 39423
rect 20913 39389 20947 39423
rect 20947 39389 20956 39423
rect 20904 39380 20956 39389
rect 21088 39380 21140 39432
rect 21272 39423 21324 39432
rect 21272 39389 21281 39423
rect 21281 39389 21315 39423
rect 21315 39389 21324 39423
rect 21272 39380 21324 39389
rect 4712 39312 4764 39321
rect 10416 39312 10468 39364
rect 11704 39312 11756 39364
rect 12256 39312 12308 39364
rect 4528 39244 4580 39296
rect 4988 39244 5040 39296
rect 5172 39244 5224 39296
rect 7288 39287 7340 39296
rect 7288 39253 7297 39287
rect 7297 39253 7331 39287
rect 7331 39253 7340 39287
rect 7288 39244 7340 39253
rect 7564 39244 7616 39296
rect 10508 39244 10560 39296
rect 21732 39423 21784 39432
rect 21732 39389 21741 39423
rect 21741 39389 21775 39423
rect 21775 39389 21784 39423
rect 21732 39380 21784 39389
rect 22008 39423 22060 39432
rect 22008 39389 22017 39423
rect 22017 39389 22051 39423
rect 22051 39389 22060 39423
rect 22008 39380 22060 39389
rect 22284 39423 22336 39432
rect 22284 39389 22293 39423
rect 22293 39389 22327 39423
rect 22327 39389 22336 39423
rect 22284 39380 22336 39389
rect 22560 39423 22612 39432
rect 22560 39389 22569 39423
rect 22569 39389 22603 39423
rect 22603 39389 22612 39423
rect 22560 39380 22612 39389
rect 23388 39423 23440 39432
rect 23388 39389 23397 39423
rect 23397 39389 23431 39423
rect 23431 39389 23440 39423
rect 23388 39380 23440 39389
rect 23848 39423 23900 39432
rect 23848 39389 23857 39423
rect 23857 39389 23891 39423
rect 23891 39389 23900 39423
rect 23848 39380 23900 39389
rect 23940 39423 23992 39432
rect 23940 39389 23949 39423
rect 23949 39389 23983 39423
rect 23983 39389 23992 39423
rect 23940 39380 23992 39389
rect 23112 39244 23164 39296
rect 23940 39244 23992 39296
rect 25228 39244 25280 39296
rect 6884 39142 6936 39194
rect 6948 39142 7000 39194
rect 7012 39142 7064 39194
rect 7076 39142 7128 39194
rect 7140 39142 7192 39194
rect 12818 39142 12870 39194
rect 12882 39142 12934 39194
rect 12946 39142 12998 39194
rect 13010 39142 13062 39194
rect 13074 39142 13126 39194
rect 18752 39142 18804 39194
rect 18816 39142 18868 39194
rect 18880 39142 18932 39194
rect 18944 39142 18996 39194
rect 19008 39142 19060 39194
rect 24686 39142 24738 39194
rect 24750 39142 24802 39194
rect 24814 39142 24866 39194
rect 24878 39142 24930 39194
rect 24942 39142 24994 39194
rect 1492 39040 1544 39092
rect 1952 39040 2004 39092
rect 3976 39040 4028 39092
rect 7288 39040 7340 39092
rect 7380 39040 7432 39092
rect 7656 39040 7708 39092
rect 8852 39040 8904 39092
rect 13452 39040 13504 39092
rect 7748 38972 7800 39024
rect 8484 38972 8536 39024
rect 11612 38972 11664 39024
rect 12532 38972 12584 39024
rect 19984 38972 20036 39024
rect 20904 39040 20956 39092
rect 21272 39040 21324 39092
rect 21364 39040 21416 39092
rect 22008 39040 22060 39092
rect 21456 38972 21508 39024
rect 23848 39040 23900 39092
rect 2872 38904 2924 38956
rect 3056 38947 3108 38956
rect 3056 38913 3065 38947
rect 3065 38913 3099 38947
rect 3099 38913 3108 38947
rect 3056 38904 3108 38913
rect 3424 38904 3476 38956
rect 2688 38836 2740 38888
rect 3792 38879 3844 38888
rect 3792 38845 3801 38879
rect 3801 38845 3835 38879
rect 3835 38845 3844 38879
rect 3792 38836 3844 38845
rect 3884 38836 3936 38888
rect 6736 38904 6788 38956
rect 7380 38904 7432 38956
rect 20628 38947 20680 38956
rect 20628 38913 20637 38947
rect 20637 38913 20671 38947
rect 20671 38913 20680 38947
rect 20628 38904 20680 38913
rect 7932 38836 7984 38888
rect 1768 38700 1820 38752
rect 2964 38768 3016 38820
rect 4988 38768 5040 38820
rect 7748 38768 7800 38820
rect 11520 38879 11572 38888
rect 11520 38845 11529 38879
rect 11529 38845 11563 38879
rect 11563 38845 11572 38879
rect 11520 38836 11572 38845
rect 16672 38768 16724 38820
rect 20996 38904 21048 38956
rect 21548 38836 21600 38888
rect 23572 38947 23624 38956
rect 23572 38913 23581 38947
rect 23581 38913 23615 38947
rect 23615 38913 23624 38947
rect 23572 38904 23624 38913
rect 23664 38904 23716 38956
rect 4344 38700 4396 38752
rect 8576 38700 8628 38752
rect 9128 38743 9180 38752
rect 9128 38709 9137 38743
rect 9137 38709 9171 38743
rect 9171 38709 9180 38743
rect 9128 38700 9180 38709
rect 12532 38743 12584 38752
rect 12532 38709 12541 38743
rect 12541 38709 12575 38743
rect 12575 38709 12584 38743
rect 12532 38700 12584 38709
rect 14464 38700 14516 38752
rect 18604 38700 18656 38752
rect 22100 38700 22152 38752
rect 22192 38700 22244 38752
rect 23848 38768 23900 38820
rect 23296 38700 23348 38752
rect 24032 38700 24084 38752
rect 24400 38743 24452 38752
rect 24400 38709 24409 38743
rect 24409 38709 24443 38743
rect 24443 38709 24452 38743
rect 24400 38700 24452 38709
rect 3917 38598 3969 38650
rect 3981 38598 4033 38650
rect 4045 38598 4097 38650
rect 4109 38598 4161 38650
rect 4173 38598 4225 38650
rect 9851 38598 9903 38650
rect 9915 38598 9967 38650
rect 9979 38598 10031 38650
rect 10043 38598 10095 38650
rect 10107 38598 10159 38650
rect 15785 38598 15837 38650
rect 15849 38598 15901 38650
rect 15913 38598 15965 38650
rect 15977 38598 16029 38650
rect 16041 38598 16093 38650
rect 21719 38598 21771 38650
rect 21783 38598 21835 38650
rect 21847 38598 21899 38650
rect 21911 38598 21963 38650
rect 21975 38598 22027 38650
rect 5356 38496 5408 38548
rect 9220 38496 9272 38548
rect 6000 38471 6052 38480
rect 6000 38437 6009 38471
rect 6009 38437 6043 38471
rect 6043 38437 6052 38471
rect 6000 38428 6052 38437
rect 1768 38292 1820 38344
rect 756 38224 808 38276
rect 2228 38267 2280 38276
rect 2228 38233 2237 38267
rect 2237 38233 2271 38267
rect 2271 38233 2280 38267
rect 2228 38224 2280 38233
rect 1216 38156 1268 38208
rect 2872 38224 2924 38276
rect 3700 38224 3752 38276
rect 5172 38292 5224 38344
rect 5356 38335 5408 38344
rect 5356 38301 5365 38335
rect 5365 38301 5399 38335
rect 5399 38301 5408 38335
rect 5356 38292 5408 38301
rect 5540 38335 5592 38344
rect 5540 38301 5549 38335
rect 5549 38301 5583 38335
rect 5583 38301 5592 38335
rect 5540 38292 5592 38301
rect 6276 38335 6328 38344
rect 6276 38301 6285 38335
rect 6285 38301 6319 38335
rect 6319 38301 6328 38335
rect 6276 38292 6328 38301
rect 6552 38335 6604 38344
rect 6552 38301 6561 38335
rect 6561 38301 6595 38335
rect 6595 38301 6604 38335
rect 6552 38292 6604 38301
rect 8484 38292 8536 38344
rect 8852 38292 8904 38344
rect 9404 38305 9456 38344
rect 5448 38224 5500 38276
rect 9404 38292 9429 38305
rect 9429 38292 9456 38305
rect 11152 38292 11204 38344
rect 11612 38428 11664 38480
rect 12532 38496 12584 38548
rect 13268 38539 13320 38548
rect 13268 38505 13277 38539
rect 13277 38505 13311 38539
rect 13311 38505 13320 38539
rect 13268 38496 13320 38505
rect 20628 38496 20680 38548
rect 21180 38496 21232 38548
rect 23572 38496 23624 38548
rect 23756 38496 23808 38548
rect 11980 38360 12032 38412
rect 12164 38360 12216 38412
rect 20720 38360 20772 38412
rect 23112 38360 23164 38412
rect 4344 38156 4396 38208
rect 4436 38156 4488 38208
rect 4712 38156 4764 38208
rect 4804 38199 4856 38208
rect 4804 38165 4813 38199
rect 4813 38165 4847 38199
rect 4847 38165 4856 38199
rect 4804 38156 4856 38165
rect 4896 38156 4948 38208
rect 10140 38199 10192 38208
rect 10140 38165 10149 38199
rect 10149 38165 10183 38199
rect 10183 38165 10192 38199
rect 10140 38156 10192 38165
rect 12440 38335 12492 38344
rect 12440 38301 12474 38335
rect 12474 38301 12492 38335
rect 12440 38292 12492 38301
rect 12624 38335 12676 38344
rect 12624 38301 12633 38335
rect 12633 38301 12667 38335
rect 12667 38301 12676 38335
rect 12624 38292 12676 38301
rect 20076 38335 20128 38344
rect 20076 38301 20085 38335
rect 20085 38301 20119 38335
rect 20119 38301 20128 38335
rect 20076 38292 20128 38301
rect 22100 38335 22152 38344
rect 22100 38301 22109 38335
rect 22109 38301 22143 38335
rect 22143 38301 22152 38335
rect 22100 38292 22152 38301
rect 22652 38335 22704 38344
rect 22652 38301 22661 38335
rect 22661 38301 22695 38335
rect 22695 38301 22704 38335
rect 22652 38292 22704 38301
rect 23204 38335 23256 38344
rect 23204 38301 23213 38335
rect 23213 38301 23247 38335
rect 23247 38301 23256 38335
rect 23204 38292 23256 38301
rect 23296 38292 23348 38344
rect 11796 38156 11848 38208
rect 12164 38156 12216 38208
rect 22192 38199 22244 38208
rect 22192 38165 22201 38199
rect 22201 38165 22235 38199
rect 22235 38165 22244 38199
rect 22192 38156 22244 38165
rect 22836 38156 22888 38208
rect 22928 38199 22980 38208
rect 22928 38165 22937 38199
rect 22937 38165 22971 38199
rect 22971 38165 22980 38199
rect 22928 38156 22980 38165
rect 23388 38224 23440 38276
rect 23940 38335 23992 38344
rect 23940 38301 23949 38335
rect 23949 38301 23983 38335
rect 23983 38301 23992 38335
rect 23940 38292 23992 38301
rect 25228 38156 25280 38208
rect 6884 38054 6936 38106
rect 6948 38054 7000 38106
rect 7012 38054 7064 38106
rect 7076 38054 7128 38106
rect 7140 38054 7192 38106
rect 12818 38054 12870 38106
rect 12882 38054 12934 38106
rect 12946 38054 12998 38106
rect 13010 38054 13062 38106
rect 13074 38054 13126 38106
rect 18752 38054 18804 38106
rect 18816 38054 18868 38106
rect 18880 38054 18932 38106
rect 18944 38054 18996 38106
rect 19008 38054 19060 38106
rect 24686 38054 24738 38106
rect 24750 38054 24802 38106
rect 24814 38054 24866 38106
rect 24878 38054 24930 38106
rect 24942 38054 24994 38106
rect 3608 37884 3660 37936
rect 4804 37952 4856 38004
rect 4988 37952 5040 38004
rect 6552 37952 6604 38004
rect 8576 37884 8628 37936
rect 8944 37927 8996 37936
rect 8944 37893 8953 37927
rect 8953 37893 8987 37927
rect 8987 37893 8996 37927
rect 8944 37884 8996 37893
rect 9220 37927 9272 37936
rect 9220 37893 9229 37927
rect 9229 37893 9263 37927
rect 9263 37893 9272 37927
rect 9220 37884 9272 37893
rect 10140 37952 10192 38004
rect 12624 37952 12676 38004
rect 14464 37952 14516 38004
rect 22100 37952 22152 38004
rect 22192 37952 22244 38004
rect 1400 37859 1452 37868
rect 1400 37825 1409 37859
rect 1409 37825 1443 37859
rect 1443 37825 1452 37859
rect 1400 37816 1452 37825
rect 1216 37748 1268 37800
rect 4160 37816 4212 37868
rect 4344 37816 4396 37868
rect 4712 37816 4764 37868
rect 4988 37859 5040 37868
rect 4988 37825 4997 37859
rect 4997 37825 5031 37859
rect 5031 37825 5040 37859
rect 4988 37816 5040 37825
rect 5356 37816 5408 37868
rect 5724 37816 5776 37868
rect 6552 37816 6604 37868
rect 6736 37816 6788 37868
rect 9680 37859 9732 37868
rect 9680 37825 9689 37859
rect 9689 37825 9723 37859
rect 9723 37825 9732 37859
rect 9680 37816 9732 37825
rect 11152 37884 11204 37936
rect 1676 37791 1728 37800
rect 1676 37757 1685 37791
rect 1685 37757 1719 37791
rect 1719 37757 1728 37791
rect 1676 37748 1728 37757
rect 1768 37748 1820 37800
rect 6184 37748 6236 37800
rect 6368 37791 6420 37800
rect 6368 37757 6377 37791
rect 6377 37757 6411 37791
rect 6411 37757 6420 37791
rect 6368 37748 6420 37757
rect 7104 37748 7156 37800
rect 7564 37748 7616 37800
rect 9128 37748 9180 37800
rect 10324 37816 10376 37868
rect 13544 37816 13596 37868
rect 15476 37816 15528 37868
rect 22468 37884 22520 37936
rect 22928 37952 22980 38004
rect 23112 37952 23164 38004
rect 24032 37859 24084 37868
rect 24032 37825 24041 37859
rect 24041 37825 24075 37859
rect 24075 37825 24084 37859
rect 24032 37816 24084 37825
rect 6276 37680 6328 37732
rect 6000 37612 6052 37664
rect 10600 37612 10652 37664
rect 11520 37680 11572 37732
rect 19524 37748 19576 37800
rect 10968 37612 11020 37664
rect 11796 37612 11848 37664
rect 20168 37680 20220 37732
rect 13912 37612 13964 37664
rect 22836 37723 22888 37732
rect 22836 37689 22845 37723
rect 22845 37689 22879 37723
rect 22879 37689 22888 37723
rect 22836 37680 22888 37689
rect 22560 37612 22612 37664
rect 22928 37612 22980 37664
rect 24400 37655 24452 37664
rect 24400 37621 24409 37655
rect 24409 37621 24443 37655
rect 24443 37621 24452 37655
rect 24400 37612 24452 37621
rect 25044 37612 25096 37664
rect 3917 37510 3969 37562
rect 3981 37510 4033 37562
rect 4045 37510 4097 37562
rect 4109 37510 4161 37562
rect 4173 37510 4225 37562
rect 9851 37510 9903 37562
rect 9915 37510 9967 37562
rect 9979 37510 10031 37562
rect 10043 37510 10095 37562
rect 10107 37510 10159 37562
rect 15785 37510 15837 37562
rect 15849 37510 15901 37562
rect 15913 37510 15965 37562
rect 15977 37510 16029 37562
rect 16041 37510 16093 37562
rect 21719 37510 21771 37562
rect 21783 37510 21835 37562
rect 21847 37510 21899 37562
rect 21911 37510 21963 37562
rect 21975 37510 22027 37562
rect 3424 37451 3476 37460
rect 3424 37417 3433 37451
rect 3433 37417 3467 37451
rect 3467 37417 3476 37451
rect 3424 37408 3476 37417
rect 3884 37408 3936 37460
rect 4988 37408 5040 37460
rect 6184 37408 6236 37460
rect 7472 37408 7524 37460
rect 7564 37340 7616 37392
rect 848 37272 900 37324
rect 2136 37272 2188 37324
rect 1032 37204 1084 37256
rect 3424 37272 3476 37324
rect 1492 37136 1544 37188
rect 2228 37179 2280 37188
rect 2228 37145 2237 37179
rect 2237 37145 2271 37179
rect 2271 37145 2280 37179
rect 2228 37136 2280 37145
rect 2780 37179 2832 37188
rect 2780 37145 2789 37179
rect 2789 37145 2823 37179
rect 2823 37145 2832 37179
rect 2780 37136 2832 37145
rect 2872 37136 2924 37188
rect 1308 37068 1360 37120
rect 4068 37179 4120 37188
rect 4068 37145 4077 37179
rect 4077 37145 4111 37179
rect 4111 37145 4120 37179
rect 4068 37136 4120 37145
rect 7288 37272 7340 37324
rect 4804 37136 4856 37188
rect 4988 37247 5040 37256
rect 4988 37213 4995 37247
rect 4995 37213 5029 37247
rect 5029 37213 5040 37247
rect 4988 37204 5040 37213
rect 5448 37204 5500 37256
rect 5540 37136 5592 37188
rect 3700 37068 3752 37120
rect 4896 37068 4948 37120
rect 5724 37111 5776 37120
rect 5724 37077 5733 37111
rect 5733 37077 5767 37111
rect 5767 37077 5776 37111
rect 5724 37068 5776 37077
rect 6736 37068 6788 37120
rect 8484 37247 8536 37256
rect 8484 37213 8493 37247
rect 8493 37213 8527 37247
rect 8527 37213 8536 37247
rect 8484 37204 8536 37213
rect 10048 37315 10100 37324
rect 10048 37281 10057 37315
rect 10057 37281 10091 37315
rect 10091 37281 10100 37315
rect 10048 37272 10100 37281
rect 20076 37408 20128 37460
rect 22652 37408 22704 37460
rect 23388 37408 23440 37460
rect 11796 37340 11848 37392
rect 23204 37340 23256 37392
rect 13728 37272 13780 37324
rect 8668 37204 8720 37256
rect 20260 37204 20312 37256
rect 20536 37204 20588 37256
rect 20720 37247 20772 37256
rect 20720 37213 20729 37247
rect 20729 37213 20763 37247
rect 20763 37213 20772 37247
rect 20720 37204 20772 37213
rect 21824 37247 21876 37256
rect 21824 37213 21833 37247
rect 21833 37213 21867 37247
rect 21867 37213 21876 37247
rect 21824 37204 21876 37213
rect 8116 37068 8168 37120
rect 11060 37111 11112 37120
rect 11060 37077 11069 37111
rect 11069 37077 11103 37111
rect 11103 37077 11112 37111
rect 11060 37068 11112 37077
rect 21916 37136 21968 37188
rect 24124 37315 24176 37324
rect 24124 37281 24133 37315
rect 24133 37281 24167 37315
rect 24167 37281 24176 37315
rect 24124 37272 24176 37281
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 22192 37136 22244 37188
rect 23112 37204 23164 37256
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 23664 37204 23716 37256
rect 24216 37204 24268 37256
rect 22928 37068 22980 37120
rect 23848 37179 23900 37188
rect 23848 37145 23857 37179
rect 23857 37145 23891 37179
rect 23891 37145 23900 37179
rect 23848 37136 23900 37145
rect 6884 36966 6936 37018
rect 6948 36966 7000 37018
rect 7012 36966 7064 37018
rect 7076 36966 7128 37018
rect 7140 36966 7192 37018
rect 12818 36966 12870 37018
rect 12882 36966 12934 37018
rect 12946 36966 12998 37018
rect 13010 36966 13062 37018
rect 13074 36966 13126 37018
rect 18752 36966 18804 37018
rect 18816 36966 18868 37018
rect 18880 36966 18932 37018
rect 18944 36966 18996 37018
rect 19008 36966 19060 37018
rect 24686 36966 24738 37018
rect 24750 36966 24802 37018
rect 24814 36966 24866 37018
rect 24878 36966 24930 37018
rect 24942 36966 24994 37018
rect 480 36864 532 36916
rect 3700 36864 3752 36916
rect 3424 36839 3476 36848
rect 3424 36805 3433 36839
rect 3433 36805 3467 36839
rect 3467 36805 3476 36839
rect 3424 36796 3476 36805
rect 3608 36796 3660 36848
rect 2780 36728 2832 36780
rect 4252 36796 4304 36848
rect 4804 36796 4856 36848
rect 4344 36728 4396 36780
rect 4620 36728 4672 36780
rect 4712 36728 4764 36780
rect 5816 36796 5868 36848
rect 8484 36864 8536 36916
rect 8576 36864 8628 36916
rect 20720 36864 20772 36916
rect 21824 36864 21876 36916
rect 21916 36864 21968 36916
rect 6920 36771 6972 36780
rect 6920 36737 6929 36771
rect 6929 36737 6963 36771
rect 6963 36737 6972 36771
rect 6920 36728 6972 36737
rect 7288 36728 7340 36780
rect 7380 36771 7432 36780
rect 7380 36737 7389 36771
rect 7389 36737 7423 36771
rect 7423 36737 7432 36771
rect 7380 36728 7432 36737
rect 7656 36728 7708 36780
rect 480 36660 532 36712
rect 940 36524 992 36576
rect 4896 36703 4948 36712
rect 4896 36669 4905 36703
rect 4905 36669 4939 36703
rect 4939 36669 4948 36703
rect 4896 36660 4948 36669
rect 9128 36728 9180 36780
rect 16672 36728 16724 36780
rect 8484 36660 8536 36712
rect 8668 36660 8720 36712
rect 10048 36660 10100 36712
rect 10416 36660 10468 36712
rect 7288 36592 7340 36644
rect 2320 36524 2372 36576
rect 5632 36524 5684 36576
rect 6736 36524 6788 36576
rect 9772 36592 9824 36644
rect 10784 36592 10836 36644
rect 8392 36524 8444 36576
rect 19248 36728 19300 36780
rect 20260 36771 20312 36780
rect 20260 36737 20269 36771
rect 20269 36737 20303 36771
rect 20303 36737 20312 36771
rect 20260 36728 20312 36737
rect 20536 36771 20588 36780
rect 20536 36737 20545 36771
rect 20545 36737 20579 36771
rect 20579 36737 20588 36771
rect 20536 36728 20588 36737
rect 20720 36728 20772 36780
rect 23848 36864 23900 36916
rect 24032 36864 24084 36916
rect 12532 36567 12584 36576
rect 12532 36533 12541 36567
rect 12541 36533 12575 36567
rect 12575 36533 12584 36567
rect 12532 36524 12584 36533
rect 17132 36524 17184 36576
rect 17408 36524 17460 36576
rect 17960 36524 18012 36576
rect 20720 36524 20772 36576
rect 21088 36524 21140 36576
rect 23112 36796 23164 36848
rect 23020 36771 23072 36780
rect 23020 36737 23029 36771
rect 23029 36737 23063 36771
rect 23063 36737 23072 36771
rect 23020 36728 23072 36737
rect 24032 36728 24084 36780
rect 22376 36660 22428 36712
rect 24492 36728 24544 36780
rect 23480 36592 23532 36644
rect 22836 36567 22888 36576
rect 22836 36533 22845 36567
rect 22845 36533 22879 36567
rect 22879 36533 22888 36567
rect 22836 36524 22888 36533
rect 24400 36567 24452 36576
rect 24400 36533 24409 36567
rect 24409 36533 24443 36567
rect 24443 36533 24452 36567
rect 24400 36524 24452 36533
rect 3917 36422 3969 36474
rect 3981 36422 4033 36474
rect 4045 36422 4097 36474
rect 4109 36422 4161 36474
rect 4173 36422 4225 36474
rect 9851 36422 9903 36474
rect 9915 36422 9967 36474
rect 9979 36422 10031 36474
rect 10043 36422 10095 36474
rect 10107 36422 10159 36474
rect 15785 36422 15837 36474
rect 15849 36422 15901 36474
rect 15913 36422 15965 36474
rect 15977 36422 16029 36474
rect 16041 36422 16093 36474
rect 21719 36422 21771 36474
rect 21783 36422 21835 36474
rect 21847 36422 21899 36474
rect 21911 36422 21963 36474
rect 21975 36422 22027 36474
rect 6920 36320 6972 36372
rect 11060 36320 11112 36372
rect 17132 36320 17184 36372
rect 21088 36320 21140 36372
rect 22376 36363 22428 36372
rect 22376 36329 22385 36363
rect 22385 36329 22419 36363
rect 22419 36329 22428 36363
rect 22376 36320 22428 36329
rect 22836 36320 22888 36372
rect 23572 36320 23624 36372
rect 1308 36116 1360 36168
rect 3884 36252 3936 36304
rect 4896 36252 4948 36304
rect 2780 36184 2832 36236
rect 5724 36295 5776 36304
rect 5724 36261 5733 36295
rect 5733 36261 5767 36295
rect 5767 36261 5776 36295
rect 5724 36252 5776 36261
rect 7288 36252 7340 36304
rect 2964 36116 3016 36168
rect 3792 36159 3844 36168
rect 3792 36125 3801 36159
rect 3801 36125 3835 36159
rect 3835 36125 3844 36159
rect 3792 36116 3844 36125
rect 4804 36116 4856 36168
rect 5172 36116 5224 36168
rect 7380 36184 7432 36236
rect 11244 36227 11296 36236
rect 11244 36193 11253 36227
rect 11253 36193 11287 36227
rect 11287 36193 11296 36227
rect 11244 36184 11296 36193
rect 388 36048 440 36100
rect 1860 36048 1912 36100
rect 2412 36048 2464 36100
rect 4068 36091 4120 36100
rect 4068 36057 4077 36091
rect 4077 36057 4111 36091
rect 4111 36057 4120 36091
rect 4068 36048 4120 36057
rect 2688 35980 2740 36032
rect 3424 35980 3476 36032
rect 4712 35980 4764 36032
rect 5172 35980 5224 36032
rect 5448 36116 5500 36168
rect 6000 36159 6052 36168
rect 6000 36125 6009 36159
rect 6009 36125 6043 36159
rect 6043 36125 6052 36159
rect 6000 36116 6052 36125
rect 6092 36159 6144 36168
rect 6092 36125 6126 36159
rect 6126 36125 6144 36159
rect 6092 36116 6144 36125
rect 6276 36159 6328 36168
rect 6276 36125 6285 36159
rect 6285 36125 6319 36159
rect 6319 36125 6328 36159
rect 6276 36116 6328 36125
rect 7288 36116 7340 36168
rect 8300 36116 8352 36168
rect 8852 36116 8904 36168
rect 9128 36116 9180 36168
rect 9772 36116 9824 36168
rect 10508 36159 10560 36168
rect 10508 36125 10517 36159
rect 10517 36125 10551 36159
rect 10551 36125 10560 36159
rect 10508 36116 10560 36125
rect 11336 36159 11388 36168
rect 12532 36184 12584 36236
rect 11336 36125 11370 36159
rect 11370 36125 11388 36159
rect 11336 36116 11388 36125
rect 17224 36116 17276 36168
rect 17868 36116 17920 36168
rect 20260 36252 20312 36304
rect 20812 36252 20864 36304
rect 17408 36091 17460 36100
rect 17408 36057 17420 36091
rect 17420 36057 17460 36091
rect 17408 36048 17460 36057
rect 17776 36048 17828 36100
rect 20536 36184 20588 36236
rect 5632 35980 5684 36032
rect 7564 35980 7616 36032
rect 8116 35980 8168 36032
rect 8576 35980 8628 36032
rect 11336 35980 11388 36032
rect 11612 35980 11664 36032
rect 12256 35980 12308 36032
rect 12624 35980 12676 36032
rect 19340 35980 19392 36032
rect 19800 35980 19852 36032
rect 23572 36159 23624 36168
rect 23572 36125 23581 36159
rect 23581 36125 23615 36159
rect 23615 36125 23624 36159
rect 23572 36116 23624 36125
rect 25136 36048 25188 36100
rect 6884 35878 6936 35930
rect 6948 35878 7000 35930
rect 7012 35878 7064 35930
rect 7076 35878 7128 35930
rect 7140 35878 7192 35930
rect 12818 35878 12870 35930
rect 12882 35878 12934 35930
rect 12946 35878 12998 35930
rect 13010 35878 13062 35930
rect 13074 35878 13126 35930
rect 18752 35878 18804 35930
rect 18816 35878 18868 35930
rect 18880 35878 18932 35930
rect 18944 35878 18996 35930
rect 19008 35878 19060 35930
rect 24686 35878 24738 35930
rect 24750 35878 24802 35930
rect 24814 35878 24866 35930
rect 24878 35878 24930 35930
rect 24942 35878 24994 35930
rect 3516 35776 3568 35828
rect 1860 35640 1912 35692
rect 2688 35683 2740 35692
rect 2688 35649 2697 35683
rect 2697 35649 2731 35683
rect 2731 35649 2740 35683
rect 2688 35640 2740 35649
rect 3424 35683 3476 35692
rect 3424 35649 3433 35683
rect 3433 35649 3467 35683
rect 3467 35649 3476 35683
rect 3424 35640 3476 35649
rect 7288 35776 7340 35828
rect 8944 35776 8996 35828
rect 9220 35776 9272 35828
rect 9588 35776 9640 35828
rect 11888 35776 11940 35828
rect 4528 35708 4580 35760
rect 6092 35708 6144 35760
rect 8576 35751 8628 35760
rect 8576 35717 8585 35751
rect 8585 35717 8619 35751
rect 8619 35717 8628 35751
rect 8576 35708 8628 35717
rect 2044 35572 2096 35624
rect 2136 35547 2188 35556
rect 2136 35513 2145 35547
rect 2145 35513 2179 35547
rect 2179 35513 2188 35547
rect 2136 35504 2188 35513
rect 1768 35436 1820 35488
rect 2044 35436 2096 35488
rect 3608 35615 3660 35624
rect 3608 35581 3617 35615
rect 3617 35581 3651 35615
rect 3651 35581 3660 35615
rect 3608 35572 3660 35581
rect 3884 35572 3936 35624
rect 3056 35436 3108 35488
rect 9404 35708 9456 35760
rect 8852 35640 8904 35692
rect 9680 35708 9732 35760
rect 4528 35615 4580 35624
rect 4528 35581 4537 35615
rect 4537 35581 4571 35615
rect 4571 35581 4580 35615
rect 4528 35572 4580 35581
rect 5264 35615 5316 35624
rect 5264 35581 5273 35615
rect 5273 35581 5307 35615
rect 5307 35581 5316 35615
rect 5264 35572 5316 35581
rect 5448 35572 5500 35624
rect 6276 35572 6328 35624
rect 8392 35572 8444 35624
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 4712 35504 4764 35556
rect 5724 35436 5776 35488
rect 5908 35436 5960 35488
rect 7472 35436 7524 35488
rect 9404 35436 9456 35488
rect 9588 35436 9640 35488
rect 11520 35708 11572 35760
rect 11704 35751 11756 35760
rect 11704 35717 11713 35751
rect 11713 35717 11747 35751
rect 11747 35717 11756 35751
rect 11704 35708 11756 35717
rect 11980 35751 12032 35760
rect 11980 35717 11989 35751
rect 11989 35717 12023 35751
rect 12023 35717 12032 35751
rect 11980 35708 12032 35717
rect 19340 35776 19392 35828
rect 12164 35708 12216 35760
rect 13820 35708 13872 35760
rect 18236 35708 18288 35760
rect 10416 35436 10468 35488
rect 11612 35640 11664 35692
rect 12624 35640 12676 35692
rect 12808 35572 12860 35624
rect 12992 35547 13044 35556
rect 12992 35513 13001 35547
rect 13001 35513 13035 35547
rect 13035 35513 13044 35547
rect 12992 35504 13044 35513
rect 11060 35436 11112 35488
rect 14188 35436 14240 35488
rect 15476 35436 15528 35488
rect 16856 35640 16908 35692
rect 17592 35615 17644 35624
rect 17592 35581 17601 35615
rect 17601 35581 17635 35615
rect 17635 35581 17644 35615
rect 17592 35572 17644 35581
rect 21272 35683 21324 35692
rect 21272 35649 21281 35683
rect 21281 35649 21315 35683
rect 21315 35649 21324 35683
rect 21272 35640 21324 35649
rect 23020 35776 23072 35828
rect 23572 35776 23624 35828
rect 25320 35708 25372 35760
rect 22376 35572 22428 35624
rect 23940 35683 23992 35692
rect 23940 35649 23949 35683
rect 23949 35649 23983 35683
rect 23983 35649 23992 35683
rect 23940 35640 23992 35649
rect 19064 35479 19116 35488
rect 19064 35445 19073 35479
rect 19073 35445 19107 35479
rect 19107 35445 19116 35479
rect 19064 35436 19116 35445
rect 21180 35436 21232 35488
rect 23756 35479 23808 35488
rect 23756 35445 23765 35479
rect 23765 35445 23799 35479
rect 23799 35445 23808 35479
rect 23756 35436 23808 35445
rect 24400 35479 24452 35488
rect 24400 35445 24409 35479
rect 24409 35445 24443 35479
rect 24443 35445 24452 35479
rect 24400 35436 24452 35445
rect 3917 35334 3969 35386
rect 3981 35334 4033 35386
rect 4045 35334 4097 35386
rect 4109 35334 4161 35386
rect 4173 35334 4225 35386
rect 9851 35334 9903 35386
rect 9915 35334 9967 35386
rect 9979 35334 10031 35386
rect 10043 35334 10095 35386
rect 10107 35334 10159 35386
rect 15785 35334 15837 35386
rect 15849 35334 15901 35386
rect 15913 35334 15965 35386
rect 15977 35334 16029 35386
rect 16041 35334 16093 35386
rect 21719 35334 21771 35386
rect 21783 35334 21835 35386
rect 21847 35334 21899 35386
rect 21911 35334 21963 35386
rect 21975 35334 22027 35386
rect 3240 35232 3292 35284
rect 5540 35232 5592 35284
rect 6184 35232 6236 35284
rect 6276 35232 6328 35284
rect 5264 35096 5316 35148
rect 756 35028 808 35080
rect 2320 35071 2372 35080
rect 2320 35037 2329 35071
rect 2329 35037 2363 35071
rect 2363 35037 2372 35071
rect 2320 35028 2372 35037
rect 2504 35028 2556 35080
rect 3240 35028 3292 35080
rect 4252 35071 4304 35080
rect 4252 35037 4261 35071
rect 4261 35037 4295 35071
rect 4295 35037 4304 35071
rect 4252 35028 4304 35037
rect 5724 35071 5776 35080
rect 5724 35037 5731 35071
rect 5731 35037 5765 35071
rect 5765 35037 5776 35071
rect 9588 35232 9640 35284
rect 10416 35232 10468 35284
rect 7932 35164 7984 35216
rect 7288 35096 7340 35148
rect 10416 35096 10468 35148
rect 11060 35232 11112 35284
rect 12808 35275 12860 35284
rect 12808 35241 12817 35275
rect 12817 35241 12851 35275
rect 12851 35241 12860 35275
rect 12808 35232 12860 35241
rect 13544 35232 13596 35284
rect 13820 35164 13872 35216
rect 11612 35096 11664 35148
rect 15476 35096 15528 35148
rect 19064 35232 19116 35284
rect 16672 35207 16724 35216
rect 16672 35173 16681 35207
rect 16681 35173 16715 35207
rect 16715 35173 16724 35207
rect 16672 35164 16724 35173
rect 17132 35164 17184 35216
rect 17592 35164 17644 35216
rect 19984 35232 20036 35284
rect 22284 35232 22336 35284
rect 23664 35232 23716 35284
rect 24584 35232 24636 35284
rect 20628 35164 20680 35216
rect 21180 35096 21232 35148
rect 5724 35028 5776 35037
rect 8944 35028 8996 35080
rect 9772 35028 9824 35080
rect 10784 35071 10836 35080
rect 10784 35037 10793 35071
rect 10793 35037 10827 35071
rect 10827 35037 10836 35071
rect 10784 35028 10836 35037
rect 11060 35071 11112 35080
rect 11060 35037 11069 35071
rect 11069 35037 11103 35071
rect 11103 35037 11112 35071
rect 11060 35028 11112 35037
rect 12072 35071 12124 35080
rect 4344 35003 4396 35012
rect 4344 34969 4353 35003
rect 4353 34969 4387 35003
rect 4387 34969 4396 35003
rect 4344 34960 4396 34969
rect 4620 34960 4672 35012
rect 3332 34892 3384 34944
rect 3792 34892 3844 34944
rect 4436 34892 4488 34944
rect 5264 34960 5316 35012
rect 5172 34892 5224 34944
rect 7564 34960 7616 35012
rect 12072 35037 12079 35071
rect 12079 35037 12113 35071
rect 12113 35037 12124 35071
rect 12072 35028 12124 35037
rect 14188 34960 14240 35012
rect 5816 34892 5868 34944
rect 14464 34892 14516 34944
rect 17960 35028 18012 35080
rect 18236 35028 18288 35080
rect 19340 35028 19392 35080
rect 16396 34960 16448 35012
rect 19248 34960 19300 35012
rect 19432 34960 19484 35012
rect 19616 34892 19668 34944
rect 22284 35096 22336 35148
rect 22652 35096 22704 35148
rect 23388 35071 23440 35080
rect 23388 35037 23397 35071
rect 23397 35037 23431 35071
rect 23431 35037 23440 35071
rect 23388 35028 23440 35037
rect 20628 34960 20680 35012
rect 24216 34960 24268 35012
rect 23480 34935 23532 34944
rect 23480 34901 23489 34935
rect 23489 34901 23523 34935
rect 23523 34901 23532 34935
rect 23480 34892 23532 34901
rect 25228 34892 25280 34944
rect 6884 34790 6936 34842
rect 6948 34790 7000 34842
rect 7012 34790 7064 34842
rect 7076 34790 7128 34842
rect 7140 34790 7192 34842
rect 12818 34790 12870 34842
rect 12882 34790 12934 34842
rect 12946 34790 12998 34842
rect 13010 34790 13062 34842
rect 13074 34790 13126 34842
rect 18752 34790 18804 34842
rect 18816 34790 18868 34842
rect 18880 34790 18932 34842
rect 18944 34790 18996 34842
rect 19008 34790 19060 34842
rect 24686 34790 24738 34842
rect 24750 34790 24802 34842
rect 24814 34790 24866 34842
rect 24878 34790 24930 34842
rect 24942 34790 24994 34842
rect 2136 34688 2188 34740
rect 2596 34688 2648 34740
rect 2780 34688 2832 34740
rect 3608 34620 3660 34672
rect 3976 34620 4028 34672
rect 4344 34688 4396 34740
rect 4620 34688 4672 34740
rect 9036 34731 9088 34740
rect 9036 34697 9045 34731
rect 9045 34697 9079 34731
rect 9079 34697 9088 34731
rect 9036 34688 9088 34697
rect 14188 34688 14240 34740
rect 15292 34688 15344 34740
rect 15384 34688 15436 34740
rect 19432 34688 19484 34740
rect 2412 34552 2464 34604
rect 2780 34595 2832 34604
rect 2780 34561 2789 34595
rect 2789 34561 2823 34595
rect 2823 34561 2832 34595
rect 2780 34552 2832 34561
rect 3332 34552 3384 34604
rect 4160 34552 4212 34604
rect 5540 34552 5592 34604
rect 6644 34595 6696 34604
rect 6644 34561 6653 34595
rect 6653 34561 6696 34595
rect 6644 34552 6696 34561
rect 9680 34620 9732 34672
rect 8484 34552 8536 34604
rect 1400 34527 1452 34536
rect 1400 34493 1409 34527
rect 1409 34493 1443 34527
rect 1443 34493 1452 34527
rect 1400 34484 1452 34493
rect 5908 34484 5960 34536
rect 6184 34484 6236 34536
rect 1768 34348 1820 34400
rect 5172 34348 5224 34400
rect 7380 34391 7432 34400
rect 7380 34357 7389 34391
rect 7389 34357 7423 34391
rect 7423 34357 7432 34391
rect 7380 34348 7432 34357
rect 9496 34595 9548 34604
rect 9496 34561 9505 34595
rect 9505 34561 9539 34595
rect 9539 34561 9548 34595
rect 9496 34552 9548 34561
rect 9588 34595 9640 34604
rect 9588 34561 9597 34595
rect 9597 34561 9631 34595
rect 9631 34561 9640 34595
rect 9588 34552 9640 34561
rect 10692 34552 10744 34604
rect 16672 34620 16724 34672
rect 16764 34620 16816 34672
rect 14832 34552 14884 34604
rect 15016 34552 15068 34604
rect 17132 34620 17184 34672
rect 19340 34663 19392 34672
rect 17500 34595 17552 34604
rect 17500 34561 17509 34595
rect 17509 34561 17543 34595
rect 17543 34561 17552 34595
rect 17500 34552 17552 34561
rect 17868 34552 17920 34604
rect 18972 34595 19024 34604
rect 18972 34561 18981 34595
rect 18981 34561 19015 34595
rect 19015 34561 19024 34595
rect 18972 34552 19024 34561
rect 19340 34629 19374 34663
rect 19374 34629 19392 34663
rect 19340 34620 19392 34629
rect 19616 34620 19668 34672
rect 20444 34620 20496 34672
rect 22192 34552 22244 34604
rect 23296 34688 23348 34740
rect 23664 34731 23716 34740
rect 23664 34697 23673 34731
rect 23673 34697 23707 34731
rect 23707 34697 23716 34731
rect 23664 34688 23716 34697
rect 23756 34688 23808 34740
rect 23940 34620 23992 34672
rect 11888 34484 11940 34536
rect 13912 34484 13964 34536
rect 11704 34416 11756 34468
rect 9772 34348 9824 34400
rect 11060 34391 11112 34400
rect 11060 34357 11069 34391
rect 11069 34357 11103 34391
rect 11103 34357 11112 34391
rect 11060 34348 11112 34357
rect 19064 34527 19116 34536
rect 17224 34416 17276 34468
rect 19064 34493 19073 34527
rect 19073 34493 19107 34527
rect 19107 34493 19116 34527
rect 19064 34484 19116 34493
rect 21088 34484 21140 34536
rect 24400 34527 24452 34536
rect 24400 34493 24409 34527
rect 24409 34493 24443 34527
rect 24443 34493 24452 34527
rect 24400 34484 24452 34493
rect 15016 34348 15068 34400
rect 19800 34348 19852 34400
rect 19984 34348 20036 34400
rect 20444 34391 20496 34400
rect 20444 34357 20453 34391
rect 20453 34357 20487 34391
rect 20487 34357 20496 34391
rect 20444 34348 20496 34357
rect 20812 34391 20864 34400
rect 20812 34357 20821 34391
rect 20821 34357 20855 34391
rect 20855 34357 20864 34391
rect 20812 34348 20864 34357
rect 23112 34348 23164 34400
rect 3917 34246 3969 34298
rect 3981 34246 4033 34298
rect 4045 34246 4097 34298
rect 4109 34246 4161 34298
rect 4173 34246 4225 34298
rect 9851 34246 9903 34298
rect 9915 34246 9967 34298
rect 9979 34246 10031 34298
rect 10043 34246 10095 34298
rect 10107 34246 10159 34298
rect 15785 34246 15837 34298
rect 15849 34246 15901 34298
rect 15913 34246 15965 34298
rect 15977 34246 16029 34298
rect 16041 34246 16093 34298
rect 21719 34246 21771 34298
rect 21783 34246 21835 34298
rect 21847 34246 21899 34298
rect 21911 34246 21963 34298
rect 21975 34246 22027 34298
rect 204 34144 256 34196
rect 1768 34144 1820 34196
rect 2964 34144 3016 34196
rect 5540 34144 5592 34196
rect 756 33940 808 33992
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 6460 34008 6512 34060
rect 6828 34051 6880 34060
rect 6828 34017 6837 34051
rect 6837 34017 6871 34051
rect 6871 34017 6880 34051
rect 6828 34008 6880 34017
rect 9404 34144 9456 34196
rect 7380 34076 7432 34128
rect 8484 34076 8536 34128
rect 9772 34144 9824 34196
rect 16212 34144 16264 34196
rect 17500 34144 17552 34196
rect 2780 33983 2832 33992
rect 2780 33949 2789 33983
rect 2789 33949 2823 33983
rect 2823 33949 2832 33983
rect 2780 33940 2832 33949
rect 1308 33872 1360 33924
rect 4068 33915 4120 33924
rect 4068 33881 4077 33915
rect 4077 33881 4111 33915
rect 4111 33881 4120 33915
rect 4068 33872 4120 33881
rect 5264 33940 5316 33992
rect 6368 33940 6420 33992
rect 4896 33872 4948 33924
rect 6184 33872 6236 33924
rect 8024 33983 8076 33992
rect 8024 33949 8033 33983
rect 8033 33949 8067 33983
rect 8067 33949 8076 33983
rect 8024 33940 8076 33949
rect 10692 34076 10744 34128
rect 10784 34076 10836 34128
rect 13728 34076 13780 34128
rect 16764 34076 16816 34128
rect 20536 34144 20588 34196
rect 20812 34144 20864 34196
rect 21088 34187 21140 34196
rect 21088 34153 21097 34187
rect 21097 34153 21131 34187
rect 21131 34153 21140 34187
rect 21088 34144 21140 34153
rect 23388 34144 23440 34196
rect 8852 34008 8904 34060
rect 11612 34008 11664 34060
rect 11888 34008 11940 34060
rect 12532 34051 12584 34060
rect 12532 34017 12541 34051
rect 12541 34017 12575 34051
rect 12575 34017 12584 34051
rect 12532 34008 12584 34017
rect 15200 34008 15252 34060
rect 15476 34008 15528 34060
rect 17316 34008 17368 34060
rect 13544 33940 13596 33992
rect 13912 33940 13964 33992
rect 296 33804 348 33856
rect 572 33804 624 33856
rect 1768 33804 1820 33856
rect 5540 33847 5592 33856
rect 5540 33813 5549 33847
rect 5549 33813 5583 33847
rect 5583 33813 5592 33847
rect 5540 33804 5592 33813
rect 6460 33804 6512 33856
rect 8668 33847 8720 33856
rect 8668 33813 8677 33847
rect 8677 33813 8711 33847
rect 8711 33813 8720 33847
rect 8668 33804 8720 33813
rect 9496 33872 9548 33924
rect 12348 33872 12400 33924
rect 12624 33872 12676 33924
rect 14004 33872 14056 33924
rect 15384 33940 15436 33992
rect 16212 33983 16264 33992
rect 16212 33949 16219 33983
rect 16219 33949 16253 33983
rect 16253 33949 16264 33983
rect 16212 33940 16264 33949
rect 16856 33940 16908 33992
rect 17500 33983 17552 33992
rect 17500 33949 17509 33983
rect 17509 33949 17543 33983
rect 17543 33949 17552 33983
rect 17500 33940 17552 33949
rect 9404 33804 9456 33856
rect 17040 33872 17092 33924
rect 19524 33872 19576 33924
rect 19800 33940 19852 33992
rect 22560 33983 22612 33992
rect 22560 33949 22569 33983
rect 22569 33949 22603 33983
rect 22603 33949 22612 33983
rect 22560 33940 22612 33949
rect 22836 33983 22888 33992
rect 22836 33949 22845 33983
rect 22845 33949 22879 33983
rect 22879 33949 22888 33983
rect 22836 33940 22888 33949
rect 14280 33804 14332 33856
rect 15016 33804 15068 33856
rect 15108 33847 15160 33856
rect 15108 33813 15117 33847
rect 15117 33813 15151 33847
rect 15151 33813 15160 33847
rect 15108 33804 15160 33813
rect 16948 33847 17000 33856
rect 16948 33813 16957 33847
rect 16957 33813 16991 33847
rect 16991 33813 17000 33847
rect 16948 33804 17000 33813
rect 18236 33847 18288 33856
rect 18236 33813 18245 33847
rect 18245 33813 18279 33847
rect 18279 33813 18288 33847
rect 18236 33804 18288 33813
rect 19892 33804 19944 33856
rect 21640 33804 21692 33856
rect 22652 33847 22704 33856
rect 22652 33813 22661 33847
rect 22661 33813 22695 33847
rect 22695 33813 22704 33847
rect 22652 33804 22704 33813
rect 23480 33940 23532 33992
rect 23204 33872 23256 33924
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 25228 33804 25280 33856
rect 6884 33702 6936 33754
rect 6948 33702 7000 33754
rect 7012 33702 7064 33754
rect 7076 33702 7128 33754
rect 7140 33702 7192 33754
rect 12818 33702 12870 33754
rect 12882 33702 12934 33754
rect 12946 33702 12998 33754
rect 13010 33702 13062 33754
rect 13074 33702 13126 33754
rect 18752 33702 18804 33754
rect 18816 33702 18868 33754
rect 18880 33702 18932 33754
rect 18944 33702 18996 33754
rect 19008 33702 19060 33754
rect 24686 33702 24738 33754
rect 24750 33702 24802 33754
rect 24814 33702 24866 33754
rect 24878 33702 24930 33754
rect 24942 33702 24994 33754
rect 1216 33600 1268 33652
rect 2688 33600 2740 33652
rect 2964 33600 3016 33652
rect 3792 33600 3844 33652
rect 5172 33600 5224 33652
rect 7104 33600 7156 33652
rect 8668 33600 8720 33652
rect 9036 33600 9088 33652
rect 9588 33600 9640 33652
rect 11612 33600 11664 33652
rect 11796 33600 11848 33652
rect 12716 33600 12768 33652
rect 13728 33600 13780 33652
rect 14004 33600 14056 33652
rect 3056 33575 3108 33584
rect 3056 33541 3065 33575
rect 3065 33541 3099 33575
rect 3099 33541 3108 33575
rect 3056 33532 3108 33541
rect 1400 33396 1452 33448
rect 3240 33464 3292 33516
rect 3424 33507 3476 33516
rect 3424 33473 3433 33507
rect 3433 33473 3467 33507
rect 3467 33473 3476 33507
rect 3424 33464 3476 33473
rect 3792 33507 3844 33516
rect 3792 33473 3801 33507
rect 3801 33473 3835 33507
rect 3835 33473 3844 33507
rect 3792 33464 3844 33473
rect 4528 33532 4580 33584
rect 4620 33464 4672 33516
rect 4344 33371 4396 33380
rect 4344 33337 4353 33371
rect 4353 33337 4387 33371
rect 4387 33337 4396 33371
rect 4344 33328 4396 33337
rect 2412 33260 2464 33312
rect 2688 33260 2740 33312
rect 4896 33507 4948 33516
rect 4896 33473 4905 33507
rect 4905 33473 4939 33507
rect 4939 33473 4948 33507
rect 4896 33464 4948 33473
rect 5356 33532 5408 33584
rect 7288 33464 7340 33516
rect 8116 33507 8168 33516
rect 8116 33473 8125 33507
rect 8125 33473 8159 33507
rect 8159 33473 8168 33507
rect 8116 33464 8168 33473
rect 10968 33532 11020 33584
rect 9772 33507 9824 33516
rect 6920 33439 6972 33448
rect 6920 33405 6929 33439
rect 6929 33405 6963 33439
rect 6963 33405 6972 33439
rect 6920 33396 6972 33405
rect 5172 33260 5224 33312
rect 5356 33260 5408 33312
rect 7196 33396 7248 33448
rect 7932 33439 7984 33448
rect 7932 33405 7966 33439
rect 7966 33405 7984 33439
rect 7932 33396 7984 33405
rect 7380 33328 7432 33380
rect 9772 33473 9797 33507
rect 9797 33473 9824 33507
rect 9772 33464 9824 33473
rect 9864 33464 9916 33516
rect 11060 33396 11112 33448
rect 12164 33464 12216 33516
rect 12716 33507 12768 33516
rect 12716 33473 12725 33507
rect 12725 33473 12759 33507
rect 12759 33473 12768 33507
rect 12716 33464 12768 33473
rect 13912 33464 13964 33516
rect 14372 33464 14424 33516
rect 15200 33507 15252 33516
rect 15200 33473 15209 33507
rect 15209 33473 15243 33507
rect 15243 33473 15252 33507
rect 15200 33464 15252 33473
rect 16764 33600 16816 33652
rect 16580 33532 16632 33584
rect 18236 33600 18288 33652
rect 17132 33507 17184 33516
rect 17132 33473 17141 33507
rect 17141 33473 17175 33507
rect 17175 33473 17184 33507
rect 17132 33464 17184 33473
rect 17224 33507 17276 33516
rect 17224 33473 17233 33507
rect 17233 33473 17267 33507
rect 17267 33473 17276 33507
rect 17224 33464 17276 33473
rect 17316 33464 17368 33516
rect 18972 33575 19024 33584
rect 18972 33541 18981 33575
rect 18981 33541 19015 33575
rect 19015 33541 19024 33575
rect 18972 33532 19024 33541
rect 18604 33396 18656 33448
rect 19156 33464 19208 33516
rect 19432 33464 19484 33516
rect 22652 33600 22704 33652
rect 22836 33600 22888 33652
rect 23664 33600 23716 33652
rect 20996 33464 21048 33516
rect 11520 33328 11572 33380
rect 12164 33328 12216 33380
rect 21548 33396 21600 33448
rect 10324 33260 10376 33312
rect 10508 33303 10560 33312
rect 10508 33269 10517 33303
rect 10517 33269 10551 33303
rect 10551 33269 10560 33303
rect 10508 33260 10560 33269
rect 12900 33260 12952 33312
rect 16212 33303 16264 33312
rect 16212 33269 16221 33303
rect 16221 33269 16255 33303
rect 16255 33269 16264 33303
rect 16212 33260 16264 33269
rect 19432 33328 19484 33380
rect 23112 33464 23164 33516
rect 20996 33260 21048 33312
rect 22192 33260 22244 33312
rect 23388 33303 23440 33312
rect 23388 33269 23397 33303
rect 23397 33269 23431 33303
rect 23431 33269 23440 33303
rect 23388 33260 23440 33269
rect 25412 33328 25464 33380
rect 24400 33303 24452 33312
rect 24400 33269 24409 33303
rect 24409 33269 24443 33303
rect 24443 33269 24452 33303
rect 24400 33260 24452 33269
rect 3917 33158 3969 33210
rect 3981 33158 4033 33210
rect 4045 33158 4097 33210
rect 4109 33158 4161 33210
rect 4173 33158 4225 33210
rect 9851 33158 9903 33210
rect 9915 33158 9967 33210
rect 9979 33158 10031 33210
rect 10043 33158 10095 33210
rect 10107 33158 10159 33210
rect 15785 33158 15837 33210
rect 15849 33158 15901 33210
rect 15913 33158 15965 33210
rect 15977 33158 16029 33210
rect 16041 33158 16093 33210
rect 21719 33158 21771 33210
rect 21783 33158 21835 33210
rect 21847 33158 21899 33210
rect 21911 33158 21963 33210
rect 21975 33158 22027 33210
rect 1400 32988 1452 33040
rect 3424 33056 3476 33108
rect 6368 33056 6420 33108
rect 8116 33056 8168 33108
rect 9404 32988 9456 33040
rect 3332 32920 3384 32972
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 4160 32920 4212 32972
rect 5540 32920 5592 32972
rect 6184 32920 6236 32972
rect 11060 33056 11112 33108
rect 1308 32716 1360 32768
rect 4528 32827 4580 32836
rect 4528 32793 4537 32827
rect 4537 32793 4571 32827
rect 4571 32793 4580 32827
rect 4528 32784 4580 32793
rect 4896 32716 4948 32768
rect 5264 32895 5316 32904
rect 5264 32861 5273 32895
rect 5273 32861 5307 32895
rect 5307 32861 5316 32895
rect 5264 32852 5316 32861
rect 5356 32895 5408 32904
rect 5356 32861 5365 32895
rect 5365 32861 5399 32895
rect 5399 32861 5408 32895
rect 5356 32852 5408 32861
rect 5448 32852 5500 32904
rect 5816 32852 5868 32904
rect 10508 32920 10560 32972
rect 10692 32920 10744 32972
rect 11336 32920 11388 32972
rect 11520 32920 11572 32972
rect 11888 32963 11940 32972
rect 11888 32929 11897 32963
rect 11897 32929 11931 32963
rect 11931 32929 11940 32963
rect 11888 32920 11940 32929
rect 12900 33099 12952 33108
rect 12900 33065 12909 33099
rect 12909 33065 12943 33099
rect 12943 33065 12952 33099
rect 12900 33056 12952 33065
rect 15108 33056 15160 33108
rect 15384 33056 15436 33108
rect 16120 33056 16172 33108
rect 18604 33099 18656 33108
rect 18604 33065 18613 33099
rect 18613 33065 18647 33099
rect 18647 33065 18656 33099
rect 18604 33056 18656 33065
rect 23388 33056 23440 33108
rect 17316 32920 17368 32972
rect 17592 32963 17644 32972
rect 17592 32929 17601 32963
rect 17601 32929 17635 32963
rect 17635 32929 17644 32963
rect 17592 32920 17644 32929
rect 7472 32895 7524 32904
rect 7472 32861 7479 32895
rect 7479 32861 7513 32895
rect 7513 32861 7524 32895
rect 7472 32852 7524 32861
rect 8116 32852 8168 32904
rect 9220 32852 9272 32904
rect 9772 32852 9824 32904
rect 11152 32895 11204 32904
rect 11152 32861 11161 32895
rect 11161 32861 11195 32895
rect 11195 32861 11204 32895
rect 11152 32852 11204 32861
rect 10140 32784 10192 32836
rect 12624 32852 12676 32904
rect 6184 32716 6236 32768
rect 12716 32784 12768 32836
rect 13544 32784 13596 32836
rect 14004 32716 14056 32768
rect 15016 32895 15068 32904
rect 15016 32861 15025 32895
rect 15025 32861 15059 32895
rect 15059 32861 15068 32895
rect 15016 32852 15068 32861
rect 15108 32895 15160 32904
rect 15108 32861 15142 32895
rect 15142 32861 15160 32895
rect 15108 32852 15160 32861
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 17408 32852 17460 32904
rect 17868 32895 17920 32904
rect 17868 32861 17877 32895
rect 17877 32861 17920 32895
rect 17868 32852 17920 32861
rect 16856 32784 16908 32836
rect 19708 32784 19760 32836
rect 15292 32716 15344 32768
rect 15384 32716 15436 32768
rect 22192 32895 22244 32904
rect 22192 32861 22201 32895
rect 22201 32861 22235 32895
rect 22235 32861 22244 32895
rect 22192 32852 22244 32861
rect 23204 32784 23256 32836
rect 23296 32784 23348 32836
rect 23940 32895 23992 32904
rect 23940 32861 23949 32895
rect 23949 32861 23983 32895
rect 23983 32861 23992 32895
rect 23940 32852 23992 32861
rect 25136 32784 25188 32836
rect 22652 32716 22704 32768
rect 25228 32716 25280 32768
rect 6884 32614 6936 32666
rect 6948 32614 7000 32666
rect 7012 32614 7064 32666
rect 7076 32614 7128 32666
rect 7140 32614 7192 32666
rect 12818 32614 12870 32666
rect 12882 32614 12934 32666
rect 12946 32614 12998 32666
rect 13010 32614 13062 32666
rect 13074 32614 13126 32666
rect 18752 32614 18804 32666
rect 18816 32614 18868 32666
rect 18880 32614 18932 32666
rect 18944 32614 18996 32666
rect 19008 32614 19060 32666
rect 24686 32614 24738 32666
rect 24750 32614 24802 32666
rect 24814 32614 24866 32666
rect 24878 32614 24930 32666
rect 24942 32614 24994 32666
rect 1216 32512 1268 32564
rect 3700 32444 3752 32496
rect 2320 32419 2372 32428
rect 2320 32385 2329 32419
rect 2329 32385 2363 32419
rect 2363 32385 2372 32419
rect 2320 32376 2372 32385
rect 1492 32308 1544 32360
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 1768 32308 1820 32360
rect 2594 32419 2646 32428
rect 2594 32385 2603 32419
rect 2603 32385 2637 32419
rect 2637 32385 2646 32419
rect 2594 32376 2646 32385
rect 3332 32419 3384 32428
rect 3332 32385 3341 32419
rect 3341 32385 3375 32419
rect 3375 32385 3384 32419
rect 3332 32376 3384 32385
rect 4528 32512 4580 32564
rect 5172 32512 5224 32564
rect 5356 32512 5408 32564
rect 6184 32512 6236 32564
rect 10140 32512 10192 32564
rect 10600 32512 10652 32564
rect 11152 32512 11204 32564
rect 6736 32444 6788 32496
rect 1860 32240 1912 32292
rect 4160 32376 4212 32428
rect 4620 32419 4672 32428
rect 4620 32385 4629 32419
rect 4629 32385 4663 32419
rect 4663 32385 4672 32419
rect 4620 32376 4672 32385
rect 4896 32376 4948 32428
rect 6092 32376 6144 32428
rect 6184 32376 6236 32428
rect 6460 32376 6512 32428
rect 8576 32444 8628 32496
rect 15016 32512 15068 32564
rect 15292 32512 15344 32564
rect 21272 32512 21324 32564
rect 8208 32376 8260 32428
rect 8392 32376 8444 32428
rect 9128 32376 9180 32428
rect 10324 32419 10376 32428
rect 10324 32385 10331 32419
rect 10331 32385 10365 32419
rect 10365 32385 10376 32419
rect 10324 32376 10376 32385
rect 10416 32376 10468 32428
rect 11980 32376 12032 32428
rect 14464 32487 14516 32496
rect 14464 32453 14473 32487
rect 14473 32453 14507 32487
rect 14507 32453 14516 32487
rect 14464 32444 14516 32453
rect 15108 32444 15160 32496
rect 14832 32419 14884 32428
rect 14832 32385 14841 32419
rect 14841 32385 14875 32419
rect 14875 32385 14884 32419
rect 14832 32376 14884 32385
rect 4068 32351 4120 32360
rect 4068 32317 4077 32351
rect 4077 32317 4111 32351
rect 4111 32317 4120 32351
rect 4068 32308 4120 32317
rect 19340 32444 19392 32496
rect 17684 32376 17736 32428
rect 19156 32419 19208 32428
rect 19156 32385 19165 32419
rect 19165 32385 19199 32419
rect 19199 32385 19208 32419
rect 19156 32376 19208 32385
rect 19708 32376 19760 32428
rect 23940 32512 23992 32564
rect 4988 32308 5040 32360
rect 5172 32308 5224 32360
rect 15108 32308 15160 32360
rect 15200 32308 15252 32360
rect 16672 32308 16724 32360
rect 16396 32240 16448 32292
rect 3056 32172 3108 32224
rect 4068 32172 4120 32224
rect 5724 32172 5776 32224
rect 9036 32215 9088 32224
rect 9036 32181 9045 32215
rect 9045 32181 9079 32215
rect 9079 32181 9088 32215
rect 9036 32172 9088 32181
rect 16580 32172 16632 32224
rect 17040 32172 17092 32224
rect 18604 32172 18656 32224
rect 20536 32215 20588 32224
rect 20536 32181 20545 32215
rect 20545 32181 20579 32215
rect 20579 32181 20588 32215
rect 20536 32172 20588 32181
rect 24124 32419 24176 32428
rect 24124 32385 24133 32419
rect 24133 32385 24167 32419
rect 24167 32385 24176 32419
rect 24124 32376 24176 32385
rect 24032 32172 24084 32224
rect 24400 32215 24452 32224
rect 24400 32181 24409 32215
rect 24409 32181 24443 32215
rect 24443 32181 24452 32215
rect 24400 32172 24452 32181
rect 3917 32070 3969 32122
rect 3981 32070 4033 32122
rect 4045 32070 4097 32122
rect 4109 32070 4161 32122
rect 4173 32070 4225 32122
rect 9851 32070 9903 32122
rect 9915 32070 9967 32122
rect 9979 32070 10031 32122
rect 10043 32070 10095 32122
rect 10107 32070 10159 32122
rect 15785 32070 15837 32122
rect 15849 32070 15901 32122
rect 15913 32070 15965 32122
rect 15977 32070 16029 32122
rect 16041 32070 16093 32122
rect 21719 32070 21771 32122
rect 21783 32070 21835 32122
rect 21847 32070 21899 32122
rect 21911 32070 21963 32122
rect 21975 32070 22027 32122
rect 1492 31968 1544 32020
rect 2596 31968 2648 32020
rect 3240 31968 3292 32020
rect 3516 31968 3568 32020
rect 5080 31968 5132 32020
rect 10508 31968 10560 32020
rect 6828 31943 6880 31952
rect 6828 31909 6837 31943
rect 6837 31909 6871 31943
rect 6871 31909 6880 31943
rect 6828 31900 6880 31909
rect 9680 31900 9732 31952
rect 10324 31900 10376 31952
rect 756 31764 808 31816
rect 1308 31764 1360 31816
rect 2136 31764 2188 31816
rect 2780 31807 2832 31816
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 3516 31832 3568 31884
rect 5816 31875 5868 31884
rect 5816 31841 5825 31875
rect 5825 31841 5859 31875
rect 5859 31841 5868 31875
rect 5816 31832 5868 31841
rect 8300 31832 8352 31884
rect 8484 31832 8536 31884
rect 13912 31968 13964 32020
rect 14004 31968 14056 32020
rect 13268 31900 13320 31952
rect 15108 32011 15160 32020
rect 15108 31977 15117 32011
rect 15117 31977 15151 32011
rect 15151 31977 15160 32011
rect 15108 31968 15160 31977
rect 15292 31968 15344 32020
rect 15752 31968 15804 32020
rect 16212 31943 16264 31952
rect 16212 31909 16221 31943
rect 16221 31909 16255 31943
rect 16255 31909 16264 31943
rect 16212 31900 16264 31909
rect 19800 31968 19852 32020
rect 20536 31968 20588 32020
rect 19340 31900 19392 31952
rect 3240 31764 3292 31816
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 4896 31807 4948 31816
rect 4896 31773 4905 31807
rect 4905 31773 4939 31807
rect 4939 31773 4948 31807
rect 4896 31764 4948 31773
rect 5540 31764 5592 31816
rect 5724 31696 5776 31748
rect 6460 31764 6512 31816
rect 12532 31764 12584 31816
rect 13820 31764 13872 31816
rect 6644 31696 6696 31748
rect 14280 31764 14332 31816
rect 15200 31764 15252 31816
rect 1768 31628 1820 31680
rect 7656 31628 7708 31680
rect 8484 31628 8536 31680
rect 9220 31628 9272 31680
rect 12072 31671 12124 31680
rect 12072 31637 12081 31671
rect 12081 31637 12115 31671
rect 12115 31637 12124 31671
rect 12072 31628 12124 31637
rect 14832 31696 14884 31748
rect 16948 31832 17000 31884
rect 17132 31832 17184 31884
rect 15476 31764 15528 31816
rect 15752 31807 15804 31816
rect 15752 31773 15761 31807
rect 15761 31773 15795 31807
rect 15795 31773 15804 31807
rect 15752 31764 15804 31773
rect 16488 31807 16540 31816
rect 16488 31773 16497 31807
rect 16497 31773 16531 31807
rect 16531 31773 16540 31807
rect 16488 31764 16540 31773
rect 20720 31900 20772 31952
rect 20904 31764 20956 31816
rect 24124 31968 24176 32020
rect 23204 31807 23256 31816
rect 23204 31773 23213 31807
rect 23213 31773 23247 31807
rect 23247 31773 23256 31807
rect 23204 31764 23256 31773
rect 25136 31764 25188 31816
rect 21548 31696 21600 31748
rect 22192 31696 22244 31748
rect 22376 31696 22428 31748
rect 15752 31628 15804 31680
rect 16028 31628 16080 31680
rect 22100 31628 22152 31680
rect 6884 31526 6936 31578
rect 6948 31526 7000 31578
rect 7012 31526 7064 31578
rect 7076 31526 7128 31578
rect 7140 31526 7192 31578
rect 12818 31526 12870 31578
rect 12882 31526 12934 31578
rect 12946 31526 12998 31578
rect 13010 31526 13062 31578
rect 13074 31526 13126 31578
rect 18752 31526 18804 31578
rect 18816 31526 18868 31578
rect 18880 31526 18932 31578
rect 18944 31526 18996 31578
rect 19008 31526 19060 31578
rect 24686 31526 24738 31578
rect 24750 31526 24802 31578
rect 24814 31526 24866 31578
rect 24878 31526 24930 31578
rect 24942 31526 24994 31578
rect 2504 31424 2556 31476
rect 3148 31424 3200 31476
rect 4160 31399 4212 31408
rect 4160 31365 4169 31399
rect 4169 31365 4203 31399
rect 4203 31365 4212 31399
rect 4160 31356 4212 31365
rect 5632 31424 5684 31476
rect 5724 31424 5776 31476
rect 4620 31356 4672 31408
rect 6000 31356 6052 31408
rect 7656 31467 7708 31476
rect 7656 31433 7665 31467
rect 7665 31433 7699 31467
rect 7699 31433 7708 31467
rect 7656 31424 7708 31433
rect 4896 31331 4948 31340
rect 4896 31297 4905 31331
rect 4905 31297 4939 31331
rect 4939 31297 4948 31331
rect 4896 31288 4948 31297
rect 5632 31288 5684 31340
rect 6184 31288 6236 31340
rect 6644 31288 6696 31340
rect 7104 31288 7156 31340
rect 9312 31356 9364 31408
rect 11152 31356 11204 31408
rect 11612 31399 11664 31408
rect 11612 31365 11621 31399
rect 11621 31365 11655 31399
rect 11655 31365 11664 31399
rect 11612 31356 11664 31365
rect 15568 31424 15620 31476
rect 17224 31424 17276 31476
rect 17960 31424 18012 31476
rect 7932 31288 7984 31340
rect 9036 31331 9088 31340
rect 9036 31297 9045 31331
rect 9045 31297 9079 31331
rect 9079 31297 9088 31331
rect 9036 31288 9088 31297
rect 9404 31331 9456 31340
rect 9404 31297 9413 31331
rect 9413 31297 9447 31331
rect 9447 31297 9456 31331
rect 9404 31288 9456 31297
rect 9772 31331 9824 31340
rect 9772 31297 9795 31331
rect 9795 31297 9824 31331
rect 9772 31288 9824 31297
rect 12440 31288 12492 31340
rect 12808 31331 12860 31340
rect 12808 31297 12815 31331
rect 12815 31297 12849 31331
rect 12849 31297 12860 31331
rect 12808 31288 12860 31297
rect 13268 31288 13320 31340
rect 1400 31263 1452 31272
rect 1400 31229 1409 31263
rect 1409 31229 1443 31263
rect 1443 31229 1452 31263
rect 1400 31220 1452 31229
rect 3332 31220 3384 31272
rect 6736 31220 6788 31272
rect 9128 31220 9180 31272
rect 1308 31084 1360 31136
rect 3700 31152 3752 31204
rect 10416 31152 10468 31204
rect 10692 31152 10744 31204
rect 2136 31084 2188 31136
rect 6092 31084 6144 31136
rect 7840 31127 7892 31136
rect 7840 31093 7849 31127
rect 7849 31093 7883 31127
rect 7883 31093 7892 31127
rect 7840 31084 7892 31093
rect 8208 31084 8260 31136
rect 8668 31084 8720 31136
rect 10324 31084 10376 31136
rect 11704 31127 11756 31136
rect 11704 31093 11713 31127
rect 11713 31093 11747 31127
rect 11747 31093 11756 31127
rect 11704 31084 11756 31093
rect 13268 31152 13320 31204
rect 13912 31331 13964 31340
rect 13912 31297 13921 31331
rect 13921 31297 13955 31331
rect 13955 31297 13964 31331
rect 13912 31288 13964 31297
rect 13728 31220 13780 31272
rect 15752 31288 15804 31340
rect 16488 31288 16540 31340
rect 17776 31288 17828 31340
rect 17960 31288 18012 31340
rect 13728 31084 13780 31136
rect 14004 31127 14056 31136
rect 14004 31093 14013 31127
rect 14013 31093 14047 31127
rect 14047 31093 14056 31127
rect 14004 31084 14056 31093
rect 19432 31288 19484 31340
rect 19340 31220 19392 31272
rect 21456 31331 21508 31340
rect 21456 31297 21465 31331
rect 21465 31297 21499 31331
rect 21499 31297 21508 31331
rect 21456 31288 21508 31297
rect 16120 31127 16172 31136
rect 16120 31093 16129 31127
rect 16129 31093 16163 31127
rect 16163 31093 16172 31127
rect 16120 31084 16172 31093
rect 17132 31084 17184 31136
rect 20628 31152 20680 31204
rect 21548 31220 21600 31272
rect 22100 31220 22152 31272
rect 21088 31195 21140 31204
rect 21088 31161 21097 31195
rect 21097 31161 21131 31195
rect 21131 31161 21140 31195
rect 21088 31152 21140 31161
rect 23296 31220 23348 31272
rect 23848 31288 23900 31340
rect 17408 31084 17460 31136
rect 18604 31127 18656 31136
rect 18604 31093 18613 31127
rect 18613 31093 18647 31127
rect 18647 31093 18656 31127
rect 18604 31084 18656 31093
rect 23940 31127 23992 31136
rect 23940 31093 23949 31127
rect 23949 31093 23983 31127
rect 23983 31093 23992 31127
rect 23940 31084 23992 31093
rect 24400 31127 24452 31136
rect 24400 31093 24409 31127
rect 24409 31093 24443 31127
rect 24443 31093 24452 31127
rect 24400 31084 24452 31093
rect 3917 30982 3969 31034
rect 3981 30982 4033 31034
rect 4045 30982 4097 31034
rect 4109 30982 4161 31034
rect 4173 30982 4225 31034
rect 9851 30982 9903 31034
rect 9915 30982 9967 31034
rect 9979 30982 10031 31034
rect 10043 30982 10095 31034
rect 10107 30982 10159 31034
rect 15785 30982 15837 31034
rect 15849 30982 15901 31034
rect 15913 30982 15965 31034
rect 15977 30982 16029 31034
rect 16041 30982 16093 31034
rect 21719 30982 21771 31034
rect 21783 30982 21835 31034
rect 21847 30982 21899 31034
rect 21911 30982 21963 31034
rect 21975 30982 22027 31034
rect 1952 30812 2004 30864
rect 3332 30923 3384 30932
rect 3332 30889 3341 30923
rect 3341 30889 3375 30923
rect 3375 30889 3384 30923
rect 3332 30880 3384 30889
rect 4620 30880 4672 30932
rect 6092 30880 6144 30932
rect 6644 30880 6696 30932
rect 7104 30880 7156 30932
rect 9036 30880 9088 30932
rect 2596 30719 2648 30728
rect 2596 30685 2603 30719
rect 2603 30685 2637 30719
rect 2637 30685 2648 30719
rect 2596 30676 2648 30685
rect 3792 30719 3844 30728
rect 3792 30685 3801 30719
rect 3801 30685 3835 30719
rect 3835 30685 3844 30719
rect 3792 30676 3844 30685
rect 4160 30676 4212 30728
rect 5816 30744 5868 30796
rect 6368 30787 6420 30796
rect 6368 30753 6377 30787
rect 6377 30753 6411 30787
rect 6411 30753 6420 30787
rect 6368 30744 6420 30753
rect 8576 30744 8628 30796
rect 4528 30719 4580 30728
rect 4528 30685 4535 30719
rect 4535 30685 4569 30719
rect 4569 30685 4580 30719
rect 4528 30676 4580 30685
rect 4620 30676 4672 30728
rect 5080 30676 5132 30728
rect 6552 30676 6604 30728
rect 9220 30719 9272 30728
rect 9220 30685 9227 30719
rect 9227 30685 9261 30719
rect 9261 30685 9272 30719
rect 9220 30676 9272 30685
rect 1492 30651 1544 30660
rect 1492 30617 1501 30651
rect 1501 30617 1535 30651
rect 1535 30617 1544 30651
rect 1492 30608 1544 30617
rect 4252 30608 4304 30660
rect 7288 30608 7340 30660
rect 8116 30608 8168 30660
rect 10968 30812 11020 30864
rect 12532 30923 12584 30932
rect 12532 30889 12541 30923
rect 12541 30889 12575 30923
rect 12575 30889 12584 30923
rect 12532 30880 12584 30889
rect 13636 30880 13688 30932
rect 14004 30880 14056 30932
rect 16120 30880 16172 30932
rect 17408 30880 17460 30932
rect 13176 30812 13228 30864
rect 11152 30787 11204 30796
rect 11152 30753 11161 30787
rect 11161 30753 11195 30787
rect 11195 30753 11204 30787
rect 11152 30744 11204 30753
rect 11244 30744 11296 30796
rect 11520 30787 11572 30796
rect 11520 30753 11554 30787
rect 11554 30753 11572 30787
rect 11520 30744 11572 30753
rect 12072 30744 12124 30796
rect 13912 30744 13964 30796
rect 14832 30812 14884 30864
rect 9772 30676 9824 30728
rect 10692 30719 10744 30728
rect 10692 30685 10701 30719
rect 10701 30685 10735 30719
rect 10735 30685 10744 30719
rect 10692 30676 10744 30685
rect 15476 30744 15528 30796
rect 572 30540 624 30592
rect 1584 30540 1636 30592
rect 4528 30540 4580 30592
rect 5264 30540 5316 30592
rect 7472 30540 7524 30592
rect 11520 30540 11572 30592
rect 12348 30540 12400 30592
rect 13820 30608 13872 30660
rect 15568 30676 15620 30728
rect 16120 30676 16172 30728
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 17960 30880 18012 30932
rect 18604 30880 18656 30932
rect 17684 30787 17736 30796
rect 17684 30753 17693 30787
rect 17693 30753 17727 30787
rect 17727 30753 17736 30787
rect 17684 30744 17736 30753
rect 20628 30880 20680 30932
rect 21456 30880 21508 30932
rect 20812 30719 20864 30728
rect 20812 30685 20821 30719
rect 20821 30685 20855 30719
rect 20855 30685 20864 30719
rect 20812 30676 20864 30685
rect 22284 30719 22336 30728
rect 22284 30685 22293 30719
rect 22293 30685 22327 30719
rect 22327 30685 22336 30719
rect 22284 30676 22336 30685
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 16396 30540 16448 30592
rect 19248 30540 19300 30592
rect 22560 30540 22612 30592
rect 25136 30608 25188 30660
rect 25688 30608 25740 30660
rect 6884 30438 6936 30490
rect 6948 30438 7000 30490
rect 7012 30438 7064 30490
rect 7076 30438 7128 30490
rect 7140 30438 7192 30490
rect 12818 30438 12870 30490
rect 12882 30438 12934 30490
rect 12946 30438 12998 30490
rect 13010 30438 13062 30490
rect 13074 30438 13126 30490
rect 18752 30438 18804 30490
rect 18816 30438 18868 30490
rect 18880 30438 18932 30490
rect 18944 30438 18996 30490
rect 19008 30438 19060 30490
rect 24686 30438 24738 30490
rect 24750 30438 24802 30490
rect 24814 30438 24866 30490
rect 24878 30438 24930 30490
rect 24942 30438 24994 30490
rect 664 30336 716 30388
rect 3700 30336 3752 30388
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 3424 30200 3476 30209
rect 4712 30268 4764 30320
rect 5908 30268 5960 30320
rect 6828 30268 6880 30320
rect 11152 30336 11204 30388
rect 13912 30336 13964 30388
rect 14372 30336 14424 30388
rect 7564 30200 7616 30252
rect 8024 30200 8076 30252
rect 10140 30200 10192 30252
rect 1676 30175 1728 30184
rect 1676 30141 1685 30175
rect 1685 30141 1719 30175
rect 1719 30141 1728 30175
rect 1676 30132 1728 30141
rect 2136 30175 2188 30184
rect 2136 30141 2145 30175
rect 2145 30141 2179 30175
rect 2179 30141 2188 30175
rect 2136 30132 2188 30141
rect 2228 30132 2280 30184
rect 2596 30132 2648 30184
rect 4160 30175 4212 30184
rect 4160 30141 4169 30175
rect 4169 30141 4203 30175
rect 4203 30141 4212 30175
rect 4160 30132 4212 30141
rect 5080 30132 5132 30184
rect 5448 30132 5500 30184
rect 5540 30132 5592 30184
rect 5908 30132 5960 30184
rect 6736 30132 6788 30184
rect 14004 30268 14056 30320
rect 14832 30268 14884 30320
rect 15016 30268 15068 30320
rect 17960 30268 18012 30320
rect 11244 30200 11296 30252
rect 1952 30064 2004 30116
rect 6000 30064 6052 30116
rect 6368 30064 6420 30116
rect 6460 30064 6512 30116
rect 5172 30039 5224 30048
rect 5172 30005 5181 30039
rect 5181 30005 5215 30039
rect 5215 30005 5224 30039
rect 5172 29996 5224 30005
rect 9036 30064 9088 30116
rect 7840 30039 7892 30048
rect 7840 30005 7849 30039
rect 7849 30005 7883 30039
rect 7883 30005 7892 30039
rect 7840 29996 7892 30005
rect 13912 30175 13964 30184
rect 13912 30141 13921 30175
rect 13921 30141 13955 30175
rect 13955 30141 13964 30175
rect 13912 30132 13964 30141
rect 16488 30200 16540 30252
rect 19248 30336 19300 30388
rect 23848 30336 23900 30388
rect 23940 30336 23992 30388
rect 19064 30200 19116 30252
rect 20536 30243 20588 30252
rect 17592 30132 17644 30184
rect 17868 30132 17920 30184
rect 12440 29996 12492 30048
rect 13820 29996 13872 30048
rect 14832 29996 14884 30048
rect 14924 30039 14976 30048
rect 14924 30005 14933 30039
rect 14933 30005 14967 30039
rect 14967 30005 14976 30039
rect 14924 29996 14976 30005
rect 17776 29996 17828 30048
rect 18236 29996 18288 30048
rect 20536 30209 20559 30243
rect 20559 30209 20588 30243
rect 20536 30200 20588 30209
rect 22100 30243 22152 30252
rect 22100 30209 22107 30243
rect 22107 30209 22141 30243
rect 22141 30209 22152 30243
rect 22100 30200 22152 30209
rect 23296 30200 23348 30252
rect 19432 30132 19484 30184
rect 19984 29996 20036 30048
rect 22284 29996 22336 30048
rect 22836 30039 22888 30048
rect 22836 30005 22845 30039
rect 22845 30005 22879 30039
rect 22879 30005 22888 30039
rect 22836 29996 22888 30005
rect 23204 30039 23256 30048
rect 23204 30005 23213 30039
rect 23213 30005 23247 30039
rect 23247 30005 23256 30039
rect 23204 29996 23256 30005
rect 24400 30039 24452 30048
rect 24400 30005 24409 30039
rect 24409 30005 24443 30039
rect 24443 30005 24452 30039
rect 24400 29996 24452 30005
rect 3917 29894 3969 29946
rect 3981 29894 4033 29946
rect 4045 29894 4097 29946
rect 4109 29894 4161 29946
rect 4173 29894 4225 29946
rect 9851 29894 9903 29946
rect 9915 29894 9967 29946
rect 9979 29894 10031 29946
rect 10043 29894 10095 29946
rect 10107 29894 10159 29946
rect 15785 29894 15837 29946
rect 15849 29894 15901 29946
rect 15913 29894 15965 29946
rect 15977 29894 16029 29946
rect 16041 29894 16093 29946
rect 21719 29894 21771 29946
rect 21783 29894 21835 29946
rect 21847 29894 21899 29946
rect 21911 29894 21963 29946
rect 21975 29894 22027 29946
rect 1124 29792 1176 29844
rect 1584 29767 1636 29776
rect 1584 29733 1593 29767
rect 1593 29733 1627 29767
rect 1627 29733 1636 29767
rect 1584 29724 1636 29733
rect 2688 29835 2740 29844
rect 2688 29801 2697 29835
rect 2697 29801 2731 29835
rect 2731 29801 2740 29835
rect 2688 29792 2740 29801
rect 2780 29792 2832 29844
rect 3056 29792 3108 29844
rect 3608 29835 3660 29844
rect 3608 29801 3617 29835
rect 3617 29801 3651 29835
rect 3651 29801 3660 29835
rect 3608 29792 3660 29801
rect 6184 29792 6236 29844
rect 7472 29792 7524 29844
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 1400 29588 1452 29597
rect 1492 29588 1544 29640
rect 1860 29588 1912 29640
rect 2412 29588 2464 29640
rect 1308 29520 1360 29572
rect 3608 29588 3660 29640
rect 7104 29724 7156 29776
rect 5172 29656 5224 29708
rect 6092 29656 6144 29708
rect 7840 29792 7892 29844
rect 8760 29835 8812 29844
rect 8760 29801 8769 29835
rect 8769 29801 8803 29835
rect 8803 29801 8812 29835
rect 8760 29792 8812 29801
rect 9036 29792 9088 29844
rect 10508 29724 10560 29776
rect 10784 29724 10836 29776
rect 11152 29767 11204 29776
rect 11152 29733 11161 29767
rect 11161 29733 11195 29767
rect 11195 29733 11204 29767
rect 11152 29724 11204 29733
rect 14648 29792 14700 29844
rect 6920 29631 6972 29640
rect 6920 29597 6929 29631
rect 6929 29597 6963 29631
rect 6963 29597 6972 29631
rect 6920 29588 6972 29597
rect 7288 29588 7340 29640
rect 10140 29656 10192 29708
rect 7932 29631 7984 29640
rect 7932 29597 7966 29631
rect 7966 29597 7984 29631
rect 7932 29588 7984 29597
rect 8116 29631 8168 29640
rect 8116 29597 8125 29631
rect 8125 29597 8159 29631
rect 8159 29597 8168 29631
rect 8116 29588 8168 29597
rect 9680 29588 9732 29640
rect 10324 29656 10376 29708
rect 11612 29656 11664 29708
rect 12072 29656 12124 29708
rect 12348 29699 12400 29708
rect 12348 29665 12357 29699
rect 12357 29665 12391 29699
rect 12391 29665 12400 29699
rect 12348 29656 12400 29665
rect 13912 29656 13964 29708
rect 15752 29699 15804 29708
rect 15752 29665 15761 29699
rect 15761 29665 15795 29699
rect 15795 29665 15804 29699
rect 15752 29656 15804 29665
rect 17500 29792 17552 29844
rect 20536 29792 20588 29844
rect 16212 29767 16264 29776
rect 16212 29733 16221 29767
rect 16221 29733 16255 29767
rect 16255 29733 16264 29767
rect 16212 29724 16264 29733
rect 17776 29724 17828 29776
rect 19892 29724 19944 29776
rect 16948 29656 17000 29708
rect 17132 29656 17184 29708
rect 10416 29588 10468 29640
rect 10600 29588 10652 29640
rect 12716 29621 12768 29640
rect 3332 29520 3384 29572
rect 4988 29495 5040 29504
rect 4988 29461 4997 29495
rect 4997 29461 5031 29495
rect 5031 29461 5040 29495
rect 4988 29452 5040 29461
rect 5264 29563 5316 29572
rect 5264 29529 5273 29563
rect 5273 29529 5307 29563
rect 5307 29529 5316 29563
rect 5264 29520 5316 29529
rect 5356 29563 5408 29572
rect 5356 29529 5365 29563
rect 5365 29529 5399 29563
rect 5399 29529 5408 29563
rect 5356 29520 5408 29529
rect 5724 29563 5776 29572
rect 5724 29529 5733 29563
rect 5733 29529 5767 29563
rect 5767 29529 5776 29563
rect 5724 29520 5776 29529
rect 6092 29495 6144 29504
rect 6092 29461 6101 29495
rect 6101 29461 6135 29495
rect 6135 29461 6144 29495
rect 6092 29452 6144 29461
rect 11980 29452 12032 29504
rect 12716 29588 12725 29621
rect 12725 29588 12768 29621
rect 14556 29588 14608 29640
rect 15936 29588 15988 29640
rect 16580 29631 16632 29640
rect 16580 29597 16614 29631
rect 16614 29597 16632 29631
rect 16580 29588 16632 29597
rect 17776 29588 17828 29640
rect 22836 29792 22888 29844
rect 23204 29792 23256 29844
rect 22560 29631 22612 29640
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 13452 29495 13504 29504
rect 13452 29461 13461 29495
rect 13461 29461 13495 29495
rect 13495 29461 13504 29495
rect 13452 29452 13504 29461
rect 14464 29452 14516 29504
rect 15936 29452 15988 29504
rect 16672 29452 16724 29504
rect 17040 29452 17092 29504
rect 17868 29452 17920 29504
rect 19984 29452 20036 29504
rect 24308 29520 24360 29572
rect 25136 29452 25188 29504
rect 6884 29350 6936 29402
rect 6948 29350 7000 29402
rect 7012 29350 7064 29402
rect 7076 29350 7128 29402
rect 7140 29350 7192 29402
rect 12818 29350 12870 29402
rect 12882 29350 12934 29402
rect 12946 29350 12998 29402
rect 13010 29350 13062 29402
rect 13074 29350 13126 29402
rect 18752 29350 18804 29402
rect 18816 29350 18868 29402
rect 18880 29350 18932 29402
rect 18944 29350 18996 29402
rect 19008 29350 19060 29402
rect 24686 29350 24738 29402
rect 24750 29350 24802 29402
rect 24814 29350 24866 29402
rect 24878 29350 24930 29402
rect 24942 29350 24994 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 940 29180 992 29232
rect 1492 29155 1544 29164
rect 1492 29121 1501 29155
rect 1501 29121 1535 29155
rect 1535 29121 1544 29155
rect 1492 29112 1544 29121
rect 3332 29180 3384 29232
rect 2504 29155 2556 29164
rect 2504 29121 2511 29155
rect 2511 29121 2545 29155
rect 2545 29121 2556 29155
rect 2504 29112 2556 29121
rect 1308 28908 1360 28960
rect 2228 29087 2280 29096
rect 2228 29053 2237 29087
rect 2237 29053 2271 29087
rect 2271 29053 2280 29087
rect 2228 29044 2280 29053
rect 1952 28976 2004 29028
rect 2044 29019 2096 29028
rect 2044 28985 2053 29019
rect 2053 28985 2087 29019
rect 2087 28985 2096 29019
rect 2044 28976 2096 28985
rect 5356 29248 5408 29300
rect 6092 29248 6144 29300
rect 7932 29180 7984 29232
rect 3608 29155 3660 29164
rect 3608 29121 3617 29155
rect 3617 29121 3651 29155
rect 3651 29121 3660 29155
rect 3608 29112 3660 29121
rect 4252 29112 4304 29164
rect 5080 29112 5132 29164
rect 7564 29112 7616 29164
rect 8116 29248 8168 29300
rect 10876 29291 10928 29300
rect 10876 29257 10885 29291
rect 10885 29257 10919 29291
rect 10919 29257 10928 29291
rect 10876 29248 10928 29257
rect 8760 29180 8812 29232
rect 11336 29248 11388 29300
rect 14004 29248 14056 29300
rect 14464 29248 14516 29300
rect 11060 29180 11112 29232
rect 11796 29180 11848 29232
rect 12164 29180 12216 29232
rect 6460 29044 6512 29096
rect 7288 29044 7340 29096
rect 2596 28908 2648 28960
rect 3240 28951 3292 28960
rect 3240 28917 3249 28951
rect 3249 28917 3283 28951
rect 3283 28917 3292 28951
rect 3240 28908 3292 28917
rect 8116 28976 8168 29028
rect 9036 29112 9088 29164
rect 9496 29155 9548 29164
rect 9496 29121 9503 29155
rect 9503 29121 9537 29155
rect 9537 29121 9548 29155
rect 9496 29112 9548 29121
rect 11336 29112 11388 29164
rect 12440 29112 12492 29164
rect 13820 29180 13872 29232
rect 14556 29223 14608 29232
rect 14556 29189 14565 29223
rect 14565 29189 14599 29223
rect 14599 29189 14608 29223
rect 14556 29180 14608 29189
rect 14832 29248 14884 29300
rect 15476 29112 15528 29164
rect 11152 28976 11204 29028
rect 11980 29044 12032 29096
rect 11796 29019 11848 29028
rect 11796 28985 11805 29019
rect 11805 28985 11839 29019
rect 11839 28985 11848 29019
rect 11796 28976 11848 28985
rect 11888 28976 11940 29028
rect 12440 28976 12492 29028
rect 14924 29044 14976 29096
rect 16856 29112 16908 29164
rect 17868 29112 17920 29164
rect 18604 29112 18656 29164
rect 9588 28908 9640 28960
rect 11428 28908 11480 28960
rect 12624 28954 12676 29006
rect 17960 28976 18012 29028
rect 18604 28976 18656 29028
rect 19616 29044 19668 29096
rect 19708 29044 19760 29096
rect 23112 28976 23164 29028
rect 13728 28908 13780 28960
rect 13820 28908 13872 28960
rect 14280 28908 14332 28960
rect 16212 28908 16264 28960
rect 17408 28908 17460 28960
rect 19616 28908 19668 28960
rect 20352 28951 20404 28960
rect 20352 28917 20361 28951
rect 20361 28917 20395 28951
rect 20395 28917 20404 28951
rect 20352 28908 20404 28917
rect 20536 28908 20588 28960
rect 21180 28908 21232 28960
rect 24400 29019 24452 29028
rect 24400 28985 24409 29019
rect 24409 28985 24443 29019
rect 24443 28985 24452 29019
rect 24400 28976 24452 28985
rect 3917 28806 3969 28858
rect 3981 28806 4033 28858
rect 4045 28806 4097 28858
rect 4109 28806 4161 28858
rect 4173 28806 4225 28858
rect 9851 28806 9903 28858
rect 9915 28806 9967 28858
rect 9979 28806 10031 28858
rect 10043 28806 10095 28858
rect 10107 28806 10159 28858
rect 15785 28806 15837 28858
rect 15849 28806 15901 28858
rect 15913 28806 15965 28858
rect 15977 28806 16029 28858
rect 16041 28806 16093 28858
rect 21719 28806 21771 28858
rect 21783 28806 21835 28858
rect 21847 28806 21899 28858
rect 21911 28806 21963 28858
rect 21975 28806 22027 28858
rect 2780 28704 2832 28756
rect 2228 28568 2280 28620
rect 9772 28704 9824 28756
rect 11152 28747 11204 28756
rect 11152 28713 11161 28747
rect 11161 28713 11195 28747
rect 11195 28713 11204 28747
rect 11152 28704 11204 28713
rect 11428 28747 11480 28756
rect 11428 28713 11437 28747
rect 11437 28713 11471 28747
rect 11471 28713 11480 28747
rect 11428 28704 11480 28713
rect 11612 28704 11664 28756
rect 13820 28704 13872 28756
rect 7288 28568 7340 28620
rect 7748 28568 7800 28620
rect 9680 28568 9732 28620
rect 19708 28704 19760 28756
rect 848 28500 900 28552
rect 2412 28432 2464 28484
rect 2964 28500 3016 28552
rect 3608 28500 3660 28552
rect 3332 28407 3384 28416
rect 3332 28373 3341 28407
rect 3341 28373 3375 28407
rect 3375 28373 3384 28407
rect 3332 28364 3384 28373
rect 3516 28364 3568 28416
rect 4896 28500 4948 28552
rect 5080 28500 5132 28552
rect 8116 28500 8168 28552
rect 8852 28500 8904 28552
rect 5356 28432 5408 28484
rect 10692 28543 10744 28552
rect 10692 28509 10701 28543
rect 10701 28509 10735 28543
rect 10735 28509 10744 28543
rect 10692 28500 10744 28509
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 11336 28543 11388 28552
rect 11336 28509 11345 28543
rect 11345 28509 11379 28543
rect 11379 28509 11388 28543
rect 11336 28500 11388 28509
rect 11612 28500 11664 28552
rect 4344 28364 4396 28416
rect 4896 28407 4948 28416
rect 4896 28373 4905 28407
rect 4905 28373 4939 28407
rect 4939 28373 4948 28407
rect 4896 28364 4948 28373
rect 5724 28364 5776 28416
rect 7472 28364 7524 28416
rect 9496 28364 9548 28416
rect 9680 28364 9732 28416
rect 10324 28364 10376 28416
rect 10876 28364 10928 28416
rect 16672 28611 16724 28620
rect 16672 28577 16681 28611
rect 16681 28577 16715 28611
rect 16715 28577 16724 28611
rect 16672 28568 16724 28577
rect 17408 28568 17460 28620
rect 19524 28636 19576 28688
rect 20352 28704 20404 28756
rect 20720 28636 20772 28688
rect 22928 28636 22980 28688
rect 12072 28432 12124 28484
rect 13912 28500 13964 28552
rect 15108 28500 15160 28552
rect 15200 28500 15252 28552
rect 15568 28500 15620 28552
rect 16120 28500 16172 28552
rect 16948 28543 17000 28552
rect 16948 28509 16957 28543
rect 16957 28509 16991 28543
rect 16991 28509 17000 28543
rect 16948 28500 17000 28509
rect 17132 28500 17184 28552
rect 17960 28500 18012 28552
rect 19156 28500 19208 28552
rect 19984 28611 20036 28620
rect 19984 28577 19993 28611
rect 19993 28577 20027 28611
rect 20027 28577 20036 28611
rect 19984 28568 20036 28577
rect 22744 28568 22796 28620
rect 19616 28543 19668 28552
rect 19616 28509 19625 28543
rect 19625 28509 19659 28543
rect 19659 28509 19668 28543
rect 19616 28500 19668 28509
rect 20352 28500 20404 28552
rect 11888 28364 11940 28416
rect 13084 28364 13136 28416
rect 13268 28364 13320 28416
rect 14004 28364 14056 28416
rect 14280 28364 14332 28416
rect 20444 28432 20496 28484
rect 23296 28500 23348 28552
rect 20996 28407 21048 28416
rect 20996 28373 21005 28407
rect 21005 28373 21039 28407
rect 21039 28373 21048 28407
rect 20996 28364 21048 28373
rect 25136 28364 25188 28416
rect 6884 28262 6936 28314
rect 6948 28262 7000 28314
rect 7012 28262 7064 28314
rect 7076 28262 7128 28314
rect 7140 28262 7192 28314
rect 12818 28262 12870 28314
rect 12882 28262 12934 28314
rect 12946 28262 12998 28314
rect 13010 28262 13062 28314
rect 13074 28262 13126 28314
rect 18752 28262 18804 28314
rect 18816 28262 18868 28314
rect 18880 28262 18932 28314
rect 18944 28262 18996 28314
rect 19008 28262 19060 28314
rect 24686 28262 24738 28314
rect 24750 28262 24802 28314
rect 24814 28262 24866 28314
rect 24878 28262 24930 28314
rect 24942 28262 24994 28314
rect 2964 28160 3016 28212
rect 3332 28160 3384 28212
rect 3792 28160 3844 28212
rect 3884 28203 3936 28212
rect 3884 28169 3893 28203
rect 3893 28169 3927 28203
rect 3927 28169 3936 28203
rect 3884 28160 3936 28169
rect 940 28092 992 28144
rect 756 28024 808 28076
rect 2044 28092 2096 28144
rect 2780 28135 2832 28144
rect 2780 28101 2789 28135
rect 2789 28101 2823 28135
rect 2823 28101 2832 28135
rect 2780 28092 2832 28101
rect 2320 28067 2372 28076
rect 2320 28033 2329 28067
rect 2329 28033 2363 28067
rect 2363 28033 2372 28067
rect 2320 28024 2372 28033
rect 4344 28092 4396 28144
rect 4528 28135 4580 28144
rect 4528 28101 4537 28135
rect 4537 28101 4571 28135
rect 4571 28101 4580 28135
rect 4528 28092 4580 28101
rect 4804 28135 4856 28144
rect 4804 28101 4813 28135
rect 4813 28101 4847 28135
rect 4847 28101 4856 28135
rect 4804 28092 4856 28101
rect 5540 28092 5592 28144
rect 9128 28160 9180 28212
rect 3516 28067 3568 28076
rect 3516 28033 3525 28067
rect 3525 28033 3559 28067
rect 3559 28033 3568 28067
rect 3516 28024 3568 28033
rect 5356 28024 5408 28076
rect 7564 28024 7616 28076
rect 8116 28024 8168 28076
rect 9956 28024 10008 28076
rect 3240 27956 3292 28008
rect 4896 27956 4948 28008
rect 6092 27956 6144 28008
rect 6368 27999 6420 28008
rect 6368 27965 6377 27999
rect 6377 27965 6411 27999
rect 6411 27965 6420 27999
rect 6368 27956 6420 27965
rect 11336 28024 11388 28076
rect 11612 28024 11664 28076
rect 11796 28024 11848 28076
rect 12072 27956 12124 28008
rect 12624 27956 12676 28008
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 1860 27888 1912 27940
rect 2688 27888 2740 27940
rect 12164 27888 12216 27940
rect 13820 27999 13872 28008
rect 13820 27965 13854 27999
rect 13854 27965 13872 27999
rect 13820 27956 13872 27965
rect 2780 27820 2832 27872
rect 6736 27820 6788 27872
rect 11060 27863 11112 27872
rect 11060 27829 11069 27863
rect 11069 27829 11103 27863
rect 11103 27829 11112 27863
rect 11060 27820 11112 27829
rect 13728 27820 13780 27872
rect 14648 27863 14700 27872
rect 14648 27829 14657 27863
rect 14657 27829 14691 27863
rect 14691 27829 14700 27863
rect 14648 27820 14700 27829
rect 16672 28160 16724 28212
rect 19156 28160 19208 28212
rect 19524 28160 19576 28212
rect 20720 28160 20772 28212
rect 20996 28160 21048 28212
rect 21456 28160 21508 28212
rect 14924 28024 14976 28076
rect 15108 27956 15160 28008
rect 17684 27956 17736 28008
rect 17960 28024 18012 28076
rect 19432 28067 19484 28076
rect 19432 28033 19441 28067
rect 19441 28033 19475 28067
rect 19475 28033 19484 28067
rect 19432 28024 19484 28033
rect 19708 28067 19760 28076
rect 19708 28033 19731 28067
rect 19731 28033 19760 28067
rect 19708 28024 19760 28033
rect 22744 28160 22796 28212
rect 16672 27888 16724 27940
rect 17316 27888 17368 27940
rect 20628 27956 20680 28008
rect 21548 27888 21600 27940
rect 22836 28067 22888 28076
rect 22836 28033 22845 28067
rect 22845 28033 22879 28067
rect 22879 28033 22888 28067
rect 22836 28024 22888 28033
rect 22928 28024 22980 28076
rect 23940 28067 23992 28076
rect 23940 28033 23949 28067
rect 23949 28033 23983 28067
rect 23983 28033 23992 28067
rect 23940 28024 23992 28033
rect 20812 27863 20864 27872
rect 20812 27829 20821 27863
rect 20821 27829 20855 27863
rect 20855 27829 20864 27863
rect 20812 27820 20864 27829
rect 22560 27820 22612 27872
rect 23480 27820 23532 27872
rect 23756 27863 23808 27872
rect 23756 27829 23765 27863
rect 23765 27829 23799 27863
rect 23799 27829 23808 27863
rect 23756 27820 23808 27829
rect 24400 27863 24452 27872
rect 24400 27829 24409 27863
rect 24409 27829 24443 27863
rect 24443 27829 24452 27863
rect 24400 27820 24452 27829
rect 3917 27718 3969 27770
rect 3981 27718 4033 27770
rect 4045 27718 4097 27770
rect 4109 27718 4161 27770
rect 4173 27718 4225 27770
rect 9851 27718 9903 27770
rect 9915 27718 9967 27770
rect 9979 27718 10031 27770
rect 10043 27718 10095 27770
rect 10107 27718 10159 27770
rect 15785 27718 15837 27770
rect 15849 27718 15901 27770
rect 15913 27718 15965 27770
rect 15977 27718 16029 27770
rect 16041 27718 16093 27770
rect 21719 27718 21771 27770
rect 21783 27718 21835 27770
rect 21847 27718 21899 27770
rect 21911 27718 21963 27770
rect 21975 27718 22027 27770
rect 1768 27616 1820 27668
rect 3792 27616 3844 27668
rect 5264 27616 5316 27668
rect 9128 27616 9180 27668
rect 7932 27480 7984 27532
rect 20 27412 72 27464
rect 1860 27344 1912 27396
rect 1124 27276 1176 27328
rect 2688 27344 2740 27396
rect 4988 27412 5040 27464
rect 6092 27412 6144 27464
rect 6736 27455 6788 27464
rect 6736 27421 6745 27455
rect 6745 27421 6779 27455
rect 6779 27421 6788 27455
rect 6736 27412 6788 27421
rect 2504 27276 2556 27328
rect 6552 27344 6604 27396
rect 6644 27387 6696 27396
rect 6644 27353 6653 27387
rect 6653 27353 6687 27387
rect 6687 27353 6696 27387
rect 6644 27344 6696 27353
rect 3792 27276 3844 27328
rect 4528 27276 4580 27328
rect 6460 27276 6512 27328
rect 7288 27276 7340 27328
rect 7656 27319 7708 27328
rect 7656 27285 7665 27319
rect 7665 27285 7699 27319
rect 7699 27285 7708 27319
rect 7656 27276 7708 27285
rect 8208 27276 8260 27328
rect 9220 27480 9272 27532
rect 9588 27523 9640 27532
rect 9588 27489 9597 27523
rect 9597 27489 9631 27523
rect 9631 27489 9640 27523
rect 9588 27480 9640 27489
rect 10048 27480 10100 27532
rect 10324 27480 10376 27532
rect 12808 27480 12860 27532
rect 9864 27455 9916 27464
rect 9864 27421 9873 27455
rect 9873 27421 9907 27455
rect 9907 27421 9916 27455
rect 9864 27412 9916 27421
rect 11520 27455 11572 27464
rect 11520 27421 11529 27455
rect 11529 27421 11563 27455
rect 11563 27421 11572 27455
rect 11520 27412 11572 27421
rect 10784 27387 10836 27396
rect 10784 27353 10793 27387
rect 10793 27353 10827 27387
rect 10827 27353 10836 27387
rect 10784 27344 10836 27353
rect 11428 27344 11480 27396
rect 12256 27412 12308 27464
rect 13820 27344 13872 27396
rect 12440 27276 12492 27328
rect 15108 27480 15160 27532
rect 16212 27523 16264 27532
rect 16212 27489 16221 27523
rect 16221 27489 16255 27523
rect 16255 27489 16264 27523
rect 16212 27480 16264 27489
rect 17316 27480 17368 27532
rect 14648 27412 14700 27464
rect 17224 27412 17276 27464
rect 20628 27616 20680 27668
rect 21456 27616 21508 27668
rect 22836 27616 22888 27668
rect 23940 27616 23992 27668
rect 19432 27480 19484 27532
rect 14648 27276 14700 27328
rect 15016 27319 15068 27328
rect 15016 27285 15025 27319
rect 15025 27285 15059 27319
rect 15059 27285 15068 27319
rect 15016 27276 15068 27285
rect 16488 27276 16540 27328
rect 19708 27412 19760 27464
rect 20812 27412 20864 27464
rect 21180 27455 21232 27464
rect 21180 27421 21189 27455
rect 21189 27421 21223 27455
rect 21223 27421 21232 27455
rect 21180 27412 21232 27421
rect 21548 27344 21600 27396
rect 22744 27412 22796 27464
rect 22836 27344 22888 27396
rect 23480 27455 23532 27464
rect 23480 27421 23489 27455
rect 23489 27421 23523 27455
rect 23523 27421 23532 27455
rect 23480 27412 23532 27421
rect 23572 27412 23624 27464
rect 17224 27319 17276 27328
rect 17224 27285 17233 27319
rect 17233 27285 17267 27319
rect 17267 27285 17276 27319
rect 17224 27276 17276 27285
rect 17868 27276 17920 27328
rect 22744 27276 22796 27328
rect 23020 27276 23072 27328
rect 25136 27276 25188 27328
rect 6884 27174 6936 27226
rect 6948 27174 7000 27226
rect 7012 27174 7064 27226
rect 7076 27174 7128 27226
rect 7140 27174 7192 27226
rect 12818 27174 12870 27226
rect 12882 27174 12934 27226
rect 12946 27174 12998 27226
rect 13010 27174 13062 27226
rect 13074 27174 13126 27226
rect 18752 27174 18804 27226
rect 18816 27174 18868 27226
rect 18880 27174 18932 27226
rect 18944 27174 18996 27226
rect 19008 27174 19060 27226
rect 24686 27174 24738 27226
rect 24750 27174 24802 27226
rect 24814 27174 24866 27226
rect 24878 27174 24930 27226
rect 24942 27174 24994 27226
rect 1216 27072 1268 27124
rect 2044 27047 2096 27056
rect 2044 27013 2053 27047
rect 2053 27013 2087 27047
rect 2087 27013 2096 27047
rect 2044 27004 2096 27013
rect 1308 26936 1360 26988
rect 2688 27004 2740 27056
rect 3056 27004 3108 27056
rect 3148 27047 3200 27056
rect 3148 27013 3157 27047
rect 3157 27013 3191 27047
rect 3191 27013 3200 27047
rect 3148 27004 3200 27013
rect 2320 26979 2372 26988
rect 2320 26945 2329 26979
rect 2329 26945 2363 26979
rect 2363 26945 2372 26979
rect 2320 26936 2372 26945
rect 2412 26979 2464 26988
rect 2412 26945 2421 26979
rect 2421 26945 2455 26979
rect 2455 26945 2464 26979
rect 2412 26936 2464 26945
rect 2964 26936 3016 26988
rect 2504 26868 2556 26920
rect 3332 26936 3384 26988
rect 6552 27072 6604 27124
rect 5356 27004 5408 27056
rect 9588 27072 9640 27124
rect 11520 27072 11572 27124
rect 12716 27072 12768 27124
rect 15200 27072 15252 27124
rect 3608 26936 3660 26988
rect 4528 26979 4580 26988
rect 4528 26945 4537 26979
rect 4537 26945 4571 26979
rect 4571 26945 4580 26979
rect 4528 26936 4580 26945
rect 4896 26936 4948 26988
rect 7748 26979 7800 26988
rect 7748 26945 7757 26979
rect 7757 26945 7791 26979
rect 7791 26945 7800 26979
rect 7748 26936 7800 26945
rect 8116 26936 8168 26988
rect 5540 26868 5592 26920
rect 20720 27072 20772 27124
rect 20812 27072 20864 27124
rect 18604 27004 18656 27056
rect 19616 27004 19668 27056
rect 22836 27115 22888 27124
rect 22836 27081 22845 27115
rect 22845 27081 22879 27115
rect 22879 27081 22888 27115
rect 22836 27072 22888 27081
rect 23020 27072 23072 27124
rect 23572 27072 23624 27124
rect 23756 27072 23808 27124
rect 10416 26936 10468 26988
rect 11612 26936 11664 26988
rect 12716 26936 12768 26988
rect 13820 26979 13872 26988
rect 13820 26945 13854 26979
rect 13854 26945 13872 26979
rect 13820 26936 13872 26945
rect 15108 26936 15160 26988
rect 12624 26868 12676 26920
rect 12900 26868 12952 26920
rect 13452 26911 13504 26920
rect 13452 26877 13461 26911
rect 13461 26877 13495 26911
rect 13495 26877 13504 26911
rect 13452 26868 13504 26877
rect 5356 26732 5408 26784
rect 5816 26800 5868 26852
rect 9312 26800 9364 26852
rect 13268 26800 13320 26852
rect 9772 26732 9824 26784
rect 11244 26732 11296 26784
rect 14648 26868 14700 26920
rect 16764 26936 16816 26988
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 22192 26936 22244 26988
rect 23756 26979 23808 26988
rect 23756 26945 23765 26979
rect 23765 26945 23799 26979
rect 23799 26945 23808 26979
rect 23756 26936 23808 26945
rect 16856 26911 16908 26920
rect 16856 26877 16865 26911
rect 16865 26877 16899 26911
rect 16899 26877 16908 26911
rect 16856 26868 16908 26877
rect 17224 26868 17276 26920
rect 17592 26911 17644 26920
rect 17592 26877 17601 26911
rect 17601 26877 17635 26911
rect 17635 26877 17644 26911
rect 17592 26868 17644 26877
rect 17776 26868 17828 26920
rect 19984 26868 20036 26920
rect 21548 26868 21600 26920
rect 17408 26732 17460 26784
rect 19432 26732 19484 26784
rect 22744 26732 22796 26784
rect 23940 26732 23992 26784
rect 24400 26775 24452 26784
rect 24400 26741 24409 26775
rect 24409 26741 24443 26775
rect 24443 26741 24452 26775
rect 24400 26732 24452 26741
rect 3917 26630 3969 26682
rect 3981 26630 4033 26682
rect 4045 26630 4097 26682
rect 4109 26630 4161 26682
rect 4173 26630 4225 26682
rect 9851 26630 9903 26682
rect 9915 26630 9967 26682
rect 9979 26630 10031 26682
rect 10043 26630 10095 26682
rect 10107 26630 10159 26682
rect 15785 26630 15837 26682
rect 15849 26630 15901 26682
rect 15913 26630 15965 26682
rect 15977 26630 16029 26682
rect 16041 26630 16093 26682
rect 21719 26630 21771 26682
rect 21783 26630 21835 26682
rect 21847 26630 21899 26682
rect 21911 26630 21963 26682
rect 21975 26630 22027 26682
rect 2412 26528 2464 26580
rect 3240 26571 3292 26580
rect 3240 26537 3249 26571
rect 3249 26537 3283 26571
rect 3283 26537 3292 26571
rect 3240 26528 3292 26537
rect 3516 26528 3568 26580
rect 2964 26460 3016 26512
rect 3608 26460 3660 26512
rect 4528 26460 4580 26512
rect 9680 26460 9732 26512
rect 10968 26528 11020 26580
rect 12900 26528 12952 26580
rect 13636 26528 13688 26580
rect 11152 26460 11204 26512
rect 15844 26528 15896 26580
rect 16028 26528 16080 26580
rect 20260 26528 20312 26580
rect 20444 26528 20496 26580
rect 23756 26528 23808 26580
rect 2320 26392 2372 26444
rect 4344 26392 4396 26444
rect 6092 26392 6144 26444
rect 6552 26435 6604 26444
rect 6552 26401 6561 26435
rect 6561 26401 6595 26435
rect 6595 26401 6604 26435
rect 6552 26392 6604 26401
rect 9956 26392 10008 26444
rect 10324 26392 10376 26444
rect 10784 26392 10836 26444
rect 1492 26324 1544 26376
rect 1768 26324 1820 26376
rect 2964 26324 3016 26376
rect 3240 26324 3292 26376
rect 3516 26367 3568 26376
rect 3516 26333 3525 26367
rect 3525 26333 3559 26367
rect 3559 26333 3568 26367
rect 3516 26324 3568 26333
rect 4068 26367 4120 26376
rect 4068 26333 4077 26367
rect 4077 26333 4111 26367
rect 4111 26333 4120 26367
rect 4068 26324 4120 26333
rect 4896 26324 4948 26376
rect 5540 26324 5592 26376
rect 6828 26367 6880 26376
rect 6828 26333 6835 26367
rect 6835 26333 6869 26367
rect 6869 26333 6880 26367
rect 6828 26324 6880 26333
rect 7840 26324 7892 26376
rect 9312 26324 9364 26376
rect 10140 26367 10192 26376
rect 10140 26333 10149 26367
rect 10149 26333 10183 26367
rect 10183 26333 10192 26367
rect 10140 26324 10192 26333
rect 10416 26367 10468 26376
rect 10416 26333 10425 26367
rect 10425 26333 10459 26367
rect 10459 26333 10468 26367
rect 10416 26324 10468 26333
rect 11060 26392 11112 26444
rect 19524 26460 19576 26512
rect 25320 26664 25372 26716
rect 15936 26392 15988 26444
rect 18696 26392 18748 26444
rect 25228 26460 25280 26512
rect 13912 26324 13964 26376
rect 14740 26324 14792 26376
rect 572 26188 624 26240
rect 2044 26188 2096 26240
rect 2596 26188 2648 26240
rect 9128 26256 9180 26308
rect 11244 26256 11296 26308
rect 11888 26299 11940 26308
rect 11888 26265 11897 26299
rect 11897 26265 11931 26299
rect 11931 26265 11940 26299
rect 11888 26256 11940 26265
rect 12256 26299 12308 26308
rect 12256 26265 12265 26299
rect 12265 26265 12299 26299
rect 12299 26265 12308 26299
rect 12256 26256 12308 26265
rect 12348 26256 12400 26308
rect 15660 26324 15712 26376
rect 4988 26188 5040 26240
rect 6184 26188 6236 26240
rect 7564 26231 7616 26240
rect 7564 26197 7573 26231
rect 7573 26197 7607 26231
rect 7607 26197 7616 26231
rect 7564 26188 7616 26197
rect 7840 26188 7892 26240
rect 12624 26231 12676 26240
rect 12624 26197 12633 26231
rect 12633 26197 12667 26231
rect 12667 26197 12676 26231
rect 12624 26188 12676 26197
rect 15844 26256 15896 26308
rect 16028 26256 16080 26308
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 23572 26324 23624 26376
rect 25136 26256 25188 26308
rect 16856 26188 16908 26240
rect 17960 26188 18012 26240
rect 19248 26231 19300 26240
rect 19248 26197 19257 26231
rect 19257 26197 19291 26231
rect 19291 26197 19300 26231
rect 19248 26188 19300 26197
rect 23664 26231 23716 26240
rect 23664 26197 23673 26231
rect 23673 26197 23707 26231
rect 23707 26197 23716 26231
rect 23664 26188 23716 26197
rect 6884 26086 6936 26138
rect 6948 26086 7000 26138
rect 7012 26086 7064 26138
rect 7076 26086 7128 26138
rect 7140 26086 7192 26138
rect 12818 26086 12870 26138
rect 12882 26086 12934 26138
rect 12946 26086 12998 26138
rect 13010 26086 13062 26138
rect 13074 26086 13126 26138
rect 18752 26086 18804 26138
rect 18816 26086 18868 26138
rect 18880 26086 18932 26138
rect 18944 26086 18996 26138
rect 19008 26086 19060 26138
rect 24686 26086 24738 26138
rect 24750 26086 24802 26138
rect 24814 26086 24866 26138
rect 24878 26086 24930 26138
rect 24942 26086 24994 26138
rect 1676 25984 1728 26036
rect 2596 25984 2648 26036
rect 1308 25916 1360 25968
rect 7840 25984 7892 26036
rect 1032 25848 1084 25900
rect 1492 25891 1544 25900
rect 1492 25857 1501 25891
rect 1501 25857 1535 25891
rect 1535 25857 1544 25891
rect 1492 25848 1544 25857
rect 1768 25891 1820 25900
rect 1768 25857 1775 25891
rect 1775 25857 1809 25891
rect 1809 25857 1820 25891
rect 1768 25848 1820 25857
rect 1860 25848 1912 25900
rect 2688 25848 2740 25900
rect 3976 25916 4028 25968
rect 2228 25712 2280 25764
rect 3332 25848 3384 25900
rect 4436 25848 4488 25900
rect 5356 25916 5408 25968
rect 6000 25916 6052 25968
rect 7104 25959 7156 25968
rect 7104 25925 7113 25959
rect 7113 25925 7147 25959
rect 7147 25925 7156 25959
rect 7104 25916 7156 25925
rect 7288 25916 7340 25968
rect 7656 25848 7708 25900
rect 10692 25984 10744 26036
rect 11152 25984 11204 26036
rect 12256 25984 12308 26036
rect 12532 25984 12584 26036
rect 13452 25984 13504 26036
rect 15016 25984 15068 26036
rect 15660 26027 15712 26036
rect 15660 25993 15669 26027
rect 15669 25993 15703 26027
rect 15703 25993 15712 26027
rect 15660 25984 15712 25993
rect 15936 25984 15988 26036
rect 16028 26027 16080 26036
rect 16028 25993 16037 26027
rect 16037 25993 16071 26027
rect 16071 25993 16080 26027
rect 16028 25984 16080 25993
rect 16488 25984 16540 26036
rect 17224 25984 17276 26036
rect 8208 25848 8260 25900
rect 10048 25891 10100 25900
rect 10048 25857 10082 25891
rect 10082 25857 10100 25891
rect 10048 25848 10100 25857
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 11888 25916 11940 25968
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 14280 25891 14332 25900
rect 14280 25857 14289 25891
rect 14289 25857 14323 25891
rect 14323 25857 14332 25891
rect 14280 25848 14332 25857
rect 19984 25984 20036 26036
rect 18696 25916 18748 25968
rect 23572 25984 23624 26036
rect 24032 25984 24084 26036
rect 7564 25780 7616 25832
rect 8300 25780 8352 25832
rect 9220 25823 9272 25832
rect 9220 25789 9229 25823
rect 9229 25789 9263 25823
rect 9263 25789 9272 25823
rect 9220 25780 9272 25789
rect 10416 25780 10468 25832
rect 12348 25780 12400 25832
rect 9588 25712 9640 25764
rect 9680 25755 9732 25764
rect 9680 25721 9689 25755
rect 9689 25721 9723 25755
rect 9723 25721 9732 25755
rect 9680 25712 9732 25721
rect 13728 25823 13780 25832
rect 13728 25789 13737 25823
rect 13737 25789 13771 25823
rect 13771 25789 13780 25823
rect 13728 25780 13780 25789
rect 14004 25823 14056 25832
rect 14004 25789 14013 25823
rect 14013 25789 14047 25823
rect 14047 25789 14056 25823
rect 14004 25780 14056 25789
rect 14096 25823 14148 25832
rect 14096 25789 14130 25823
rect 14130 25789 14148 25823
rect 14096 25780 14148 25789
rect 20628 25848 20680 25900
rect 21364 25891 21416 25900
rect 21364 25857 21373 25891
rect 21373 25857 21407 25891
rect 21407 25857 21416 25891
rect 21364 25848 21416 25857
rect 21548 25891 21600 25900
rect 21548 25857 21557 25891
rect 21557 25857 21591 25891
rect 21591 25857 21600 25891
rect 21548 25848 21600 25857
rect 24124 25959 24176 25968
rect 24124 25925 24133 25959
rect 24133 25925 24167 25959
rect 24167 25925 24176 25959
rect 24124 25916 24176 25925
rect 23572 25848 23624 25900
rect 22100 25780 22152 25832
rect 23388 25780 23440 25832
rect 23940 25712 23992 25764
rect 1952 25644 2004 25696
rect 2596 25644 2648 25696
rect 3056 25644 3108 25696
rect 3332 25644 3384 25696
rect 4252 25644 4304 25696
rect 4436 25687 4488 25696
rect 4436 25653 4445 25687
rect 4445 25653 4479 25687
rect 4479 25653 4488 25687
rect 4436 25644 4488 25653
rect 4896 25644 4948 25696
rect 5816 25687 5868 25696
rect 5816 25653 5825 25687
rect 5825 25653 5859 25687
rect 5859 25653 5868 25687
rect 5816 25644 5868 25653
rect 6092 25644 6144 25696
rect 7104 25644 7156 25696
rect 12348 25644 12400 25696
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 13268 25644 13320 25696
rect 20076 25687 20128 25696
rect 20076 25653 20085 25687
rect 20085 25653 20119 25687
rect 20119 25653 20128 25687
rect 20076 25644 20128 25653
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 23112 25687 23164 25696
rect 23112 25653 23121 25687
rect 23121 25653 23155 25687
rect 23155 25653 23164 25687
rect 23112 25644 23164 25653
rect 24400 25687 24452 25696
rect 24400 25653 24409 25687
rect 24409 25653 24443 25687
rect 24443 25653 24452 25687
rect 24400 25644 24452 25653
rect 3917 25542 3969 25594
rect 3981 25542 4033 25594
rect 4045 25542 4097 25594
rect 4109 25542 4161 25594
rect 4173 25542 4225 25594
rect 9851 25542 9903 25594
rect 9915 25542 9967 25594
rect 9979 25542 10031 25594
rect 10043 25542 10095 25594
rect 10107 25542 10159 25594
rect 15785 25542 15837 25594
rect 15849 25542 15901 25594
rect 15913 25542 15965 25594
rect 15977 25542 16029 25594
rect 16041 25542 16093 25594
rect 21719 25542 21771 25594
rect 21783 25542 21835 25594
rect 21847 25542 21899 25594
rect 21911 25542 21963 25594
rect 21975 25542 22027 25594
rect 1216 25440 1268 25492
rect 2228 25440 2280 25492
rect 2136 25372 2188 25424
rect 3240 25440 3292 25492
rect 5448 25440 5500 25492
rect 7748 25440 7800 25492
rect 8484 25440 8536 25492
rect 8852 25440 8904 25492
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 2136 25279 2188 25288
rect 2136 25245 2145 25279
rect 2145 25245 2179 25279
rect 2179 25245 2188 25279
rect 2136 25236 2188 25245
rect 2688 25236 2740 25288
rect 4068 25236 4120 25288
rect 4436 25236 4488 25288
rect 4528 25236 4580 25288
rect 6552 25304 6604 25356
rect 7288 25347 7340 25356
rect 7288 25313 7297 25347
rect 7297 25313 7331 25347
rect 7331 25313 7340 25347
rect 7288 25304 7340 25313
rect 8852 25304 8904 25356
rect 9404 25304 9456 25356
rect 10416 25440 10468 25492
rect 18236 25440 18288 25492
rect 20076 25440 20128 25492
rect 19524 25372 19576 25424
rect 20628 25440 20680 25492
rect 21364 25483 21416 25492
rect 21364 25449 21373 25483
rect 21373 25449 21407 25483
rect 21407 25449 21416 25483
rect 21364 25440 21416 25449
rect 23112 25440 23164 25492
rect 23572 25440 23624 25492
rect 23664 25440 23716 25492
rect 1860 25143 1912 25152
rect 1860 25109 1869 25143
rect 1869 25109 1903 25143
rect 1903 25109 1912 25143
rect 1860 25100 1912 25109
rect 4620 25168 4672 25220
rect 5448 25279 5500 25288
rect 5448 25245 5457 25279
rect 5457 25245 5491 25279
rect 5491 25245 5500 25279
rect 5448 25236 5500 25245
rect 6920 25236 6972 25288
rect 7564 25279 7616 25288
rect 7564 25245 7571 25279
rect 7571 25245 7605 25279
rect 7605 25245 7616 25279
rect 7564 25236 7616 25245
rect 10876 25236 10928 25288
rect 3516 25100 3568 25152
rect 3792 25100 3844 25152
rect 3976 25143 4028 25152
rect 3976 25109 3985 25143
rect 3985 25109 4019 25143
rect 4019 25109 4028 25143
rect 3976 25100 4028 25109
rect 4160 25100 4212 25152
rect 8668 25168 8720 25220
rect 9036 25168 9088 25220
rect 9588 25168 9640 25220
rect 10140 25168 10192 25220
rect 12532 25304 12584 25356
rect 15384 25304 15436 25356
rect 16764 25304 16816 25356
rect 17316 25347 17368 25356
rect 17316 25313 17325 25347
rect 17325 25313 17359 25347
rect 17359 25313 17368 25347
rect 17316 25304 17368 25313
rect 17408 25304 17460 25356
rect 18512 25304 18564 25356
rect 11704 25211 11756 25220
rect 11704 25177 11713 25211
rect 11713 25177 11747 25211
rect 11747 25177 11756 25211
rect 11704 25168 11756 25177
rect 12348 25236 12400 25288
rect 6092 25100 6144 25152
rect 6368 25100 6420 25152
rect 8116 25100 8168 25152
rect 11520 25100 11572 25152
rect 12072 25100 12124 25152
rect 12440 25168 12492 25220
rect 12256 25100 12308 25152
rect 12348 25100 12400 25152
rect 12624 25168 12676 25220
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 19708 25304 19760 25356
rect 19984 25304 20036 25356
rect 21180 25304 21232 25356
rect 23480 25304 23532 25356
rect 20628 25279 20680 25288
rect 20628 25245 20635 25279
rect 20635 25245 20669 25279
rect 20669 25245 20680 25279
rect 20628 25236 20680 25245
rect 22560 25236 22612 25288
rect 16672 25168 16724 25220
rect 22100 25211 22152 25220
rect 22100 25177 22134 25211
rect 22134 25177 22152 25211
rect 22100 25168 22152 25177
rect 25136 25168 25188 25220
rect 19248 25100 19300 25152
rect 21180 25100 21232 25152
rect 23756 25100 23808 25152
rect 6884 24998 6936 25050
rect 6948 24998 7000 25050
rect 7012 24998 7064 25050
rect 7076 24998 7128 25050
rect 7140 24998 7192 25050
rect 12818 24998 12870 25050
rect 12882 24998 12934 25050
rect 12946 24998 12998 25050
rect 13010 24998 13062 25050
rect 13074 24998 13126 25050
rect 18752 24998 18804 25050
rect 18816 24998 18868 25050
rect 18880 24998 18932 25050
rect 18944 24998 18996 25050
rect 19008 24998 19060 25050
rect 24686 24998 24738 25050
rect 24750 24998 24802 25050
rect 24814 24998 24866 25050
rect 24878 24998 24930 25050
rect 24942 24998 24994 25050
rect 1308 24828 1360 24880
rect 2044 24896 2096 24948
rect 2964 24896 3016 24948
rect 3056 24896 3108 24948
rect 756 24760 808 24812
rect 1492 24760 1544 24812
rect 1124 24692 1176 24744
rect 2780 24760 2832 24812
rect 3240 24803 3292 24812
rect 3240 24769 3249 24803
rect 3249 24769 3283 24803
rect 3283 24769 3292 24803
rect 3240 24760 3292 24769
rect 3516 24828 3568 24880
rect 4160 24896 4212 24948
rect 8208 24896 8260 24948
rect 8300 24896 8352 24948
rect 12256 24896 12308 24948
rect 15016 24896 15068 24948
rect 3792 24760 3844 24812
rect 3976 24760 4028 24812
rect 4528 24803 4580 24812
rect 4528 24769 4537 24803
rect 4537 24769 4571 24803
rect 4571 24769 4580 24803
rect 4528 24760 4580 24769
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 6460 24760 6512 24812
rect 8024 24760 8076 24812
rect 8852 24828 8904 24880
rect 9220 24828 9272 24880
rect 12164 24828 12216 24880
rect 8668 24760 8720 24812
rect 11336 24760 11388 24812
rect 11520 24760 11572 24812
rect 12716 24828 12768 24880
rect 3516 24692 3568 24744
rect 4068 24692 4120 24744
rect 4436 24692 4488 24744
rect 2596 24624 2648 24676
rect 4160 24667 4212 24676
rect 4160 24633 4169 24667
rect 4169 24633 4203 24667
rect 4203 24633 4212 24667
rect 4160 24624 4212 24633
rect 4252 24624 4304 24676
rect 6368 24692 6420 24744
rect 11796 24692 11848 24744
rect 12072 24692 12124 24744
rect 16764 24828 16816 24880
rect 17316 24896 17368 24948
rect 21364 24896 21416 24948
rect 21548 24896 21600 24948
rect 23480 24939 23532 24948
rect 23480 24905 23489 24939
rect 23489 24905 23523 24939
rect 23523 24905 23532 24939
rect 23480 24896 23532 24905
rect 16580 24760 16632 24812
rect 18604 24828 18656 24880
rect 19248 24828 19300 24880
rect 17868 24760 17920 24812
rect 18236 24760 18288 24812
rect 18696 24760 18748 24812
rect 19984 24760 20036 24812
rect 21640 24828 21692 24880
rect 21456 24692 21508 24744
rect 2412 24599 2464 24608
rect 2412 24565 2421 24599
rect 2421 24565 2455 24599
rect 2455 24565 2464 24599
rect 2412 24556 2464 24565
rect 8300 24624 8352 24676
rect 9680 24624 9732 24676
rect 10140 24624 10192 24676
rect 10968 24624 11020 24676
rect 11704 24624 11756 24676
rect 5724 24556 5776 24608
rect 5908 24556 5960 24608
rect 6184 24599 6236 24608
rect 6184 24565 6193 24599
rect 6193 24565 6227 24599
rect 6227 24565 6236 24599
rect 6184 24556 6236 24565
rect 8760 24556 8812 24608
rect 13176 24599 13228 24608
rect 13176 24565 13185 24599
rect 13185 24565 13219 24599
rect 13219 24565 13228 24599
rect 13176 24556 13228 24565
rect 22376 24760 22428 24812
rect 24308 24760 24360 24812
rect 22100 24692 22152 24744
rect 17776 24556 17828 24608
rect 18512 24556 18564 24608
rect 19892 24556 19944 24608
rect 20628 24556 20680 24608
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 21548 24599 21600 24608
rect 21548 24565 21557 24599
rect 21557 24565 21591 24599
rect 21591 24565 21600 24599
rect 21548 24556 21600 24565
rect 24400 24599 24452 24608
rect 24400 24565 24409 24599
rect 24409 24565 24443 24599
rect 24443 24565 24452 24599
rect 24400 24556 24452 24565
rect 3917 24454 3969 24506
rect 3981 24454 4033 24506
rect 4045 24454 4097 24506
rect 4109 24454 4161 24506
rect 4173 24454 4225 24506
rect 9851 24454 9903 24506
rect 9915 24454 9967 24506
rect 9979 24454 10031 24506
rect 10043 24454 10095 24506
rect 10107 24454 10159 24506
rect 15785 24454 15837 24506
rect 15849 24454 15901 24506
rect 15913 24454 15965 24506
rect 15977 24454 16029 24506
rect 16041 24454 16093 24506
rect 21719 24454 21771 24506
rect 21783 24454 21835 24506
rect 21847 24454 21899 24506
rect 21911 24454 21963 24506
rect 21975 24454 22027 24506
rect 2780 24352 2832 24404
rect 5908 24352 5960 24404
rect 6184 24352 6236 24404
rect 2596 24216 2648 24268
rect 388 24148 440 24200
rect 2964 24216 3016 24268
rect 4252 24216 4304 24268
rect 4804 24216 4856 24268
rect 5080 24216 5132 24268
rect 5816 24327 5868 24336
rect 5816 24293 5825 24327
rect 5825 24293 5859 24327
rect 5859 24293 5868 24327
rect 5816 24284 5868 24293
rect 5908 24216 5960 24268
rect 6368 24259 6420 24268
rect 6368 24225 6377 24259
rect 6377 24225 6411 24259
rect 6411 24225 6420 24259
rect 6368 24216 6420 24225
rect 6184 24191 6236 24200
rect 6184 24157 6218 24191
rect 6218 24157 6236 24191
rect 8576 24352 8628 24404
rect 9680 24352 9732 24404
rect 10048 24284 10100 24336
rect 6184 24148 6236 24157
rect 1584 24123 1636 24132
rect 1584 24089 1593 24123
rect 1593 24089 1627 24123
rect 1627 24089 1636 24123
rect 1584 24080 1636 24089
rect 1952 24123 2004 24132
rect 1952 24089 1961 24123
rect 1961 24089 1995 24123
rect 1995 24089 2004 24123
rect 1952 24080 2004 24089
rect 2320 24123 2372 24132
rect 2320 24089 2329 24123
rect 2329 24089 2363 24123
rect 2363 24089 2372 24123
rect 2320 24080 2372 24089
rect 2688 24055 2740 24064
rect 2688 24021 2697 24055
rect 2697 24021 2731 24055
rect 2731 24021 2740 24055
rect 2688 24012 2740 24021
rect 4620 24080 4672 24132
rect 5172 24080 5224 24132
rect 8944 24191 8996 24200
rect 8944 24157 8953 24191
rect 8953 24157 8987 24191
rect 8987 24157 8996 24191
rect 8944 24148 8996 24157
rect 9588 24148 9640 24200
rect 10784 24148 10836 24200
rect 13084 24352 13136 24404
rect 15016 24352 15068 24404
rect 13912 24284 13964 24336
rect 19248 24352 19300 24404
rect 19432 24352 19484 24404
rect 20444 24352 20496 24404
rect 21456 24352 21508 24404
rect 23388 24395 23440 24404
rect 23388 24361 23397 24395
rect 23397 24361 23431 24395
rect 23431 24361 23440 24395
rect 23388 24352 23440 24361
rect 23848 24395 23900 24404
rect 23848 24361 23857 24395
rect 23857 24361 23891 24395
rect 23891 24361 23900 24395
rect 23848 24352 23900 24361
rect 12072 24216 12124 24268
rect 14832 24216 14884 24268
rect 15660 24259 15712 24268
rect 15660 24225 15669 24259
rect 15669 24225 15703 24259
rect 15703 24225 15712 24259
rect 15660 24216 15712 24225
rect 17684 24284 17736 24336
rect 17868 24284 17920 24336
rect 18696 24284 18748 24336
rect 12348 24148 12400 24200
rect 6184 24012 6236 24064
rect 7656 24080 7708 24132
rect 11336 24080 11388 24132
rect 7564 24055 7616 24064
rect 7564 24021 7573 24055
rect 7573 24021 7607 24055
rect 7607 24021 7616 24055
rect 7564 24012 7616 24021
rect 8116 24012 8168 24064
rect 8576 24012 8628 24064
rect 9496 24012 9548 24064
rect 12164 24012 12216 24064
rect 13820 24012 13872 24064
rect 14372 24012 14424 24064
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 17316 24148 17368 24200
rect 19432 24148 19484 24200
rect 19616 24148 19668 24200
rect 19708 24191 19760 24200
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 16764 24080 16816 24132
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 23940 24191 23992 24200
rect 23940 24157 23949 24191
rect 23949 24157 23983 24191
rect 23983 24157 23992 24191
rect 23940 24148 23992 24157
rect 15476 24012 15528 24064
rect 17500 24012 17552 24064
rect 19892 24055 19944 24064
rect 19892 24021 19901 24055
rect 19901 24021 19935 24055
rect 19935 24021 19944 24055
rect 19892 24012 19944 24021
rect 25872 24080 25924 24132
rect 20628 24012 20680 24064
rect 23388 24012 23440 24064
rect 25136 24012 25188 24064
rect 6884 23910 6936 23962
rect 6948 23910 7000 23962
rect 7012 23910 7064 23962
rect 7076 23910 7128 23962
rect 7140 23910 7192 23962
rect 12818 23910 12870 23962
rect 12882 23910 12934 23962
rect 12946 23910 12998 23962
rect 13010 23910 13062 23962
rect 13074 23910 13126 23962
rect 18752 23910 18804 23962
rect 18816 23910 18868 23962
rect 18880 23910 18932 23962
rect 18944 23910 18996 23962
rect 19008 23910 19060 23962
rect 24686 23910 24738 23962
rect 24750 23910 24802 23962
rect 24814 23910 24866 23962
rect 24878 23910 24930 23962
rect 24942 23910 24994 23962
rect 2412 23808 2464 23860
rect 3516 23851 3568 23860
rect 3516 23817 3525 23851
rect 3525 23817 3559 23851
rect 3559 23817 3568 23851
rect 3516 23808 3568 23817
rect 4068 23851 4120 23860
rect 4068 23817 4077 23851
rect 4077 23817 4111 23851
rect 4111 23817 4120 23851
rect 4068 23808 4120 23817
rect 7656 23808 7708 23860
rect 2044 23672 2096 23724
rect 2228 23672 2280 23724
rect 3332 23672 3384 23724
rect 3792 23672 3844 23724
rect 3976 23672 4028 23724
rect 8116 23740 8168 23792
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 848 23536 900 23588
rect 1032 23536 1084 23588
rect 3424 23604 3476 23656
rect 5356 23604 5408 23656
rect 5448 23604 5500 23656
rect 8208 23672 8260 23724
rect 8760 23740 8812 23792
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 9956 23783 10008 23792
rect 9956 23749 9965 23783
rect 9965 23749 9999 23783
rect 9999 23749 10008 23783
rect 9956 23740 10008 23749
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 11980 23808 12032 23860
rect 12440 23808 12492 23860
rect 13452 23808 13504 23860
rect 11796 23740 11848 23792
rect 9772 23672 9824 23724
rect 11704 23672 11756 23724
rect 14832 23740 14884 23792
rect 2228 23536 2280 23588
rect 2504 23536 2556 23588
rect 3700 23536 3752 23588
rect 6460 23536 6512 23588
rect 6736 23468 6788 23520
rect 8576 23604 8628 23656
rect 10048 23604 10100 23656
rect 11152 23604 11204 23656
rect 12256 23672 12308 23724
rect 12624 23715 12676 23724
rect 12624 23681 12633 23715
rect 12633 23681 12667 23715
rect 12667 23681 12676 23715
rect 12624 23672 12676 23681
rect 13636 23715 13688 23724
rect 13636 23681 13670 23715
rect 13670 23681 13688 23715
rect 13636 23672 13688 23681
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 15660 23851 15712 23860
rect 15660 23817 15669 23851
rect 15669 23817 15703 23851
rect 15703 23817 15712 23851
rect 15660 23808 15712 23817
rect 15936 23808 15988 23860
rect 19708 23808 19760 23860
rect 12532 23604 12584 23656
rect 13176 23604 13228 23656
rect 7656 23468 7708 23520
rect 7840 23468 7892 23520
rect 8208 23468 8260 23520
rect 8392 23511 8444 23520
rect 8392 23477 8401 23511
rect 8401 23477 8435 23511
rect 8435 23477 8444 23511
rect 8392 23468 8444 23477
rect 12072 23511 12124 23520
rect 12072 23477 12081 23511
rect 12081 23477 12115 23511
rect 12115 23477 12124 23511
rect 12072 23468 12124 23477
rect 13268 23468 13320 23520
rect 14004 23604 14056 23656
rect 16488 23740 16540 23792
rect 22376 23808 22428 23860
rect 23296 23808 23348 23860
rect 17868 23715 17920 23724
rect 17868 23681 17877 23715
rect 17877 23681 17911 23715
rect 17911 23681 17920 23715
rect 17868 23672 17920 23681
rect 18512 23672 18564 23724
rect 19524 23672 19576 23724
rect 20536 23672 20588 23724
rect 21640 23672 21692 23724
rect 22744 23672 22796 23724
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 23940 23715 23992 23724
rect 23940 23681 23949 23715
rect 23949 23681 23983 23715
rect 23983 23681 23992 23715
rect 23940 23672 23992 23681
rect 14004 23468 14056 23520
rect 14280 23468 14332 23520
rect 19616 23468 19668 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 23572 23511 23624 23520
rect 23572 23477 23581 23511
rect 23581 23477 23615 23511
rect 23615 23477 23624 23511
rect 23572 23468 23624 23477
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 3917 23366 3969 23418
rect 3981 23366 4033 23418
rect 4045 23366 4097 23418
rect 4109 23366 4161 23418
rect 4173 23366 4225 23418
rect 9851 23366 9903 23418
rect 9915 23366 9967 23418
rect 9979 23366 10031 23418
rect 10043 23366 10095 23418
rect 10107 23366 10159 23418
rect 15785 23366 15837 23418
rect 15849 23366 15901 23418
rect 15913 23366 15965 23418
rect 15977 23366 16029 23418
rect 16041 23366 16093 23418
rect 21719 23366 21771 23418
rect 21783 23366 21835 23418
rect 21847 23366 21899 23418
rect 21911 23366 21963 23418
rect 21975 23366 22027 23418
rect 2044 23264 2096 23316
rect 2228 23307 2280 23316
rect 2228 23273 2237 23307
rect 2237 23273 2271 23307
rect 2271 23273 2280 23307
rect 2228 23264 2280 23273
rect 2596 23264 2648 23316
rect 3240 23264 3292 23316
rect 9220 23264 9272 23316
rect 12348 23264 12400 23316
rect 1032 23060 1084 23112
rect 848 22992 900 23044
rect 2504 22992 2556 23044
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 11060 23128 11112 23180
rect 14832 23264 14884 23316
rect 15016 23264 15068 23316
rect 16764 23264 16816 23316
rect 19892 23264 19944 23316
rect 23940 23264 23992 23316
rect 3332 23060 3384 23112
rect 3332 22924 3384 22976
rect 4160 23060 4212 23112
rect 6000 23060 6052 23112
rect 6184 23060 6236 23112
rect 6552 23060 6604 23112
rect 7564 23060 7616 23112
rect 8392 23060 8444 23112
rect 8944 23103 8996 23112
rect 8944 23069 8953 23103
rect 8953 23069 8987 23103
rect 8987 23069 8996 23103
rect 8944 23060 8996 23069
rect 4252 22924 4304 22976
rect 6736 22992 6788 23044
rect 10048 22992 10100 23044
rect 4896 22924 4948 22976
rect 9404 22924 9456 22976
rect 10876 23103 10928 23112
rect 10876 23069 10885 23103
rect 10885 23069 10919 23103
rect 10919 23069 10928 23103
rect 10876 23060 10928 23069
rect 12164 23060 12216 23112
rect 14280 23060 14332 23112
rect 15108 23060 15160 23112
rect 16764 23060 16816 23112
rect 17408 23060 17460 23112
rect 18512 23060 18564 23112
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 19984 23060 20036 23112
rect 20628 23103 20680 23112
rect 20628 23069 20637 23103
rect 20637 23069 20671 23103
rect 20671 23069 20680 23103
rect 20628 23060 20680 23069
rect 11152 22992 11204 23044
rect 11336 23035 11388 23044
rect 11336 23001 11345 23035
rect 11345 23001 11379 23035
rect 11379 23001 11388 23035
rect 11336 22992 11388 23001
rect 11428 22992 11480 23044
rect 11796 22992 11848 23044
rect 19432 22992 19484 23044
rect 20720 22992 20772 23044
rect 21732 23060 21784 23112
rect 22376 23103 22428 23112
rect 22376 23069 22385 23103
rect 22385 23069 22419 23103
rect 22419 23069 22428 23103
rect 22376 23060 22428 23069
rect 23756 23060 23808 23112
rect 22744 22992 22796 23044
rect 11520 22924 11572 22976
rect 11888 22967 11940 22976
rect 11888 22933 11897 22967
rect 11897 22933 11931 22967
rect 11931 22933 11940 22967
rect 11888 22924 11940 22933
rect 14556 22924 14608 22976
rect 15108 22967 15160 22976
rect 15108 22933 15117 22967
rect 15117 22933 15151 22967
rect 15151 22933 15160 22967
rect 15108 22924 15160 22933
rect 17132 22924 17184 22976
rect 17408 22924 17460 22976
rect 21364 22924 21416 22976
rect 22100 22924 22152 22976
rect 22192 22967 22244 22976
rect 22192 22933 22201 22967
rect 22201 22933 22235 22967
rect 22235 22933 22244 22967
rect 22192 22924 22244 22933
rect 25136 22924 25188 22976
rect 6884 22822 6936 22874
rect 6948 22822 7000 22874
rect 7012 22822 7064 22874
rect 7076 22822 7128 22874
rect 7140 22822 7192 22874
rect 12818 22822 12870 22874
rect 12882 22822 12934 22874
rect 12946 22822 12998 22874
rect 13010 22822 13062 22874
rect 13074 22822 13126 22874
rect 18752 22822 18804 22874
rect 18816 22822 18868 22874
rect 18880 22822 18932 22874
rect 18944 22822 18996 22874
rect 19008 22822 19060 22874
rect 24686 22822 24738 22874
rect 24750 22822 24802 22874
rect 24814 22822 24866 22874
rect 24878 22822 24930 22874
rect 24942 22822 24994 22874
rect 2688 22720 2740 22772
rect 1308 22652 1360 22704
rect 3516 22720 3568 22772
rect 6092 22720 6144 22772
rect 8116 22720 8168 22772
rect 10784 22720 10836 22772
rect 11060 22763 11112 22772
rect 11060 22729 11069 22763
rect 11069 22729 11103 22763
rect 11103 22729 11112 22763
rect 11060 22720 11112 22729
rect 11428 22720 11480 22772
rect 12256 22720 12308 22772
rect 13820 22720 13872 22772
rect 14464 22720 14516 22772
rect 14740 22720 14792 22772
rect 15384 22720 15436 22772
rect 19432 22720 19484 22772
rect 19892 22720 19944 22772
rect 20720 22720 20772 22772
rect 21732 22720 21784 22772
rect 22284 22720 22336 22772
rect 23204 22720 23256 22772
rect 848 22584 900 22636
rect 2872 22584 2924 22636
rect 5448 22652 5500 22704
rect 7840 22652 7892 22704
rect 6736 22584 6788 22636
rect 9680 22584 9732 22636
rect 10324 22623 10349 22636
rect 10349 22623 10376 22636
rect 1400 22448 1452 22500
rect 2596 22448 2648 22500
rect 4068 22448 4120 22500
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 6184 22516 6236 22568
rect 4896 22380 4948 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 6736 22380 6788 22432
rect 10324 22584 10376 22623
rect 12624 22584 12676 22636
rect 12900 22584 12952 22636
rect 13176 22652 13228 22704
rect 13452 22652 13504 22704
rect 16672 22652 16724 22704
rect 16580 22584 16632 22636
rect 17776 22584 17828 22636
rect 22744 22652 22796 22704
rect 16764 22516 16816 22568
rect 17316 22491 17368 22500
rect 17316 22457 17325 22491
rect 17325 22457 17359 22491
rect 17359 22457 17368 22491
rect 17316 22448 17368 22457
rect 10968 22380 11020 22432
rect 12348 22380 12400 22432
rect 12624 22380 12676 22432
rect 14832 22423 14884 22432
rect 14832 22389 14841 22423
rect 14841 22389 14875 22423
rect 14875 22389 14884 22423
rect 14832 22380 14884 22389
rect 15660 22380 15712 22432
rect 16948 22380 17000 22432
rect 17868 22559 17920 22568
rect 17868 22525 17877 22559
rect 17877 22525 17911 22559
rect 17911 22525 17920 22559
rect 17868 22516 17920 22525
rect 21640 22627 21692 22636
rect 21640 22593 21649 22627
rect 21649 22593 21683 22627
rect 21683 22593 21692 22627
rect 21640 22584 21692 22593
rect 21732 22516 21784 22568
rect 19984 22448 20036 22500
rect 22008 22584 22060 22636
rect 22652 22584 22704 22636
rect 23480 22627 23532 22636
rect 23480 22593 23487 22627
rect 23487 22593 23521 22627
rect 23521 22593 23532 22627
rect 23480 22584 23532 22593
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 19248 22380 19300 22432
rect 20628 22380 20680 22432
rect 22284 22380 22336 22432
rect 22836 22423 22888 22432
rect 22836 22389 22845 22423
rect 22845 22389 22879 22423
rect 22879 22389 22888 22423
rect 22836 22380 22888 22389
rect 3917 22278 3969 22330
rect 3981 22278 4033 22330
rect 4045 22278 4097 22330
rect 4109 22278 4161 22330
rect 4173 22278 4225 22330
rect 9851 22278 9903 22330
rect 9915 22278 9967 22330
rect 9979 22278 10031 22330
rect 10043 22278 10095 22330
rect 10107 22278 10159 22330
rect 15785 22278 15837 22330
rect 15849 22278 15901 22330
rect 15913 22278 15965 22330
rect 15977 22278 16029 22330
rect 16041 22278 16093 22330
rect 21719 22278 21771 22330
rect 21783 22278 21835 22330
rect 21847 22278 21899 22330
rect 21911 22278 21963 22330
rect 21975 22278 22027 22330
rect 3056 22219 3108 22228
rect 3056 22185 3065 22219
rect 3065 22185 3099 22219
rect 3099 22185 3108 22219
rect 3056 22176 3108 22185
rect 3608 22176 3660 22228
rect 3792 22176 3844 22228
rect 6000 22151 6052 22160
rect 6000 22117 6009 22151
rect 6009 22117 6043 22151
rect 6043 22117 6052 22151
rect 6000 22108 6052 22117
rect 6552 22151 6604 22160
rect 6552 22117 6561 22151
rect 6561 22117 6595 22151
rect 6595 22117 6604 22151
rect 6552 22108 6604 22117
rect 8484 22108 8536 22160
rect 9496 22108 9548 22160
rect 2320 22040 2372 22092
rect 5172 22040 5224 22092
rect 6184 22040 6236 22092
rect 9404 22040 9456 22092
rect 9864 22040 9916 22092
rect 12900 22219 12952 22228
rect 12900 22185 12909 22219
rect 12909 22185 12943 22219
rect 12943 22185 12952 22219
rect 12900 22176 12952 22185
rect 13636 22176 13688 22228
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 14832 22040 14884 22092
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 17316 22219 17368 22228
rect 17316 22185 17325 22219
rect 17325 22185 17359 22219
rect 17359 22185 17368 22219
rect 17316 22176 17368 22185
rect 18512 22176 18564 22228
rect 22192 22176 22244 22228
rect 1032 21972 1084 22024
rect 1216 21972 1268 22024
rect 2412 21972 2464 22024
rect 3148 21972 3200 22024
rect 3240 22015 3292 22024
rect 3240 21981 3249 22015
rect 3249 21981 3283 22015
rect 3283 21981 3292 22015
rect 3240 21972 3292 21981
rect 1768 21947 1820 21956
rect 1768 21913 1777 21947
rect 1777 21913 1811 21947
rect 1811 21913 1820 21947
rect 1768 21904 1820 21913
rect 2044 21947 2096 21956
rect 2044 21913 2053 21947
rect 2053 21913 2087 21947
rect 2087 21913 2096 21947
rect 2044 21904 2096 21913
rect 1216 21836 1268 21888
rect 3976 21904 4028 21956
rect 5080 21947 5132 21956
rect 5080 21913 5089 21947
rect 5089 21913 5123 21947
rect 5123 21913 5132 21947
rect 5080 21904 5132 21913
rect 5448 22015 5500 22024
rect 5448 21981 5457 22015
rect 5457 21981 5491 22015
rect 5491 21981 5500 22015
rect 5448 21972 5500 21981
rect 5816 22015 5868 22024
rect 5816 21981 5839 22015
rect 5839 21981 5868 22015
rect 5816 21972 5868 21981
rect 6552 21972 6604 22024
rect 6828 21972 6880 22024
rect 8208 21972 8260 22024
rect 8576 21972 8628 22024
rect 9036 21972 9088 22024
rect 2872 21879 2924 21888
rect 2872 21845 2881 21879
rect 2881 21845 2915 21879
rect 2915 21845 2924 21879
rect 2872 21836 2924 21845
rect 3148 21836 3200 21888
rect 4620 21836 4672 21888
rect 5632 21904 5684 21956
rect 13360 21972 13412 22024
rect 5908 21836 5960 21888
rect 6184 21836 6236 21888
rect 7380 21836 7432 21888
rect 8392 21836 8444 21888
rect 8668 21836 8720 21888
rect 9772 21836 9824 21888
rect 11244 21836 11296 21888
rect 11796 21904 11848 21956
rect 11980 21947 12032 21956
rect 11980 21913 11989 21947
rect 11989 21913 12023 21947
rect 12023 21913 12032 21947
rect 11980 21904 12032 21913
rect 12072 21904 12124 21956
rect 15108 22015 15160 22024
rect 15108 21981 15142 22015
rect 15142 21981 15160 22015
rect 15108 21972 15160 21981
rect 16120 21972 16172 22024
rect 16488 21972 16540 22024
rect 17224 21972 17276 22024
rect 21640 22108 21692 22160
rect 22836 22176 22888 22228
rect 23572 22176 23624 22228
rect 19248 22083 19300 22092
rect 19248 22049 19257 22083
rect 19257 22049 19291 22083
rect 19291 22049 19300 22083
rect 19248 22040 19300 22049
rect 20352 22040 20404 22092
rect 20260 21972 20312 22024
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 15384 21836 15436 21888
rect 17684 21836 17736 21888
rect 18604 21836 18656 21888
rect 19616 21904 19668 21956
rect 20444 21904 20496 21956
rect 20720 21904 20772 21956
rect 22468 22108 22520 22160
rect 25688 22108 25740 22160
rect 22284 22083 22336 22092
rect 22284 22049 22293 22083
rect 22293 22049 22327 22083
rect 22327 22049 22336 22083
rect 22284 22040 22336 22049
rect 23296 22040 23348 22092
rect 22100 21972 22152 22024
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 25688 21972 25740 22024
rect 23480 21904 23532 21956
rect 25136 21904 25188 21956
rect 20904 21836 20956 21888
rect 20996 21879 21048 21888
rect 20996 21845 21005 21879
rect 21005 21845 21039 21879
rect 21039 21845 21048 21879
rect 20996 21836 21048 21845
rect 21364 21836 21416 21888
rect 21640 21836 21692 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 23388 21879 23440 21888
rect 23388 21845 23397 21879
rect 23397 21845 23431 21879
rect 23431 21845 23440 21879
rect 23388 21836 23440 21845
rect 23756 21836 23808 21888
rect 6884 21734 6936 21786
rect 6948 21734 7000 21786
rect 7012 21734 7064 21786
rect 7076 21734 7128 21786
rect 7140 21734 7192 21786
rect 12818 21734 12870 21786
rect 12882 21734 12934 21786
rect 12946 21734 12998 21786
rect 13010 21734 13062 21786
rect 13074 21734 13126 21786
rect 18752 21734 18804 21786
rect 18816 21734 18868 21786
rect 18880 21734 18932 21786
rect 18944 21734 18996 21786
rect 19008 21734 19060 21786
rect 24686 21734 24738 21786
rect 24750 21734 24802 21786
rect 24814 21734 24866 21786
rect 24878 21734 24930 21786
rect 24942 21734 24994 21786
rect 848 21632 900 21684
rect 1768 21632 1820 21684
rect 2320 21632 2372 21684
rect 2504 21632 2556 21684
rect 1308 21564 1360 21616
rect 4160 21632 4212 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 2596 21496 2648 21548
rect 3976 21564 4028 21616
rect 5080 21632 5132 21684
rect 5172 21632 5224 21684
rect 6184 21632 6236 21684
rect 7104 21632 7156 21684
rect 6644 21564 6696 21616
rect 7380 21564 7432 21616
rect 7656 21607 7708 21616
rect 7656 21573 7665 21607
rect 7665 21573 7699 21607
rect 7699 21573 7708 21607
rect 7656 21564 7708 21573
rect 8484 21675 8536 21684
rect 8484 21641 8493 21675
rect 8493 21641 8527 21675
rect 8527 21641 8536 21675
rect 8484 21632 8536 21641
rect 9680 21632 9732 21684
rect 11060 21632 11112 21684
rect 11980 21632 12032 21684
rect 14740 21632 14792 21684
rect 20352 21632 20404 21684
rect 20812 21632 20864 21684
rect 4896 21496 4948 21548
rect 5908 21496 5960 21548
rect 6092 21496 6144 21548
rect 8668 21496 8720 21548
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 9220 21539 9272 21548
rect 9220 21505 9229 21539
rect 9229 21505 9263 21539
rect 9263 21505 9272 21539
rect 9220 21496 9272 21505
rect 9404 21496 9456 21548
rect 15200 21564 15252 21616
rect 12624 21496 12676 21548
rect 13636 21496 13688 21548
rect 14280 21496 14332 21548
rect 15016 21496 15068 21548
rect 15384 21539 15436 21548
rect 15384 21505 15391 21539
rect 15391 21505 15425 21539
rect 15425 21505 15436 21539
rect 15384 21496 15436 21505
rect 15476 21496 15528 21548
rect 15844 21496 15896 21548
rect 16120 21564 16172 21616
rect 16764 21564 16816 21616
rect 18604 21564 18656 21616
rect 6736 21428 6788 21480
rect 8484 21428 8536 21480
rect 9588 21428 9640 21480
rect 11336 21428 11388 21480
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 1308 21292 1360 21344
rect 4528 21360 4580 21412
rect 3700 21292 3752 21344
rect 4344 21292 4396 21344
rect 5816 21292 5868 21344
rect 8392 21292 8444 21344
rect 11428 21292 11480 21344
rect 13544 21292 13596 21344
rect 15016 21335 15068 21344
rect 15016 21301 15025 21335
rect 15025 21301 15059 21335
rect 15059 21301 15068 21335
rect 15016 21292 15068 21301
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 17776 21496 17828 21548
rect 19616 21564 19668 21616
rect 19984 21564 20036 21616
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 19064 21360 19116 21412
rect 19800 21360 19852 21412
rect 20260 21496 20312 21548
rect 20996 21632 21048 21684
rect 21272 21632 21324 21684
rect 22284 21632 22336 21684
rect 24492 21632 24544 21684
rect 21456 21496 21508 21548
rect 23572 21539 23624 21548
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 24216 21496 24268 21548
rect 23756 21428 23808 21480
rect 23664 21360 23716 21412
rect 17132 21292 17184 21344
rect 17224 21292 17276 21344
rect 17776 21292 17828 21344
rect 18788 21292 18840 21344
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 23848 21335 23900 21344
rect 23848 21301 23857 21335
rect 23857 21301 23891 21335
rect 23891 21301 23900 21335
rect 23848 21292 23900 21301
rect 3917 21190 3969 21242
rect 3981 21190 4033 21242
rect 4045 21190 4097 21242
rect 4109 21190 4161 21242
rect 4173 21190 4225 21242
rect 9851 21190 9903 21242
rect 9915 21190 9967 21242
rect 9979 21190 10031 21242
rect 10043 21190 10095 21242
rect 10107 21190 10159 21242
rect 15785 21190 15837 21242
rect 15849 21190 15901 21242
rect 15913 21190 15965 21242
rect 15977 21190 16029 21242
rect 16041 21190 16093 21242
rect 21719 21190 21771 21242
rect 21783 21190 21835 21242
rect 21847 21190 21899 21242
rect 21911 21190 21963 21242
rect 21975 21190 22027 21242
rect 7104 21088 7156 21140
rect 2964 21020 3016 21072
rect 1216 20952 1268 21004
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 8852 21088 8904 21140
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 1768 20884 1820 20936
rect 1308 20816 1360 20868
rect 2136 20748 2188 20800
rect 3976 20884 4028 20936
rect 3332 20816 3384 20868
rect 8208 20952 8260 21004
rect 8484 20952 8536 21004
rect 8944 20995 8996 21004
rect 8944 20961 8953 20995
rect 8953 20961 8987 20995
rect 8987 20961 8996 20995
rect 8944 20952 8996 20961
rect 9772 20952 9824 21004
rect 10140 20952 10192 21004
rect 5080 20884 5132 20936
rect 5632 20884 5684 20936
rect 5908 20884 5960 20936
rect 7840 20884 7892 20936
rect 4068 20748 4120 20800
rect 6092 20748 6144 20800
rect 6368 20748 6420 20800
rect 9128 20884 9180 20936
rect 9864 20884 9916 20936
rect 8944 20816 8996 20868
rect 15016 21020 15068 21072
rect 17868 21088 17920 21140
rect 19340 21088 19392 21140
rect 19616 21088 19668 21140
rect 21364 21088 21416 21140
rect 11796 20952 11848 21004
rect 11980 20995 12032 21004
rect 11980 20961 11989 20995
rect 11989 20961 12023 20995
rect 12023 20961 12032 20995
rect 11980 20952 12032 20961
rect 13360 20952 13412 21004
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 15752 20995 15804 21004
rect 15752 20961 15786 20995
rect 15786 20961 15804 20995
rect 15752 20952 15804 20961
rect 16120 20952 16172 21004
rect 16764 20952 16816 21004
rect 16948 20995 17000 21004
rect 16948 20961 16957 20995
rect 16957 20961 16991 20995
rect 16991 20961 17000 20995
rect 16948 20952 17000 20961
rect 11152 20884 11204 20936
rect 12164 20884 12216 20936
rect 14832 20884 14884 20936
rect 16672 20884 16724 20936
rect 18788 20952 18840 21004
rect 19064 20952 19116 21004
rect 19156 20884 19208 20936
rect 11060 20816 11112 20868
rect 11520 20816 11572 20868
rect 12624 20816 12676 20868
rect 13636 20816 13688 20868
rect 20720 21063 20772 21072
rect 20720 21029 20729 21063
rect 20729 21029 20763 21063
rect 20763 21029 20772 21063
rect 20720 21020 20772 21029
rect 20904 21020 20956 21072
rect 22376 20884 22428 20936
rect 22468 20884 22520 20936
rect 20168 20816 20220 20868
rect 21180 20816 21232 20868
rect 22652 20816 22704 20868
rect 8208 20748 8260 20800
rect 9128 20748 9180 20800
rect 9680 20748 9732 20800
rect 10140 20748 10192 20800
rect 10692 20748 10744 20800
rect 10968 20748 11020 20800
rect 12716 20748 12768 20800
rect 13452 20748 13504 20800
rect 13820 20748 13872 20800
rect 14096 20748 14148 20800
rect 15108 20748 15160 20800
rect 20812 20748 20864 20800
rect 23296 20748 23348 20800
rect 24216 20748 24268 20800
rect 6884 20646 6936 20698
rect 6948 20646 7000 20698
rect 7012 20646 7064 20698
rect 7076 20646 7128 20698
rect 7140 20646 7192 20698
rect 12818 20646 12870 20698
rect 12882 20646 12934 20698
rect 12946 20646 12998 20698
rect 13010 20646 13062 20698
rect 13074 20646 13126 20698
rect 18752 20646 18804 20698
rect 18816 20646 18868 20698
rect 18880 20646 18932 20698
rect 18944 20646 18996 20698
rect 19008 20646 19060 20698
rect 24686 20646 24738 20698
rect 24750 20646 24802 20698
rect 24814 20646 24866 20698
rect 24878 20646 24930 20698
rect 24942 20646 24994 20698
rect 3976 20544 4028 20596
rect 7840 20544 7892 20596
rect 2044 20408 2096 20460
rect 2596 20408 2648 20460
rect 3792 20451 3844 20460
rect 3792 20417 3801 20451
rect 3801 20417 3835 20451
rect 3835 20417 3844 20451
rect 3792 20408 3844 20417
rect 3884 20451 3936 20460
rect 3884 20417 3918 20451
rect 3918 20417 3936 20451
rect 3884 20408 3936 20417
rect 4068 20451 4120 20460
rect 4068 20417 4077 20451
rect 4077 20417 4111 20451
rect 4111 20417 4120 20451
rect 4068 20408 4120 20417
rect 4896 20476 4948 20528
rect 6644 20476 6696 20528
rect 9956 20519 10008 20528
rect 9956 20485 9965 20519
rect 9965 20485 9999 20519
rect 9999 20485 10008 20519
rect 9956 20476 10008 20485
rect 10232 20519 10284 20528
rect 10232 20485 10241 20519
rect 10241 20485 10275 20519
rect 10275 20485 10284 20519
rect 10232 20476 10284 20485
rect 10508 20476 10560 20528
rect 11244 20544 11296 20596
rect 11152 20476 11204 20528
rect 12532 20544 12584 20596
rect 15384 20587 15436 20596
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 16672 20544 16724 20596
rect 17132 20544 17184 20596
rect 19156 20544 19208 20596
rect 19432 20544 19484 20596
rect 19616 20544 19668 20596
rect 20444 20544 20496 20596
rect 22468 20587 22520 20596
rect 22468 20553 22477 20587
rect 22477 20553 22511 20587
rect 22511 20553 22520 20587
rect 22468 20544 22520 20553
rect 23756 20587 23808 20596
rect 23756 20553 23765 20587
rect 23765 20553 23799 20587
rect 23799 20553 23808 20587
rect 23756 20544 23808 20553
rect 11796 20476 11848 20528
rect 12440 20476 12492 20528
rect 8576 20408 8628 20460
rect 10600 20408 10652 20460
rect 15108 20476 15160 20528
rect 18236 20476 18288 20528
rect 13360 20451 13412 20460
rect 13360 20417 13394 20451
rect 13394 20417 13412 20451
rect 13360 20408 13412 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 14280 20408 14332 20460
rect 14556 20408 14608 20460
rect 14740 20408 14792 20460
rect 16948 20408 17000 20460
rect 22100 20408 22152 20460
rect 22652 20451 22704 20460
rect 22652 20417 22661 20451
rect 22661 20417 22695 20451
rect 22695 20417 22704 20451
rect 22652 20408 22704 20417
rect 22744 20451 22796 20460
rect 22744 20417 22753 20451
rect 22753 20417 22787 20451
rect 22787 20417 22796 20451
rect 22744 20408 22796 20417
rect 22928 20408 22980 20460
rect 24216 20451 24268 20460
rect 24216 20417 24225 20451
rect 24225 20417 24259 20451
rect 24259 20417 24268 20451
rect 24216 20408 24268 20417
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 3148 20340 3200 20392
rect 3516 20315 3568 20324
rect 3516 20281 3525 20315
rect 3525 20281 3559 20315
rect 3559 20281 3568 20315
rect 3516 20272 3568 20281
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 10968 20340 11020 20392
rect 11336 20340 11388 20392
rect 12256 20340 12308 20392
rect 9404 20272 9456 20324
rect 11244 20315 11296 20324
rect 11244 20281 11253 20315
rect 11253 20281 11287 20315
rect 11287 20281 11296 20315
rect 11244 20272 11296 20281
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 5816 20204 5868 20213
rect 5908 20204 5960 20256
rect 7288 20204 7340 20256
rect 11336 20204 11388 20256
rect 12716 20340 12768 20392
rect 13912 20340 13964 20392
rect 14188 20340 14240 20392
rect 22284 20340 22336 20392
rect 23480 20340 23532 20392
rect 22652 20272 22704 20324
rect 14832 20204 14884 20256
rect 16396 20204 16448 20256
rect 18512 20204 18564 20256
rect 22836 20204 22888 20256
rect 23848 20204 23900 20256
rect 24308 20247 24360 20256
rect 24308 20213 24317 20247
rect 24317 20213 24351 20247
rect 24351 20213 24360 20247
rect 24308 20204 24360 20213
rect 3917 20102 3969 20154
rect 3981 20102 4033 20154
rect 4045 20102 4097 20154
rect 4109 20102 4161 20154
rect 4173 20102 4225 20154
rect 9851 20102 9903 20154
rect 9915 20102 9967 20154
rect 9979 20102 10031 20154
rect 10043 20102 10095 20154
rect 10107 20102 10159 20154
rect 15785 20102 15837 20154
rect 15849 20102 15901 20154
rect 15913 20102 15965 20154
rect 15977 20102 16029 20154
rect 16041 20102 16093 20154
rect 21719 20102 21771 20154
rect 21783 20102 21835 20154
rect 21847 20102 21899 20154
rect 21911 20102 21963 20154
rect 21975 20102 22027 20154
rect 1860 20000 1912 20052
rect 3516 20000 3568 20052
rect 4344 20000 4396 20052
rect 9772 20000 9824 20052
rect 10600 20000 10652 20052
rect 11980 20000 12032 20052
rect 2136 19864 2188 19916
rect 756 19796 808 19848
rect 2044 19796 2096 19848
rect 5816 19864 5868 19916
rect 7656 19864 7708 19916
rect 8024 19864 8076 19916
rect 13268 20000 13320 20052
rect 13544 20043 13596 20052
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 14280 20000 14332 20052
rect 16120 20000 16172 20052
rect 16580 20000 16632 20052
rect 14464 19932 14516 19984
rect 15384 19932 15436 19984
rect 20904 20000 20956 20052
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 16396 19864 16448 19916
rect 17776 19932 17828 19984
rect 17684 19864 17736 19916
rect 19248 19907 19300 19916
rect 19248 19873 19257 19907
rect 19257 19873 19291 19907
rect 19291 19873 19300 19907
rect 19248 19864 19300 19873
rect 1308 19728 1360 19780
rect 5632 19796 5684 19848
rect 7288 19796 7340 19848
rect 7380 19796 7432 19848
rect 10876 19796 10928 19848
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12860 19839
rect 12808 19796 12860 19805
rect 14280 19796 14332 19848
rect 4988 19728 5040 19780
rect 5356 19728 5408 19780
rect 5816 19728 5868 19780
rect 6736 19728 6788 19780
rect 6828 19728 6880 19780
rect 6460 19703 6512 19712
rect 6460 19669 6469 19703
rect 6469 19669 6503 19703
rect 6503 19669 6512 19703
rect 6460 19660 6512 19669
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 9128 19728 9180 19780
rect 15016 19728 15068 19780
rect 16856 19839 16908 19848
rect 16856 19805 16865 19839
rect 16865 19805 16899 19839
rect 16899 19805 16908 19839
rect 16856 19796 16908 19805
rect 20812 19796 20864 19848
rect 21272 19796 21324 19848
rect 22100 20043 22152 20052
rect 22100 20009 22109 20043
rect 22109 20009 22143 20043
rect 22143 20009 22152 20043
rect 22100 20000 22152 20009
rect 22284 20000 22336 20052
rect 22468 20000 22520 20052
rect 24032 20000 24084 20052
rect 23664 19839 23716 19848
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 21088 19728 21140 19780
rect 24216 19728 24268 19780
rect 11336 19660 11388 19712
rect 12716 19660 12768 19712
rect 14096 19660 14148 19712
rect 16948 19660 17000 19712
rect 18144 19660 18196 19712
rect 19156 19660 19208 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 6884 19558 6936 19610
rect 6948 19558 7000 19610
rect 7012 19558 7064 19610
rect 7076 19558 7128 19610
rect 7140 19558 7192 19610
rect 12818 19558 12870 19610
rect 12882 19558 12934 19610
rect 12946 19558 12998 19610
rect 13010 19558 13062 19610
rect 13074 19558 13126 19610
rect 18752 19558 18804 19610
rect 18816 19558 18868 19610
rect 18880 19558 18932 19610
rect 18944 19558 18996 19610
rect 19008 19558 19060 19610
rect 24686 19558 24738 19610
rect 24750 19558 24802 19610
rect 24814 19558 24866 19610
rect 24878 19558 24930 19610
rect 24942 19558 24994 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 1952 19456 2004 19508
rect 4620 19456 4672 19508
rect 4712 19456 4764 19508
rect 5816 19456 5868 19508
rect 6368 19456 6420 19508
rect 7748 19456 7800 19508
rect 8208 19499 8260 19508
rect 8208 19465 8217 19499
rect 8217 19465 8251 19499
rect 8251 19465 8260 19499
rect 8208 19456 8260 19465
rect 848 19320 900 19372
rect 1860 19320 1912 19372
rect 2044 19320 2096 19372
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 3792 19320 3844 19372
rect 4620 19320 4672 19372
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 4896 19320 4948 19329
rect 7196 19320 7248 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 7840 19431 7892 19440
rect 7840 19397 7849 19431
rect 7849 19397 7883 19431
rect 7883 19397 7892 19431
rect 7840 19388 7892 19397
rect 9128 19456 9180 19508
rect 9220 19456 9272 19508
rect 14280 19456 14332 19508
rect 16856 19456 16908 19508
rect 19248 19456 19300 19508
rect 19984 19456 20036 19508
rect 8024 19320 8076 19372
rect 12716 19388 12768 19440
rect 13544 19388 13596 19440
rect 13912 19388 13964 19440
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 7656 19252 7708 19304
rect 10600 19320 10652 19372
rect 11796 19363 11848 19372
rect 11796 19329 11803 19363
rect 11803 19329 11837 19363
rect 11837 19329 11848 19363
rect 11796 19320 11848 19329
rect 16396 19320 16448 19372
rect 11244 19252 11296 19304
rect 11520 19295 11572 19304
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 5816 19116 5868 19168
rect 8300 19116 8352 19168
rect 11060 19184 11112 19236
rect 9680 19116 9732 19168
rect 10140 19116 10192 19168
rect 10416 19116 10468 19168
rect 12532 19159 12584 19168
rect 12532 19125 12541 19159
rect 12541 19125 12575 19159
rect 12575 19125 12584 19159
rect 12532 19116 12584 19125
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 16120 19116 16172 19168
rect 19064 19320 19116 19372
rect 19800 19388 19852 19440
rect 19432 19363 19484 19372
rect 19432 19329 19439 19363
rect 19439 19329 19473 19363
rect 19473 19329 19484 19363
rect 19432 19320 19484 19329
rect 21088 19456 21140 19508
rect 20444 19388 20496 19440
rect 22192 19456 22244 19508
rect 23204 19456 23256 19508
rect 23296 19456 23348 19508
rect 23572 19456 23624 19508
rect 23848 19456 23900 19508
rect 21272 19320 21324 19372
rect 22652 19363 22704 19372
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 22928 19320 22980 19372
rect 23296 19252 23348 19304
rect 24124 19431 24176 19440
rect 24124 19397 24133 19431
rect 24133 19397 24167 19431
rect 24167 19397 24176 19431
rect 24124 19388 24176 19397
rect 25504 19320 25556 19372
rect 25136 19252 25188 19304
rect 25504 19184 25556 19236
rect 20260 19116 20312 19168
rect 20812 19116 20864 19168
rect 23848 19159 23900 19168
rect 23848 19125 23857 19159
rect 23857 19125 23891 19159
rect 23891 19125 23900 19159
rect 23848 19116 23900 19125
rect 3917 19014 3969 19066
rect 3981 19014 4033 19066
rect 4045 19014 4097 19066
rect 4109 19014 4161 19066
rect 4173 19014 4225 19066
rect 9851 19014 9903 19066
rect 9915 19014 9967 19066
rect 9979 19014 10031 19066
rect 10043 19014 10095 19066
rect 10107 19014 10159 19066
rect 15785 19014 15837 19066
rect 15849 19014 15901 19066
rect 15913 19014 15965 19066
rect 15977 19014 16029 19066
rect 16041 19014 16093 19066
rect 21719 19014 21771 19066
rect 21783 19014 21835 19066
rect 21847 19014 21899 19066
rect 21911 19014 21963 19066
rect 21975 19014 22027 19066
rect 1400 18912 1452 18964
rect 4528 18912 4580 18964
rect 7472 18912 7524 18964
rect 10508 18912 10560 18964
rect 12716 18912 12768 18964
rect 16120 18912 16172 18964
rect 16304 18912 16356 18964
rect 20260 18912 20312 18964
rect 20444 18912 20496 18964
rect 21548 18912 21600 18964
rect 4620 18844 4672 18896
rect 5908 18844 5960 18896
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 6736 18776 6788 18828
rect 9128 18776 9180 18828
rect 14464 18776 14516 18828
rect 19156 18776 19208 18828
rect 23480 18844 23532 18896
rect 25136 18844 25188 18896
rect 2320 18708 2372 18760
rect 1308 18640 1360 18692
rect 3976 18708 4028 18760
rect 4528 18708 4580 18760
rect 4712 18708 4764 18760
rect 6368 18708 6420 18760
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 9680 18708 9732 18760
rect 9772 18708 9824 18760
rect 10416 18708 10468 18760
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 7104 18640 7156 18692
rect 7840 18640 7892 18692
rect 9956 18640 10008 18692
rect 2872 18572 2924 18624
rect 4068 18572 4120 18624
rect 4804 18615 4856 18624
rect 4804 18581 4813 18615
rect 4813 18581 4847 18615
rect 4847 18581 4856 18615
rect 4804 18572 4856 18581
rect 8668 18572 8720 18624
rect 10876 18640 10928 18692
rect 11428 18640 11480 18692
rect 10416 18615 10468 18624
rect 10416 18581 10425 18615
rect 10425 18581 10459 18615
rect 10459 18581 10468 18615
rect 10416 18572 10468 18581
rect 14924 18708 14976 18760
rect 15016 18751 15068 18760
rect 15016 18717 15025 18751
rect 15025 18717 15059 18751
rect 15059 18717 15068 18751
rect 15016 18708 15068 18717
rect 16212 18708 16264 18760
rect 17132 18708 17184 18760
rect 11980 18572 12032 18624
rect 12256 18615 12308 18624
rect 12256 18581 12265 18615
rect 12265 18581 12299 18615
rect 12299 18581 12308 18615
rect 12256 18572 12308 18581
rect 14280 18683 14332 18692
rect 14280 18649 14289 18683
rect 14289 18649 14323 18683
rect 14323 18649 14332 18683
rect 14280 18640 14332 18649
rect 14648 18683 14700 18692
rect 14648 18649 14657 18683
rect 14657 18649 14691 18683
rect 14691 18649 14700 18683
rect 14648 18640 14700 18649
rect 15752 18640 15804 18692
rect 20628 18708 20680 18760
rect 21180 18640 21232 18692
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 23112 18708 23164 18760
rect 23388 18751 23440 18760
rect 23388 18717 23397 18751
rect 23397 18717 23431 18751
rect 23431 18717 23440 18751
rect 23388 18708 23440 18717
rect 23756 18640 23808 18692
rect 15568 18615 15620 18624
rect 15568 18581 15577 18615
rect 15577 18581 15611 18615
rect 15611 18581 15620 18615
rect 15568 18572 15620 18581
rect 16580 18572 16632 18624
rect 18328 18572 18380 18624
rect 23020 18615 23072 18624
rect 23020 18581 23029 18615
rect 23029 18581 23063 18615
rect 23063 18581 23072 18615
rect 23020 18572 23072 18581
rect 25320 18572 25372 18624
rect 6884 18470 6936 18522
rect 6948 18470 7000 18522
rect 7012 18470 7064 18522
rect 7076 18470 7128 18522
rect 7140 18470 7192 18522
rect 12818 18470 12870 18522
rect 12882 18470 12934 18522
rect 12946 18470 12998 18522
rect 13010 18470 13062 18522
rect 13074 18470 13126 18522
rect 18752 18470 18804 18522
rect 18816 18470 18868 18522
rect 18880 18470 18932 18522
rect 18944 18470 18996 18522
rect 19008 18470 19060 18522
rect 24686 18470 24738 18522
rect 24750 18470 24802 18522
rect 24814 18470 24866 18522
rect 24878 18470 24930 18522
rect 24942 18470 24994 18522
rect 940 18368 992 18420
rect 5632 18368 5684 18420
rect 1216 18300 1268 18352
rect 4068 18300 4120 18352
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 1860 18232 1912 18284
rect 2320 18275 2372 18284
rect 2320 18241 2327 18275
rect 2327 18241 2361 18275
rect 2361 18241 2372 18275
rect 2320 18232 2372 18241
rect 4160 18232 4212 18284
rect 4712 18300 4764 18352
rect 4344 18232 4396 18284
rect 5632 18232 5684 18284
rect 8300 18368 8352 18420
rect 9128 18368 9180 18420
rect 11612 18368 11664 18420
rect 8024 18300 8076 18352
rect 8484 18275 8536 18284
rect 8484 18241 8491 18275
rect 8491 18241 8525 18275
rect 8525 18241 8536 18275
rect 8484 18232 8536 18241
rect 8944 18300 8996 18352
rect 12256 18300 12308 18352
rect 12624 18300 12676 18352
rect 14648 18368 14700 18420
rect 21364 18368 21416 18420
rect 23112 18300 23164 18352
rect 10324 18232 10376 18284
rect 12164 18232 12216 18284
rect 14096 18232 14148 18284
rect 1584 18164 1636 18216
rect 4988 18164 5040 18216
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 12532 18164 12584 18216
rect 12900 18164 12952 18216
rect 1492 18028 1544 18080
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 2964 18028 3016 18080
rect 4988 18071 5040 18080
rect 4988 18037 4997 18071
rect 4997 18037 5031 18071
rect 5031 18037 5040 18071
rect 4988 18028 5040 18037
rect 5540 18028 5592 18080
rect 6460 18028 6512 18080
rect 11152 18096 11204 18148
rect 13084 18096 13136 18148
rect 15752 18232 15804 18284
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 19248 18232 19300 18284
rect 22376 18232 22428 18284
rect 23296 18232 23348 18284
rect 17040 18164 17092 18216
rect 17408 18164 17460 18216
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 17684 18096 17736 18148
rect 17868 18096 17920 18148
rect 10508 18028 10560 18080
rect 10692 18028 10744 18080
rect 11704 18028 11756 18080
rect 13728 18028 13780 18080
rect 14556 18028 14608 18080
rect 16120 18028 16172 18080
rect 24400 18164 24452 18216
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 23572 18028 23624 18080
rect 24400 18071 24452 18080
rect 24400 18037 24409 18071
rect 24409 18037 24443 18071
rect 24443 18037 24452 18071
rect 24400 18028 24452 18037
rect 3917 17926 3969 17978
rect 3981 17926 4033 17978
rect 4045 17926 4097 17978
rect 4109 17926 4161 17978
rect 4173 17926 4225 17978
rect 9851 17926 9903 17978
rect 9915 17926 9967 17978
rect 9979 17926 10031 17978
rect 10043 17926 10095 17978
rect 10107 17926 10159 17978
rect 15785 17926 15837 17978
rect 15849 17926 15901 17978
rect 15913 17926 15965 17978
rect 15977 17926 16029 17978
rect 16041 17926 16093 17978
rect 21719 17926 21771 17978
rect 21783 17926 21835 17978
rect 21847 17926 21899 17978
rect 21911 17926 21963 17978
rect 21975 17926 22027 17978
rect 1860 17824 1912 17876
rect 2136 17824 2188 17876
rect 2688 17824 2740 17876
rect 4804 17824 4856 17876
rect 3792 17731 3844 17740
rect 3792 17697 3801 17731
rect 3801 17697 3835 17731
rect 3835 17697 3844 17731
rect 3792 17688 3844 17697
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 2136 17620 2188 17672
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 2780 17663 2832 17672
rect 2780 17629 2814 17663
rect 2814 17629 2832 17663
rect 2780 17620 2832 17629
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3608 17620 3660 17672
rect 3516 17552 3568 17604
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 3240 17484 3292 17536
rect 3424 17484 3476 17536
rect 4620 17484 4672 17536
rect 4804 17484 4856 17536
rect 5540 17484 5592 17536
rect 6368 17552 6420 17604
rect 6920 17620 6972 17672
rect 8392 17620 8444 17672
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 10784 17824 10836 17876
rect 11060 17824 11112 17876
rect 10508 17756 10560 17808
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 9312 17620 9364 17672
rect 11152 17688 11204 17740
rect 12256 17756 12308 17808
rect 10140 17620 10192 17672
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 12164 17688 12216 17740
rect 12716 17731 12768 17740
rect 12716 17697 12725 17731
rect 12725 17697 12759 17731
rect 12759 17697 12768 17731
rect 12716 17688 12768 17697
rect 12440 17620 12492 17672
rect 13084 17663 13136 17672
rect 13084 17629 13118 17663
rect 13118 17629 13136 17663
rect 13084 17620 13136 17629
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 13268 17620 13320 17629
rect 13912 17620 13964 17672
rect 17132 17731 17184 17740
rect 17132 17697 17141 17731
rect 17141 17697 17175 17731
rect 17175 17697 17184 17731
rect 17132 17688 17184 17697
rect 14832 17620 14884 17672
rect 15292 17620 15344 17672
rect 16304 17620 16356 17672
rect 17868 17824 17920 17876
rect 18052 17756 18104 17808
rect 22376 17824 22428 17876
rect 22836 17824 22888 17876
rect 23756 17867 23808 17876
rect 23756 17833 23765 17867
rect 23765 17833 23799 17867
rect 23799 17833 23808 17867
rect 23756 17824 23808 17833
rect 22192 17756 22244 17808
rect 12072 17484 12124 17536
rect 18052 17552 18104 17604
rect 17868 17484 17920 17536
rect 18972 17620 19024 17672
rect 22100 17688 22152 17740
rect 22468 17688 22520 17740
rect 22192 17663 22244 17672
rect 22192 17629 22201 17663
rect 22201 17629 22235 17663
rect 22235 17629 22244 17663
rect 22192 17620 22244 17629
rect 19432 17552 19484 17604
rect 20904 17552 20956 17604
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 22284 17527 22336 17536
rect 22284 17493 22293 17527
rect 22293 17493 22327 17527
rect 22327 17493 22336 17527
rect 22284 17484 22336 17493
rect 22468 17527 22520 17536
rect 22468 17493 22477 17527
rect 22477 17493 22511 17527
rect 22511 17493 22520 17527
rect 22468 17484 22520 17493
rect 22652 17484 22704 17536
rect 23112 17552 23164 17604
rect 24492 17484 24544 17536
rect 25044 17484 25096 17536
rect 6884 17382 6936 17434
rect 6948 17382 7000 17434
rect 7012 17382 7064 17434
rect 7076 17382 7128 17434
rect 7140 17382 7192 17434
rect 12818 17382 12870 17434
rect 12882 17382 12934 17434
rect 12946 17382 12998 17434
rect 13010 17382 13062 17434
rect 13074 17382 13126 17434
rect 18752 17382 18804 17434
rect 18816 17382 18868 17434
rect 18880 17382 18932 17434
rect 18944 17382 18996 17434
rect 19008 17382 19060 17434
rect 24686 17382 24738 17434
rect 24750 17382 24802 17434
rect 24814 17382 24866 17434
rect 24878 17382 24930 17434
rect 24942 17382 24994 17434
rect 388 17212 440 17264
rect 1032 17212 1084 17264
rect 3332 17280 3384 17332
rect 4528 17280 4580 17332
rect 6736 17280 6788 17332
rect 6920 17280 6972 17332
rect 3424 17212 3476 17264
rect 5172 17217 5224 17264
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 3792 17187 3844 17196
rect 3792 17153 3801 17187
rect 3801 17153 3835 17187
rect 3835 17153 3844 17187
rect 3792 17144 3844 17153
rect 4804 17144 4856 17196
rect 5172 17212 5197 17217
rect 5197 17212 5224 17217
rect 6644 17212 6696 17264
rect 9128 17280 9180 17332
rect 9772 17280 9824 17332
rect 10784 17280 10836 17332
rect 10968 17280 11020 17332
rect 8116 17212 8168 17264
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7196 17144 7248 17196
rect 7840 17144 7892 17196
rect 2044 17076 2096 17128
rect 2412 17076 2464 17128
rect 2596 17119 2648 17128
rect 2596 17085 2605 17119
rect 2605 17085 2639 17119
rect 2639 17085 2648 17119
rect 2596 17076 2648 17085
rect 4344 17076 4396 17128
rect 6184 17076 6236 17128
rect 2136 17008 2188 17060
rect 3700 17008 3752 17060
rect 7656 17076 7708 17128
rect 10600 17212 10652 17264
rect 12808 17280 12860 17332
rect 13268 17280 13320 17332
rect 14372 17280 14424 17332
rect 17040 17280 17092 17332
rect 17868 17280 17920 17332
rect 19432 17280 19484 17332
rect 9220 17144 9272 17196
rect 9588 17144 9640 17196
rect 10324 17187 10376 17196
rect 10324 17153 10331 17187
rect 10331 17153 10365 17187
rect 10365 17153 10376 17187
rect 10324 17144 10376 17153
rect 11060 17144 11112 17196
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 17132 17212 17184 17264
rect 11704 17076 11756 17128
rect 12072 17076 12124 17128
rect 12808 17144 12860 17196
rect 13452 17144 13504 17196
rect 15016 17144 15068 17196
rect 16304 17144 16356 17196
rect 14096 17076 14148 17128
rect 16856 17144 16908 17196
rect 17040 17144 17092 17196
rect 9588 17008 9640 17060
rect 2596 16940 2648 16992
rect 2688 16940 2740 16992
rect 6184 16940 6236 16992
rect 8392 16940 8444 16992
rect 11244 16940 11296 16992
rect 12532 16940 12584 16992
rect 14464 16983 14516 16992
rect 14464 16949 14473 16983
rect 14473 16949 14507 16983
rect 14507 16949 14516 16983
rect 14464 16940 14516 16949
rect 17684 17076 17736 17128
rect 20444 17280 20496 17332
rect 20628 17280 20680 17332
rect 20904 17280 20956 17332
rect 22192 17280 22244 17332
rect 22468 17280 22520 17332
rect 23020 17280 23072 17332
rect 25136 17280 25188 17332
rect 20536 17144 20588 17196
rect 20352 17076 20404 17128
rect 22836 17144 22888 17196
rect 23848 17187 23900 17196
rect 23848 17153 23857 17187
rect 23857 17153 23891 17187
rect 23891 17153 23900 17187
rect 23848 17144 23900 17153
rect 21824 17119 21876 17128
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 21640 17008 21692 17060
rect 16212 16983 16264 16992
rect 16212 16949 16221 16983
rect 16221 16949 16255 16983
rect 16255 16949 16264 16983
rect 16212 16940 16264 16949
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 18236 16940 18288 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 21548 16983 21600 16992
rect 21548 16949 21557 16983
rect 21557 16949 21591 16983
rect 21591 16949 21600 16983
rect 21548 16940 21600 16949
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 3917 16838 3969 16890
rect 3981 16838 4033 16890
rect 4045 16838 4097 16890
rect 4109 16838 4161 16890
rect 4173 16838 4225 16890
rect 9851 16838 9903 16890
rect 9915 16838 9967 16890
rect 9979 16838 10031 16890
rect 10043 16838 10095 16890
rect 10107 16838 10159 16890
rect 15785 16838 15837 16890
rect 15849 16838 15901 16890
rect 15913 16838 15965 16890
rect 15977 16838 16029 16890
rect 16041 16838 16093 16890
rect 21719 16838 21771 16890
rect 21783 16838 21835 16890
rect 21847 16838 21899 16890
rect 21911 16838 21963 16890
rect 21975 16838 22027 16890
rect 388 16736 440 16788
rect 3516 16736 3568 16788
rect 3792 16736 3844 16788
rect 9588 16736 9640 16788
rect 10324 16736 10376 16788
rect 11244 16736 11296 16788
rect 3240 16668 3292 16720
rect 6828 16668 6880 16720
rect 7564 16711 7616 16720
rect 7564 16677 7573 16711
rect 7573 16677 7607 16711
rect 7607 16677 7616 16711
rect 7564 16668 7616 16677
rect 1676 16600 1728 16652
rect 2228 16600 2280 16652
rect 3148 16600 3200 16652
rect 4528 16600 4580 16652
rect 5908 16600 5960 16652
rect 6368 16600 6420 16652
rect 6736 16600 6788 16652
rect 7012 16600 7064 16652
rect 7196 16600 7248 16652
rect 1584 16532 1636 16584
rect 3516 16532 3568 16584
rect 5356 16532 5408 16584
rect 6644 16532 6696 16584
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8668 16600 8720 16652
rect 11980 16600 12032 16652
rect 13360 16736 13412 16788
rect 16120 16736 16172 16788
rect 16212 16736 16264 16788
rect 16304 16736 16356 16788
rect 16764 16736 16816 16788
rect 16856 16736 16908 16788
rect 17316 16736 17368 16788
rect 17684 16736 17736 16788
rect 20168 16736 20220 16788
rect 21548 16736 21600 16788
rect 22284 16736 22336 16788
rect 15660 16600 15712 16652
rect 13636 16532 13688 16584
rect 14464 16532 14516 16584
rect 15568 16532 15620 16584
rect 16028 16600 16080 16652
rect 16764 16643 16816 16652
rect 16764 16609 16798 16643
rect 16798 16609 16816 16643
rect 16764 16600 16816 16609
rect 19616 16600 19668 16652
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 18236 16532 18288 16584
rect 2228 16464 2280 16516
rect 3056 16439 3108 16448
rect 3056 16405 3065 16439
rect 3065 16405 3099 16439
rect 3099 16405 3108 16439
rect 3056 16396 3108 16405
rect 4620 16464 4672 16516
rect 5264 16464 5316 16516
rect 13176 16464 13228 16516
rect 14004 16464 14056 16516
rect 14924 16464 14976 16516
rect 3976 16439 4028 16448
rect 3976 16405 3985 16439
rect 3985 16405 4019 16439
rect 4019 16405 4028 16439
rect 3976 16396 4028 16405
rect 4988 16396 5040 16448
rect 6276 16396 6328 16448
rect 8392 16396 8444 16448
rect 12256 16396 12308 16448
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 17408 16396 17460 16448
rect 17868 16439 17920 16448
rect 17868 16405 17877 16439
rect 17877 16405 17911 16439
rect 17911 16405 17920 16439
rect 17868 16396 17920 16405
rect 20720 16396 20772 16448
rect 21640 16532 21692 16584
rect 22928 16532 22980 16584
rect 23572 16532 23624 16584
rect 25228 16464 25280 16516
rect 23664 16396 23716 16448
rect 572 16328 624 16380
rect 6884 16294 6936 16346
rect 6948 16294 7000 16346
rect 7012 16294 7064 16346
rect 7076 16294 7128 16346
rect 7140 16294 7192 16346
rect 12818 16294 12870 16346
rect 12882 16294 12934 16346
rect 12946 16294 12998 16346
rect 13010 16294 13062 16346
rect 13074 16294 13126 16346
rect 18752 16294 18804 16346
rect 18816 16294 18868 16346
rect 18880 16294 18932 16346
rect 18944 16294 18996 16346
rect 19008 16294 19060 16346
rect 24686 16294 24738 16346
rect 24750 16294 24802 16346
rect 24814 16294 24866 16346
rect 24878 16294 24930 16346
rect 24942 16294 24994 16346
rect 572 16124 624 16176
rect 2044 16167 2096 16176
rect 2044 16133 2053 16167
rect 2053 16133 2087 16167
rect 2087 16133 2096 16167
rect 2044 16124 2096 16133
rect 1860 16056 1912 16108
rect 3332 16124 3384 16176
rect 5356 16167 5408 16176
rect 5356 16133 5365 16167
rect 5365 16133 5399 16167
rect 5399 16133 5408 16167
rect 5356 16124 5408 16133
rect 6276 16124 6328 16176
rect 8116 16192 8168 16244
rect 12716 16192 12768 16244
rect 14924 16192 14976 16244
rect 17868 16192 17920 16244
rect 18144 16167 18196 16176
rect 18144 16133 18178 16167
rect 18178 16133 18196 16167
rect 18144 16124 18196 16133
rect 20444 16192 20496 16244
rect 21456 16192 21508 16244
rect 21548 16192 21600 16244
rect 23296 16192 23348 16244
rect 23756 16192 23808 16244
rect 23848 16192 23900 16244
rect 2780 16056 2832 16108
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 9036 16056 9088 16108
rect 3608 15988 3660 16040
rect 4620 15988 4672 16040
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 4896 15988 4948 16040
rect 6276 15988 6328 16040
rect 7288 15988 7340 16040
rect 3516 15852 3568 15904
rect 8208 15920 8260 15972
rect 8668 15920 8720 15972
rect 9680 15988 9732 16040
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 12072 16099 12124 16108
rect 12072 16065 12081 16099
rect 12081 16065 12115 16099
rect 12115 16065 12124 16099
rect 12072 16056 12124 16065
rect 12256 16056 12308 16108
rect 13636 16056 13688 16108
rect 14280 16056 14332 16108
rect 15016 16056 15068 16108
rect 19340 16099 19392 16108
rect 19340 16065 19349 16099
rect 19349 16065 19383 16099
rect 19383 16065 19392 16099
rect 19340 16056 19392 16065
rect 20720 16056 20772 16108
rect 21272 16124 21324 16176
rect 13360 15988 13412 16040
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 13912 15920 13964 15972
rect 9680 15852 9732 15904
rect 10324 15852 10376 15904
rect 10508 15852 10560 15904
rect 14280 15852 14332 15904
rect 15752 15852 15804 15904
rect 16856 15852 16908 15904
rect 20168 15920 20220 15972
rect 19524 15852 19576 15904
rect 19984 15852 20036 15904
rect 22100 15852 22152 15904
rect 24400 16056 24452 16108
rect 23480 15988 23532 16040
rect 23572 15852 23624 15904
rect 23848 15852 23900 15904
rect 3917 15750 3969 15802
rect 3981 15750 4033 15802
rect 4045 15750 4097 15802
rect 4109 15750 4161 15802
rect 4173 15750 4225 15802
rect 9851 15750 9903 15802
rect 9915 15750 9967 15802
rect 9979 15750 10031 15802
rect 10043 15750 10095 15802
rect 10107 15750 10159 15802
rect 15785 15750 15837 15802
rect 15849 15750 15901 15802
rect 15913 15750 15965 15802
rect 15977 15750 16029 15802
rect 16041 15750 16093 15802
rect 21719 15750 21771 15802
rect 21783 15750 21835 15802
rect 21847 15750 21899 15802
rect 21911 15750 21963 15802
rect 21975 15750 22027 15802
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 2136 15648 2188 15700
rect 2780 15648 2832 15700
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 1584 15580 1636 15632
rect 3700 15580 3752 15632
rect 4712 15648 4764 15700
rect 1860 15512 1912 15564
rect 1952 15444 2004 15496
rect 2412 15444 2464 15496
rect 3700 15444 3752 15496
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 7288 15648 7340 15700
rect 7564 15648 7616 15700
rect 9680 15648 9732 15700
rect 10600 15648 10652 15700
rect 12440 15648 12492 15700
rect 16856 15648 16908 15700
rect 19340 15648 19392 15700
rect 8208 15580 8260 15632
rect 9220 15580 9272 15632
rect 4068 15487 4120 15496
rect 4068 15453 4075 15487
rect 4075 15453 4109 15487
rect 4109 15453 4120 15487
rect 4068 15444 4120 15453
rect 4160 15444 4212 15496
rect 5264 15444 5316 15496
rect 6276 15444 6328 15496
rect 9680 15512 9732 15564
rect 9956 15555 10008 15564
rect 9956 15521 9990 15555
rect 9990 15521 10008 15555
rect 9956 15512 10008 15521
rect 10324 15512 10376 15564
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 7288 15308 7340 15360
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 9036 15308 9088 15360
rect 9312 15308 9364 15360
rect 9680 15308 9732 15360
rect 12072 15512 12124 15564
rect 18328 15512 18380 15564
rect 19156 15512 19208 15564
rect 20812 15512 20864 15564
rect 22376 15555 22428 15564
rect 22376 15521 22385 15555
rect 22385 15521 22419 15555
rect 22419 15521 22428 15555
rect 22376 15512 22428 15521
rect 11152 15487 11204 15496
rect 11152 15453 11159 15487
rect 11159 15453 11193 15487
rect 11193 15453 11204 15487
rect 11152 15444 11204 15453
rect 11244 15376 11296 15428
rect 15016 15444 15068 15496
rect 17224 15444 17276 15496
rect 17684 15444 17736 15496
rect 18144 15444 18196 15496
rect 13268 15376 13320 15428
rect 14464 15376 14516 15428
rect 17132 15376 17184 15428
rect 17776 15376 17828 15428
rect 19340 15376 19392 15428
rect 19616 15444 19668 15496
rect 21732 15444 21784 15496
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 24124 15691 24176 15700
rect 24124 15657 24133 15691
rect 24133 15657 24167 15691
rect 24167 15657 24176 15691
rect 24124 15648 24176 15657
rect 22284 15444 22336 15453
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 11980 15308 12032 15360
rect 14280 15308 14332 15360
rect 17224 15308 17276 15360
rect 17868 15308 17920 15360
rect 18144 15308 18196 15360
rect 19800 15308 19852 15360
rect 20444 15308 20496 15360
rect 20996 15308 21048 15360
rect 22100 15351 22152 15360
rect 22100 15317 22109 15351
rect 22109 15317 22143 15351
rect 22143 15317 22152 15351
rect 22100 15308 22152 15317
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 6884 15206 6936 15258
rect 6948 15206 7000 15258
rect 7012 15206 7064 15258
rect 7076 15206 7128 15258
rect 7140 15206 7192 15258
rect 12818 15206 12870 15258
rect 12882 15206 12934 15258
rect 12946 15206 12998 15258
rect 13010 15206 13062 15258
rect 13074 15206 13126 15258
rect 18752 15206 18804 15258
rect 18816 15206 18868 15258
rect 18880 15206 18932 15258
rect 18944 15206 18996 15258
rect 19008 15206 19060 15258
rect 24686 15206 24738 15258
rect 24750 15206 24802 15258
rect 24814 15206 24866 15258
rect 24878 15206 24930 15258
rect 24942 15206 24994 15258
rect 1308 15104 1360 15156
rect 2228 15104 2280 15156
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 2320 14764 2372 14816
rect 3056 15104 3108 15156
rect 3976 15147 4028 15156
rect 3976 15113 3985 15147
rect 3985 15113 4019 15147
rect 4019 15113 4028 15147
rect 3976 15104 4028 15113
rect 4160 15104 4212 15156
rect 3240 15036 3292 15088
rect 6460 15104 6512 15156
rect 4344 15036 4396 15088
rect 3792 14968 3844 15020
rect 4252 14968 4304 15020
rect 5264 15036 5316 15088
rect 4988 14968 5040 15020
rect 7380 15104 7432 15156
rect 9404 15104 9456 15156
rect 10140 15104 10192 15156
rect 11612 15104 11664 15156
rect 11796 15104 11848 15156
rect 12624 15104 12676 15156
rect 13452 15104 13504 15156
rect 16948 15104 17000 15156
rect 7472 14968 7524 15020
rect 9220 15011 9272 15020
rect 9220 14977 9229 15011
rect 9229 14977 9263 15011
rect 9263 14977 9272 15011
rect 9220 14968 9272 14977
rect 11152 15036 11204 15088
rect 11796 14968 11848 15020
rect 11980 15011 12032 15020
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14968 12032 14977
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 13452 14968 13504 15020
rect 20812 15104 20864 15156
rect 22100 15104 22152 15156
rect 22744 15104 22796 15156
rect 23572 15104 23624 15156
rect 18144 15036 18196 15088
rect 19616 15036 19668 15088
rect 15292 14968 15344 15020
rect 17224 14968 17276 15020
rect 17408 15011 17460 15020
rect 17408 14977 17442 15011
rect 17442 14977 17460 15011
rect 17408 14968 17460 14977
rect 17868 14968 17920 15020
rect 19340 14968 19392 15020
rect 2780 14832 2832 14884
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 3240 14764 3292 14816
rect 6644 14900 6696 14952
rect 4712 14764 4764 14816
rect 4804 14764 4856 14816
rect 6460 14832 6512 14884
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 11888 14900 11940 14952
rect 12808 14900 12860 14952
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 20352 15036 20404 15088
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 5448 14764 5500 14816
rect 5908 14764 5960 14816
rect 6828 14764 6880 14816
rect 7288 14764 7340 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 14004 14764 14056 14816
rect 22192 14968 22244 15020
rect 22468 14968 22520 15020
rect 14648 14832 14700 14884
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 16212 14832 16264 14884
rect 16672 14832 16724 14884
rect 21732 14900 21784 14952
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 18696 14764 18748 14816
rect 19892 14764 19944 14816
rect 21640 14807 21692 14816
rect 21640 14773 21649 14807
rect 21649 14773 21683 14807
rect 21683 14773 21692 14807
rect 21640 14764 21692 14773
rect 24308 15036 24360 15088
rect 23020 14900 23072 14952
rect 22284 14764 22336 14816
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 3917 14662 3969 14714
rect 3981 14662 4033 14714
rect 4045 14662 4097 14714
rect 4109 14662 4161 14714
rect 4173 14662 4225 14714
rect 9851 14662 9903 14714
rect 9915 14662 9967 14714
rect 9979 14662 10031 14714
rect 10043 14662 10095 14714
rect 10107 14662 10159 14714
rect 15785 14662 15837 14714
rect 15849 14662 15901 14714
rect 15913 14662 15965 14714
rect 15977 14662 16029 14714
rect 16041 14662 16093 14714
rect 21719 14662 21771 14714
rect 21783 14662 21835 14714
rect 21847 14662 21899 14714
rect 21911 14662 21963 14714
rect 21975 14662 22027 14714
rect 2872 14560 2924 14612
rect 3792 14560 3844 14612
rect 2872 14424 2924 14476
rect 4344 14492 4396 14544
rect 5356 14492 5408 14544
rect 7564 14560 7616 14612
rect 8208 14560 8260 14612
rect 8852 14560 8904 14612
rect 11152 14560 11204 14612
rect 10140 14492 10192 14544
rect 10508 14492 10560 14544
rect 940 14356 992 14408
rect 1860 14356 1912 14408
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 6460 14424 6512 14476
rect 6828 14467 6880 14476
rect 6828 14433 6837 14467
rect 6837 14433 6871 14467
rect 6871 14433 6880 14467
rect 6828 14424 6880 14433
rect 8116 14424 8168 14476
rect 10416 14424 10468 14476
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 4804 14356 4856 14408
rect 4988 14356 5040 14408
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 6736 14356 6788 14408
rect 7656 14356 7708 14408
rect 8024 14356 8076 14408
rect 9404 14356 9456 14408
rect 10048 14356 10100 14408
rect 2504 14220 2556 14272
rect 3516 14220 3568 14272
rect 4804 14220 4856 14272
rect 7380 14288 7432 14340
rect 11244 14467 11296 14476
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 6920 14220 6972 14272
rect 11060 14220 11112 14272
rect 11152 14220 11204 14272
rect 11428 14356 11480 14408
rect 12072 14560 12124 14612
rect 13636 14560 13688 14612
rect 14648 14560 14700 14612
rect 14924 14560 14976 14612
rect 15292 14560 15344 14612
rect 18512 14560 18564 14612
rect 20812 14560 20864 14612
rect 23296 14560 23348 14612
rect 13452 14492 13504 14544
rect 15016 14424 15068 14476
rect 16212 14492 16264 14544
rect 16028 14424 16080 14476
rect 16488 14424 16540 14476
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 17224 14467 17276 14476
rect 17224 14433 17258 14467
rect 17258 14433 17276 14467
rect 17224 14424 17276 14433
rect 12072 14356 12124 14408
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 12900 14399 12952 14408
rect 12900 14365 12907 14399
rect 12907 14365 12941 14399
rect 12941 14365 12952 14399
rect 12900 14356 12952 14365
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 13176 14220 13228 14272
rect 17500 14220 17552 14272
rect 21640 14424 21692 14476
rect 20352 14356 20404 14408
rect 22192 14356 22244 14408
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 19156 14220 19208 14272
rect 22100 14263 22152 14272
rect 22100 14229 22109 14263
rect 22109 14229 22143 14263
rect 22143 14229 22152 14263
rect 22100 14220 22152 14229
rect 25136 14492 25188 14544
rect 23756 14424 23808 14476
rect 24216 14356 24268 14408
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 25320 14220 25372 14272
rect 6884 14118 6936 14170
rect 6948 14118 7000 14170
rect 7012 14118 7064 14170
rect 7076 14118 7128 14170
rect 7140 14118 7192 14170
rect 12818 14118 12870 14170
rect 12882 14118 12934 14170
rect 12946 14118 12998 14170
rect 13010 14118 13062 14170
rect 13074 14118 13126 14170
rect 18752 14118 18804 14170
rect 18816 14118 18868 14170
rect 18880 14118 18932 14170
rect 18944 14118 18996 14170
rect 19008 14118 19060 14170
rect 24686 14118 24738 14170
rect 24750 14118 24802 14170
rect 24814 14118 24866 14170
rect 24878 14118 24930 14170
rect 24942 14118 24994 14170
rect 25320 14084 25372 14136
rect 25872 14084 25924 14136
rect 2964 14016 3016 14068
rect 3332 14016 3384 14068
rect 1584 13948 1636 14000
rect 4804 14016 4856 14068
rect 6092 14016 6144 14068
rect 6736 14016 6788 14068
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 1492 13812 1544 13864
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 4712 13880 4764 13932
rect 5080 13880 5132 13932
rect 5908 13880 5960 13932
rect 6460 13880 6512 13932
rect 7656 14016 7708 14068
rect 7840 14016 7892 14068
rect 9772 14016 9824 14068
rect 10048 14016 10100 14068
rect 10324 14016 10376 14068
rect 7012 13948 7064 14000
rect 8024 13948 8076 14000
rect 9680 13948 9732 14000
rect 9864 13953 9916 14000
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 2320 13676 2372 13728
rect 3332 13676 3384 13728
rect 4436 13719 4488 13728
rect 4436 13685 4445 13719
rect 4445 13685 4479 13719
rect 4479 13685 4488 13719
rect 4436 13676 4488 13685
rect 8024 13744 8076 13796
rect 7840 13719 7892 13728
rect 7840 13685 7849 13719
rect 7849 13685 7883 13719
rect 7883 13685 7892 13719
rect 7840 13676 7892 13685
rect 9404 13880 9456 13932
rect 9864 13948 9889 13953
rect 9889 13948 9916 13953
rect 15476 14016 15528 14068
rect 17408 14016 17460 14068
rect 18052 14016 18104 14068
rect 19156 14016 19208 14068
rect 19616 14016 19668 14068
rect 21180 14016 21232 14068
rect 14464 13948 14516 14000
rect 16672 13948 16724 14000
rect 9496 13744 9548 13796
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 13636 13923 13688 13932
rect 13636 13889 13645 13923
rect 13645 13889 13679 13923
rect 13679 13889 13688 13923
rect 13636 13880 13688 13889
rect 14280 13880 14332 13932
rect 16948 13923 17000 13932
rect 16948 13889 16955 13923
rect 16955 13889 16989 13923
rect 16989 13889 17000 13923
rect 16948 13880 17000 13889
rect 17408 13880 17460 13932
rect 19064 13880 19116 13932
rect 19984 13948 20036 14000
rect 21640 13948 21692 14000
rect 23112 14016 23164 14068
rect 23296 14016 23348 14068
rect 25780 14016 25832 14068
rect 21548 13880 21600 13932
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 22744 13880 22796 13889
rect 12992 13812 13044 13864
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 13176 13812 13228 13864
rect 13544 13812 13596 13864
rect 14004 13812 14056 13864
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 11888 13676 11940 13728
rect 14924 13676 14976 13728
rect 15476 13676 15528 13728
rect 16028 13676 16080 13728
rect 16764 13676 16816 13728
rect 18328 13676 18380 13728
rect 19156 13744 19208 13796
rect 19984 13812 20036 13864
rect 23204 13923 23256 13932
rect 23204 13889 23213 13923
rect 23213 13889 23247 13923
rect 23247 13889 23256 13923
rect 23204 13880 23256 13889
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 23480 13880 23532 13889
rect 23572 13855 23624 13864
rect 19064 13719 19116 13728
rect 19064 13685 19073 13719
rect 19073 13685 19107 13719
rect 19107 13685 19116 13719
rect 19064 13676 19116 13685
rect 19524 13719 19576 13728
rect 19524 13685 19533 13719
rect 19533 13685 19567 13719
rect 19567 13685 19576 13719
rect 19524 13676 19576 13685
rect 22192 13744 22244 13796
rect 23572 13821 23581 13855
rect 23581 13821 23615 13855
rect 23615 13821 23624 13855
rect 23572 13812 23624 13821
rect 25780 13812 25832 13864
rect 23020 13744 23072 13796
rect 22100 13676 22152 13728
rect 23296 13676 23348 13728
rect 24400 13719 24452 13728
rect 24400 13685 24409 13719
rect 24409 13685 24443 13719
rect 24443 13685 24452 13719
rect 24400 13676 24452 13685
rect 3917 13574 3969 13626
rect 3981 13574 4033 13626
rect 4045 13574 4097 13626
rect 4109 13574 4161 13626
rect 4173 13574 4225 13626
rect 9851 13574 9903 13626
rect 9915 13574 9967 13626
rect 9979 13574 10031 13626
rect 10043 13574 10095 13626
rect 10107 13574 10159 13626
rect 15785 13574 15837 13626
rect 15849 13574 15901 13626
rect 15913 13574 15965 13626
rect 15977 13574 16029 13626
rect 16041 13574 16093 13626
rect 21719 13574 21771 13626
rect 21783 13574 21835 13626
rect 21847 13574 21899 13626
rect 21911 13574 21963 13626
rect 21975 13574 22027 13626
rect 1216 13472 1268 13524
rect 1308 13404 1360 13456
rect 1400 13336 1452 13388
rect 2136 13336 2188 13388
rect 5080 13404 5132 13456
rect 5724 13404 5776 13456
rect 5908 13404 5960 13456
rect 8392 13404 8444 13456
rect 9496 13404 9548 13456
rect 9864 13404 9916 13456
rect 10232 13404 10284 13456
rect 10324 13404 10376 13456
rect 1492 13311 1544 13320
rect 1492 13277 1501 13311
rect 1501 13277 1535 13311
rect 1535 13277 1544 13311
rect 1492 13268 1544 13277
rect 3332 13268 3384 13320
rect 2596 13243 2648 13252
rect 2596 13209 2605 13243
rect 2605 13209 2639 13243
rect 2639 13209 2648 13243
rect 2596 13200 2648 13209
rect 3148 13243 3200 13252
rect 3148 13209 3157 13243
rect 3157 13209 3191 13243
rect 3191 13209 3200 13243
rect 3148 13200 3200 13209
rect 3976 13268 4028 13320
rect 6092 13336 6144 13388
rect 9128 13336 9180 13388
rect 10140 13336 10192 13388
rect 13452 13472 13504 13524
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 13636 13336 13688 13388
rect 13912 13336 13964 13388
rect 16856 13472 16908 13524
rect 18512 13472 18564 13524
rect 20812 13472 20864 13524
rect 22560 13472 22612 13524
rect 23480 13472 23532 13524
rect 17132 13336 17184 13388
rect 17684 13336 17736 13388
rect 19524 13336 19576 13388
rect 5540 13268 5592 13320
rect 5908 13268 5960 13320
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 8024 13200 8076 13252
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 11888 13268 11940 13320
rect 11980 13268 12032 13320
rect 12256 13268 12308 13320
rect 9956 13200 10008 13252
rect 14372 13268 14424 13320
rect 14648 13268 14700 13320
rect 15292 13268 15344 13320
rect 16764 13268 16816 13320
rect 2780 13132 2832 13184
rect 4436 13132 4488 13184
rect 5356 13132 5408 13184
rect 6276 13132 6328 13184
rect 7288 13132 7340 13184
rect 17684 13200 17736 13252
rect 18236 13200 18288 13252
rect 19064 13268 19116 13320
rect 19524 13200 19576 13252
rect 13176 13132 13228 13184
rect 14740 13132 14792 13184
rect 18052 13132 18104 13184
rect 19984 13404 20036 13456
rect 21272 13404 21324 13456
rect 22376 13404 22428 13456
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 20536 13268 20588 13320
rect 21548 13268 21600 13320
rect 20168 13243 20220 13252
rect 20168 13209 20177 13243
rect 20177 13209 20211 13243
rect 20211 13209 20220 13243
rect 20168 13200 20220 13209
rect 19984 13132 20036 13184
rect 22560 13311 22612 13320
rect 22560 13277 22569 13311
rect 22569 13277 22603 13311
rect 22603 13277 22612 13311
rect 22560 13268 22612 13277
rect 23480 13200 23532 13252
rect 6884 13030 6936 13082
rect 6948 13030 7000 13082
rect 7012 13030 7064 13082
rect 7076 13030 7128 13082
rect 7140 13030 7192 13082
rect 12818 13030 12870 13082
rect 12882 13030 12934 13082
rect 12946 13030 12998 13082
rect 13010 13030 13062 13082
rect 13074 13030 13126 13082
rect 18752 13030 18804 13082
rect 18816 13030 18868 13082
rect 18880 13030 18932 13082
rect 18944 13030 18996 13082
rect 19008 13030 19060 13082
rect 24686 13030 24738 13082
rect 24750 13030 24802 13082
rect 24814 13030 24866 13082
rect 24878 13030 24930 13082
rect 24942 13030 24994 13082
rect 1768 12971 1820 12980
rect 1768 12937 1777 12971
rect 1777 12937 1811 12971
rect 1811 12937 1820 12971
rect 1768 12928 1820 12937
rect 6368 12928 6420 12980
rect 2228 12792 2280 12844
rect 3240 12792 3292 12844
rect 3608 12792 3660 12844
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 6092 12792 6144 12844
rect 7288 12928 7340 12980
rect 7380 12928 7432 12980
rect 7932 12928 7984 12980
rect 6736 12792 6788 12844
rect 9128 12928 9180 12980
rect 9496 12928 9548 12980
rect 10968 12928 11020 12980
rect 11612 12928 11664 12980
rect 20168 12928 20220 12980
rect 10508 12860 10560 12912
rect 1768 12724 1820 12776
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 3792 12724 3844 12776
rect 4436 12724 4488 12776
rect 4620 12767 4672 12776
rect 4620 12733 4647 12767
rect 4647 12733 4672 12767
rect 4620 12724 4672 12733
rect 4737 12767 4789 12776
rect 4737 12733 4746 12767
rect 4746 12733 4780 12767
rect 4780 12733 4789 12767
rect 4737 12724 4789 12733
rect 3240 12656 3292 12708
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 3792 12588 3844 12640
rect 6092 12588 6144 12640
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 9864 12792 9916 12844
rect 19156 12860 19208 12912
rect 7840 12724 7892 12776
rect 8024 12767 8076 12776
rect 8024 12733 8033 12767
rect 8033 12733 8067 12767
rect 8067 12733 8076 12767
rect 8024 12724 8076 12733
rect 8392 12724 8444 12776
rect 9036 12767 9088 12776
rect 9036 12733 9070 12767
rect 9070 12733 9088 12767
rect 9036 12724 9088 12733
rect 11336 12792 11388 12844
rect 11980 12835 12032 12844
rect 11980 12801 11987 12835
rect 11987 12801 12021 12835
rect 12021 12801 12032 12835
rect 11980 12792 12032 12801
rect 12072 12792 12124 12844
rect 14832 12792 14884 12844
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17092 12835
rect 17040 12792 17092 12801
rect 17684 12792 17736 12844
rect 11244 12656 11296 12708
rect 11612 12656 11664 12708
rect 11980 12588 12032 12640
rect 12072 12588 12124 12640
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 16120 12724 16172 12776
rect 19984 12860 20036 12912
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 20536 12860 20588 12912
rect 22468 12928 22520 12980
rect 22836 12928 22888 12980
rect 23572 12928 23624 12980
rect 20996 12724 21048 12776
rect 22192 12792 22244 12844
rect 22468 12802 22520 12854
rect 24492 12860 24544 12912
rect 21548 12656 21600 12708
rect 14648 12588 14700 12640
rect 17776 12631 17828 12640
rect 17776 12597 17785 12631
rect 17785 12597 17819 12631
rect 17819 12597 17828 12631
rect 17776 12588 17828 12597
rect 18328 12588 18380 12640
rect 20352 12588 20404 12640
rect 21180 12588 21232 12640
rect 22100 12588 22152 12640
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 3917 12486 3969 12538
rect 3981 12486 4033 12538
rect 4045 12486 4097 12538
rect 4109 12486 4161 12538
rect 4173 12486 4225 12538
rect 9851 12486 9903 12538
rect 9915 12486 9967 12538
rect 9979 12486 10031 12538
rect 10043 12486 10095 12538
rect 10107 12486 10159 12538
rect 15785 12486 15837 12538
rect 15849 12486 15901 12538
rect 15913 12486 15965 12538
rect 15977 12486 16029 12538
rect 16041 12486 16093 12538
rect 21719 12486 21771 12538
rect 21783 12486 21835 12538
rect 21847 12486 21899 12538
rect 21911 12486 21963 12538
rect 21975 12486 22027 12538
rect 3608 12384 3660 12436
rect 4252 12384 4304 12436
rect 4712 12384 4764 12436
rect 5356 12384 5408 12436
rect 4436 12316 4488 12368
rect 940 12248 992 12300
rect 2044 12248 2096 12300
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 2780 12248 2832 12300
rect 3332 12248 3384 12300
rect 4252 12248 4304 12300
rect 2688 12223 2740 12232
rect 2688 12189 2697 12223
rect 2697 12189 2731 12223
rect 2731 12189 2740 12223
rect 2688 12180 2740 12189
rect 3700 12180 3752 12232
rect 4160 12180 4212 12232
rect 1952 12044 2004 12096
rect 4804 12180 4856 12232
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 6920 12384 6972 12436
rect 7380 12384 7432 12436
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 7932 12384 7984 12436
rect 15476 12384 15528 12436
rect 8484 12316 8536 12368
rect 12532 12248 12584 12300
rect 13912 12248 13964 12300
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 17592 12291 17644 12300
rect 17592 12257 17601 12291
rect 17601 12257 17635 12291
rect 17635 12257 17644 12291
rect 17592 12248 17644 12257
rect 18328 12248 18380 12300
rect 18604 12248 18656 12300
rect 20996 12384 21048 12436
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 4988 12180 5040 12232
rect 6092 12223 6144 12232
rect 6092 12189 6101 12223
rect 6101 12189 6135 12223
rect 6135 12189 6144 12223
rect 6092 12180 6144 12189
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 12716 12180 12768 12232
rect 12808 12180 12860 12232
rect 14372 12180 14424 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 14740 12180 14792 12232
rect 15384 12180 15436 12232
rect 15476 12180 15528 12232
rect 16488 12180 16540 12232
rect 16764 12180 16816 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20220 12223
rect 20168 12180 20220 12189
rect 20536 12180 20588 12232
rect 20812 12180 20864 12232
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 25136 12384 25188 12436
rect 25228 12316 25280 12368
rect 23848 12248 23900 12300
rect 3792 12044 3844 12096
rect 6092 12044 6144 12096
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 9036 12112 9088 12164
rect 9680 12044 9732 12096
rect 11244 12044 11296 12096
rect 11612 12044 11664 12096
rect 11980 12112 12032 12164
rect 12164 12112 12216 12164
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 14188 12112 14240 12164
rect 13176 12044 13228 12096
rect 13728 12044 13780 12096
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 14372 12044 14424 12096
rect 14648 12044 14700 12096
rect 15108 12044 15160 12096
rect 21548 12155 21600 12164
rect 15752 12044 15804 12096
rect 21548 12121 21582 12155
rect 21582 12121 21600 12155
rect 21548 12112 21600 12121
rect 23664 12180 23716 12232
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 20720 12044 20772 12096
rect 21824 12044 21876 12096
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 23112 12087 23164 12096
rect 23112 12053 23121 12087
rect 23121 12053 23155 12087
rect 23155 12053 23164 12087
rect 23112 12044 23164 12053
rect 6884 11942 6936 11994
rect 6948 11942 7000 11994
rect 7012 11942 7064 11994
rect 7076 11942 7128 11994
rect 7140 11942 7192 11994
rect 12818 11942 12870 11994
rect 12882 11942 12934 11994
rect 12946 11942 12998 11994
rect 13010 11942 13062 11994
rect 13074 11942 13126 11994
rect 18752 11942 18804 11994
rect 18816 11942 18868 11994
rect 18880 11942 18932 11994
rect 18944 11942 18996 11994
rect 19008 11942 19060 11994
rect 24686 11942 24738 11994
rect 24750 11942 24802 11994
rect 24814 11942 24866 11994
rect 24878 11942 24930 11994
rect 24942 11942 24994 11994
rect 2412 11840 2464 11892
rect 2044 11772 2096 11824
rect 4160 11840 4212 11892
rect 4896 11840 4948 11892
rect 5540 11840 5592 11892
rect 6368 11840 6420 11892
rect 3056 11772 3108 11824
rect 1768 11636 1820 11688
rect 1492 11500 1544 11552
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 3976 11772 4028 11824
rect 4896 11679 4948 11688
rect 4896 11645 4905 11679
rect 4905 11645 4939 11679
rect 4939 11645 4948 11679
rect 4896 11636 4948 11645
rect 4436 11500 4488 11552
rect 8024 11840 8076 11892
rect 12164 11840 12216 11892
rect 12440 11840 12492 11892
rect 12532 11883 12584 11892
rect 12532 11849 12541 11883
rect 12541 11849 12575 11883
rect 12575 11849 12584 11883
rect 12532 11840 12584 11849
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 15384 11840 15436 11892
rect 17040 11840 17092 11892
rect 17868 11772 17920 11824
rect 7288 11704 7340 11756
rect 8576 11747 8628 11756
rect 8576 11713 8583 11747
rect 8583 11713 8617 11747
rect 8617 11713 8628 11747
rect 8576 11704 8628 11713
rect 9036 11704 9088 11756
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 12808 11704 12860 11756
rect 13176 11747 13228 11756
rect 13176 11713 13183 11747
rect 13183 11713 13217 11747
rect 13217 11713 13228 11747
rect 13176 11704 13228 11713
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 15200 11747 15252 11756
rect 15200 11713 15207 11747
rect 15207 11713 15241 11747
rect 15241 11713 15252 11747
rect 15200 11704 15252 11713
rect 15292 11704 15344 11756
rect 16304 11704 16356 11756
rect 22744 11840 22796 11892
rect 22836 11840 22888 11892
rect 23112 11840 23164 11892
rect 18328 11777 18380 11824
rect 18328 11772 18353 11777
rect 18353 11772 18380 11777
rect 18604 11772 18656 11824
rect 21824 11772 21876 11824
rect 20352 11704 20404 11756
rect 21548 11704 21600 11756
rect 23480 11704 23532 11756
rect 23572 11747 23624 11756
rect 23572 11713 23581 11747
rect 23581 11713 23615 11747
rect 23615 11713 23624 11747
rect 23572 11704 23624 11713
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 11060 11568 11112 11620
rect 11428 11568 11480 11620
rect 7012 11500 7064 11552
rect 8208 11500 8260 11552
rect 9128 11500 9180 11552
rect 9312 11543 9364 11552
rect 9312 11509 9321 11543
rect 9321 11509 9355 11543
rect 9355 11509 9364 11543
rect 9312 11500 9364 11509
rect 11888 11500 11940 11552
rect 13728 11636 13780 11688
rect 12992 11500 13044 11552
rect 13912 11500 13964 11552
rect 15752 11636 15804 11688
rect 15844 11636 15896 11688
rect 16120 11636 16172 11688
rect 22928 11636 22980 11688
rect 19156 11568 19208 11620
rect 25044 11704 25096 11756
rect 25320 11704 25372 11756
rect 16948 11500 17000 11552
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19064 11500 19116 11509
rect 22560 11500 22612 11552
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 25228 11500 25280 11552
rect 3917 11398 3969 11450
rect 3981 11398 4033 11450
rect 4045 11398 4097 11450
rect 4109 11398 4161 11450
rect 4173 11398 4225 11450
rect 9851 11398 9903 11450
rect 9915 11398 9967 11450
rect 9979 11398 10031 11450
rect 10043 11398 10095 11450
rect 10107 11398 10159 11450
rect 15785 11398 15837 11450
rect 15849 11398 15901 11450
rect 15913 11398 15965 11450
rect 15977 11398 16029 11450
rect 16041 11398 16093 11450
rect 21719 11398 21771 11450
rect 21783 11398 21835 11450
rect 21847 11398 21899 11450
rect 21911 11398 21963 11450
rect 21975 11398 22027 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 3056 11296 3108 11348
rect 3884 11296 3936 11348
rect 1676 11271 1728 11280
rect 1676 11237 1685 11271
rect 1685 11237 1719 11271
rect 1719 11237 1728 11271
rect 1676 11228 1728 11237
rect 1860 11228 1912 11280
rect 3240 11228 3292 11280
rect 6736 11296 6788 11348
rect 7472 11296 7524 11348
rect 9312 11296 9364 11348
rect 9680 11296 9732 11348
rect 9864 11296 9916 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 2504 11092 2556 11144
rect 3792 11160 3844 11212
rect 3976 11160 4028 11212
rect 4528 11160 4580 11212
rect 3332 11092 3384 11144
rect 4344 11092 4396 11144
rect 7748 11160 7800 11212
rect 13820 11296 13872 11348
rect 15384 11296 15436 11348
rect 16764 11296 16816 11348
rect 17040 11271 17092 11280
rect 17040 11237 17049 11271
rect 17049 11237 17083 11271
rect 17083 11237 17092 11271
rect 17040 11228 17092 11237
rect 16212 11203 16264 11212
rect 16212 11169 16246 11203
rect 16246 11169 16264 11203
rect 16212 11160 16264 11169
rect 18236 11296 18288 11348
rect 18604 11296 18656 11348
rect 19064 11296 19116 11348
rect 23480 11296 23532 11348
rect 17868 11228 17920 11280
rect 20720 11271 20772 11280
rect 20720 11237 20729 11271
rect 20729 11237 20763 11271
rect 20763 11237 20772 11271
rect 20720 11228 20772 11237
rect 22284 11228 22336 11280
rect 2044 11067 2096 11076
rect 2044 11033 2053 11067
rect 2053 11033 2087 11067
rect 2087 11033 2096 11067
rect 2044 11024 2096 11033
rect 2596 11024 2648 11076
rect 940 10956 992 11008
rect 3332 10956 3384 11008
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 4436 11067 4488 11076
rect 4436 11033 4445 11067
rect 4445 11033 4479 11067
rect 4479 11033 4488 11067
rect 4436 11024 4488 11033
rect 7380 11092 7432 11144
rect 7012 11024 7064 11076
rect 7932 11092 7984 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 9956 11135 10008 11144
rect 9956 11101 9990 11135
rect 9990 11101 10008 11135
rect 9956 11092 10008 11101
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 12716 11092 12768 11144
rect 13176 11092 13228 11144
rect 7748 11024 7800 11076
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 17408 11135 17460 11144
rect 17408 11101 17415 11135
rect 17415 11101 17449 11135
rect 17449 11101 17460 11135
rect 17408 11092 17460 11101
rect 18604 11092 18656 11144
rect 19524 11160 19576 11212
rect 22376 11160 22428 11212
rect 22744 11203 22796 11212
rect 22744 11169 22753 11203
rect 22753 11169 22787 11203
rect 22787 11169 22796 11203
rect 22744 11160 22796 11169
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 21180 11092 21232 11144
rect 22928 11092 22980 11144
rect 15384 11024 15436 11076
rect 16948 11024 17000 11076
rect 17224 11024 17276 11076
rect 17592 11024 17644 11076
rect 13176 10956 13228 11008
rect 15292 10956 15344 11008
rect 16304 10956 16356 11008
rect 19800 11024 19852 11076
rect 19524 10956 19576 11008
rect 20628 10956 20680 11008
rect 21456 10956 21508 11008
rect 23572 10956 23624 11008
rect 6884 10854 6936 10906
rect 6948 10854 7000 10906
rect 7012 10854 7064 10906
rect 7076 10854 7128 10906
rect 7140 10854 7192 10906
rect 12818 10854 12870 10906
rect 12882 10854 12934 10906
rect 12946 10854 12998 10906
rect 13010 10854 13062 10906
rect 13074 10854 13126 10906
rect 18752 10854 18804 10906
rect 18816 10854 18868 10906
rect 18880 10854 18932 10906
rect 18944 10854 18996 10906
rect 19008 10854 19060 10906
rect 24686 10854 24738 10906
rect 24750 10854 24802 10906
rect 24814 10854 24866 10906
rect 24878 10854 24930 10906
rect 24942 10854 24994 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2044 10752 2096 10804
rect 1492 10727 1544 10736
rect 1492 10693 1501 10727
rect 1501 10693 1535 10727
rect 1535 10693 1544 10727
rect 1492 10684 1544 10693
rect 4344 10752 4396 10804
rect 4528 10752 4580 10804
rect 5632 10752 5684 10804
rect 5816 10752 5868 10804
rect 6460 10752 6512 10804
rect 7472 10752 7524 10804
rect 8668 10752 8720 10804
rect 9772 10752 9824 10804
rect 10140 10752 10192 10804
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 7564 10684 7616 10736
rect 11796 10752 11848 10804
rect 12256 10752 12308 10804
rect 13268 10752 13320 10804
rect 10876 10684 10928 10736
rect 13176 10684 13228 10736
rect 4344 10659 4396 10668
rect 4344 10625 4351 10659
rect 4351 10625 4385 10659
rect 4385 10625 4396 10659
rect 4344 10616 4396 10625
rect 5816 10616 5868 10668
rect 6184 10616 6236 10668
rect 8576 10616 8628 10668
rect 9404 10616 9456 10668
rect 11244 10616 11296 10668
rect 1308 10548 1360 10600
rect 1768 10548 1820 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4988 10548 5040 10600
rect 5172 10548 5224 10600
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 2964 10412 3016 10464
rect 4988 10412 5040 10464
rect 8300 10548 8352 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 6828 10412 6880 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 8024 10412 8076 10464
rect 13452 10684 13504 10736
rect 14280 10752 14332 10804
rect 16212 10752 16264 10804
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 14188 10684 14240 10736
rect 14648 10684 14700 10736
rect 14740 10727 14792 10736
rect 14740 10693 14749 10727
rect 14749 10693 14783 10727
rect 14783 10693 14792 10727
rect 14740 10684 14792 10693
rect 15108 10684 15160 10736
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 11428 10548 11480 10600
rect 11888 10548 11940 10600
rect 18328 10616 18380 10668
rect 19524 10659 19576 10668
rect 19524 10625 19531 10659
rect 19531 10625 19565 10659
rect 19565 10625 19576 10659
rect 19524 10616 19576 10625
rect 19616 10616 19668 10668
rect 20076 10752 20128 10804
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 20996 10752 21048 10804
rect 20720 10616 20772 10668
rect 13176 10412 13228 10464
rect 13636 10412 13688 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 19156 10455 19208 10464
rect 19156 10421 19165 10455
rect 19165 10421 19199 10455
rect 19199 10421 19208 10455
rect 19156 10412 19208 10421
rect 20720 10412 20772 10464
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 20996 10412 21048 10464
rect 22560 10412 22612 10464
rect 22744 10659 22796 10668
rect 22744 10625 22753 10659
rect 22753 10625 22787 10659
rect 22787 10625 22796 10659
rect 22744 10616 22796 10625
rect 23204 10684 23256 10736
rect 3917 10310 3969 10362
rect 3981 10310 4033 10362
rect 4045 10310 4097 10362
rect 4109 10310 4161 10362
rect 4173 10310 4225 10362
rect 9851 10310 9903 10362
rect 9915 10310 9967 10362
rect 9979 10310 10031 10362
rect 10043 10310 10095 10362
rect 10107 10310 10159 10362
rect 15785 10310 15837 10362
rect 15849 10310 15901 10362
rect 15913 10310 15965 10362
rect 15977 10310 16029 10362
rect 16041 10310 16093 10362
rect 21719 10310 21771 10362
rect 21783 10310 21835 10362
rect 21847 10310 21899 10362
rect 21911 10310 21963 10362
rect 21975 10310 22027 10362
rect 2136 10208 2188 10260
rect 4068 10208 4120 10260
rect 6000 10208 6052 10260
rect 6368 10208 6420 10260
rect 7288 10208 7340 10260
rect 7380 10208 7432 10260
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 14004 10208 14056 10260
rect 17500 10208 17552 10260
rect 18604 10208 18656 10260
rect 19156 10208 19208 10260
rect 20260 10208 20312 10260
rect 20720 10208 20772 10260
rect 2136 10072 2188 10124
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 6184 10140 6236 10192
rect 4804 10115 4856 10124
rect 4804 10081 4838 10115
rect 4838 10081 4856 10115
rect 4804 10072 4856 10081
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 5172 10072 5224 10124
rect 480 10004 532 10056
rect 2872 10004 2924 10056
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 3608 10004 3660 10056
rect 6092 10072 6144 10124
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6460 10072 6512 10124
rect 6736 10115 6788 10124
rect 6736 10081 6770 10115
rect 6770 10081 6788 10115
rect 6736 10072 6788 10081
rect 10876 10072 10928 10124
rect 10692 10004 10744 10056
rect 4896 9868 4948 9920
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 11428 9936 11480 9988
rect 6828 9868 6880 9920
rect 9036 9868 9088 9920
rect 10508 9868 10560 9920
rect 10692 9868 10744 9920
rect 11612 9868 11664 9920
rect 12624 10004 12676 10056
rect 14004 10004 14056 10056
rect 11980 9936 12032 9988
rect 12164 9936 12216 9988
rect 14372 9983 14397 9988
rect 14397 9983 14424 9988
rect 12532 9868 12584 9920
rect 14372 9936 14424 9983
rect 19432 10004 19484 10056
rect 20444 10140 20496 10192
rect 22468 10208 22520 10260
rect 22100 10140 22152 10192
rect 22744 10140 22796 10192
rect 22284 10072 22336 10124
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 24584 10140 24636 10192
rect 25136 10140 25188 10192
rect 20536 9868 20588 9920
rect 22192 9868 22244 9920
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 22744 9868 22796 9920
rect 23020 9868 23072 9920
rect 23756 9911 23808 9920
rect 23756 9877 23765 9911
rect 23765 9877 23799 9911
rect 23799 9877 23808 9911
rect 23756 9868 23808 9877
rect 6884 9766 6936 9818
rect 6948 9766 7000 9818
rect 7012 9766 7064 9818
rect 7076 9766 7128 9818
rect 7140 9766 7192 9818
rect 12818 9766 12870 9818
rect 12882 9766 12934 9818
rect 12946 9766 12998 9818
rect 13010 9766 13062 9818
rect 13074 9766 13126 9818
rect 18752 9766 18804 9818
rect 18816 9766 18868 9818
rect 18880 9766 18932 9818
rect 18944 9766 18996 9818
rect 19008 9766 19060 9818
rect 24686 9766 24738 9818
rect 24750 9766 24802 9818
rect 24814 9766 24866 9818
rect 24878 9766 24930 9818
rect 24942 9766 24994 9818
rect 2412 9664 2464 9716
rect 4160 9664 4212 9716
rect 4436 9664 4488 9716
rect 6368 9664 6420 9716
rect 7380 9664 7432 9716
rect 7840 9664 7892 9716
rect 10140 9664 10192 9716
rect 10600 9664 10652 9716
rect 10692 9664 10744 9716
rect 10876 9664 10928 9716
rect 11244 9707 11296 9716
rect 11244 9673 11253 9707
rect 11253 9673 11287 9707
rect 11287 9673 11296 9707
rect 11244 9664 11296 9673
rect 20 9596 72 9648
rect 1308 9528 1360 9580
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 1584 9528 1636 9537
rect 3148 9596 3200 9648
rect 3516 9596 3568 9648
rect 4712 9528 4764 9580
rect 7840 9528 7892 9580
rect 8390 9571 8442 9580
rect 8390 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8442 9571
rect 8390 9528 8442 9537
rect 1584 9392 1636 9444
rect 2780 9392 2832 9444
rect 3148 9392 3200 9444
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 6368 9460 6420 9512
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 8484 9460 8536 9512
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10508 9528 10560 9580
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 9588 9503 9640 9512
rect 8116 9435 8168 9444
rect 8116 9401 8125 9435
rect 8125 9401 8159 9435
rect 8159 9401 8168 9435
rect 8116 9392 8168 9401
rect 9588 9469 9597 9503
rect 9597 9469 9631 9503
rect 9631 9469 9640 9503
rect 9588 9460 9640 9469
rect 10140 9460 10192 9512
rect 12624 9664 12676 9716
rect 11428 9528 11480 9580
rect 12072 9571 12124 9580
rect 9404 9324 9456 9376
rect 9588 9324 9640 9376
rect 10324 9324 10376 9376
rect 12072 9537 12079 9571
rect 12079 9537 12113 9571
rect 12113 9537 12124 9571
rect 12072 9528 12124 9537
rect 12348 9596 12400 9648
rect 13268 9664 13320 9716
rect 14004 9664 14056 9716
rect 15108 9664 15160 9716
rect 15292 9664 15344 9716
rect 16304 9664 16356 9716
rect 16580 9664 16632 9716
rect 17960 9664 18012 9716
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 22284 9664 22336 9716
rect 22376 9664 22428 9716
rect 23664 9664 23716 9716
rect 18144 9596 18196 9648
rect 12624 9324 12676 9376
rect 14004 9324 14056 9376
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 19800 9596 19852 9648
rect 20536 9528 20588 9580
rect 19340 9460 19392 9512
rect 19524 9460 19576 9512
rect 19616 9460 19668 9512
rect 15108 9392 15160 9444
rect 17960 9392 18012 9444
rect 22192 9528 22244 9580
rect 23848 9596 23900 9648
rect 25688 9596 25740 9648
rect 22376 9528 22428 9580
rect 19524 9324 19576 9376
rect 19708 9324 19760 9376
rect 22100 9324 22152 9376
rect 22192 9367 22244 9376
rect 22192 9333 22201 9367
rect 22201 9333 22235 9367
rect 22235 9333 22244 9367
rect 22192 9324 22244 9333
rect 24584 9460 24636 9512
rect 23020 9324 23072 9376
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 3917 9222 3969 9274
rect 3981 9222 4033 9274
rect 4045 9222 4097 9274
rect 4109 9222 4161 9274
rect 4173 9222 4225 9274
rect 9851 9222 9903 9274
rect 9915 9222 9967 9274
rect 9979 9222 10031 9274
rect 10043 9222 10095 9274
rect 10107 9222 10159 9274
rect 15785 9222 15837 9274
rect 15849 9222 15901 9274
rect 15913 9222 15965 9274
rect 15977 9222 16029 9274
rect 16041 9222 16093 9274
rect 21719 9222 21771 9274
rect 21783 9222 21835 9274
rect 21847 9222 21899 9274
rect 21911 9222 21963 9274
rect 21975 9222 22027 9274
rect 1308 9120 1360 9172
rect 3056 9120 3108 9172
rect 1492 9052 1544 9104
rect 2228 9095 2280 9104
rect 2228 9061 2237 9095
rect 2237 9061 2271 9095
rect 2271 9061 2280 9095
rect 2228 9052 2280 9061
rect 940 8984 992 9036
rect 1952 8916 2004 8968
rect 1860 8848 1912 8900
rect 3240 9120 3292 9172
rect 7472 9120 7524 9172
rect 7840 9120 7892 9172
rect 9588 9120 9640 9172
rect 9036 8984 9088 9036
rect 10600 9120 10652 9172
rect 2412 8848 2464 8900
rect 2596 8891 2648 8900
rect 2596 8857 2605 8891
rect 2605 8857 2639 8891
rect 2639 8857 2648 8891
rect 2596 8848 2648 8857
rect 3424 8916 3476 8968
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 7840 8916 7892 8968
rect 12440 8916 12492 8968
rect 13544 8916 13596 8968
rect 13268 8848 13320 8900
rect 8484 8780 8536 8832
rect 12440 8780 12492 8832
rect 14004 8984 14056 9036
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14424 8959
rect 14372 8916 14424 8925
rect 15752 8959 15804 8968
rect 15752 8925 15759 8959
rect 15759 8925 15793 8959
rect 15793 8925 15804 8959
rect 15752 8916 15804 8925
rect 17224 9120 17276 9172
rect 17684 9120 17736 9172
rect 22468 9120 22520 9172
rect 23296 9120 23348 9172
rect 24032 9120 24084 9172
rect 24124 9120 24176 9172
rect 19616 8984 19668 9036
rect 21272 9027 21324 9036
rect 21272 8993 21281 9027
rect 21281 8993 21315 9027
rect 21315 8993 21324 9027
rect 21272 8984 21324 8993
rect 19156 8916 19208 8968
rect 23848 8984 23900 9036
rect 23940 8984 23992 9036
rect 22560 8916 22612 8968
rect 23572 8916 23624 8968
rect 20444 8848 20496 8900
rect 22376 8848 22428 8900
rect 14832 8780 14884 8832
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 16120 8780 16172 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 17132 8780 17184 8832
rect 17960 8780 18012 8832
rect 22008 8780 22060 8832
rect 6884 8678 6936 8730
rect 6948 8678 7000 8730
rect 7012 8678 7064 8730
rect 7076 8678 7128 8730
rect 7140 8678 7192 8730
rect 12818 8678 12870 8730
rect 12882 8678 12934 8730
rect 12946 8678 12998 8730
rect 13010 8678 13062 8730
rect 13074 8678 13126 8730
rect 18752 8678 18804 8730
rect 18816 8678 18868 8730
rect 18880 8678 18932 8730
rect 18944 8678 18996 8730
rect 19008 8678 19060 8730
rect 24686 8678 24738 8730
rect 24750 8678 24802 8730
rect 24814 8678 24866 8730
rect 24878 8678 24930 8730
rect 24942 8678 24994 8730
rect 1216 8576 1268 8628
rect 1492 8551 1544 8560
rect 1492 8517 1501 8551
rect 1501 8517 1535 8551
rect 1535 8517 1544 8551
rect 1492 8508 1544 8517
rect 1676 8508 1728 8560
rect 8116 8576 8168 8628
rect 10324 8576 10376 8628
rect 10876 8576 10928 8628
rect 12072 8576 12124 8628
rect 12440 8576 12492 8628
rect 13544 8576 13596 8628
rect 13728 8576 13780 8628
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 2228 8440 2280 8492
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 2320 8372 2372 8424
rect 3332 8347 3384 8356
rect 3332 8313 3341 8347
rect 3341 8313 3375 8347
rect 3375 8313 3384 8347
rect 3332 8304 3384 8313
rect 6092 8372 6144 8424
rect 7472 8508 7524 8560
rect 11612 8508 11664 8560
rect 7564 8440 7616 8492
rect 8024 8440 8076 8492
rect 8300 8440 8352 8492
rect 12716 8508 12768 8560
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12164 8440 12216 8492
rect 12348 8440 12400 8492
rect 12532 8440 12584 8492
rect 13452 8508 13504 8560
rect 15108 8576 15160 8628
rect 16304 8576 16356 8628
rect 17040 8576 17092 8628
rect 13912 8440 13964 8492
rect 14648 8440 14700 8492
rect 14740 8440 14792 8492
rect 15660 8508 15712 8560
rect 17316 8508 17368 8560
rect 22100 8576 22152 8628
rect 22192 8576 22244 8628
rect 23756 8576 23808 8628
rect 18604 8508 18656 8560
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 18328 8440 18380 8492
rect 19340 8440 19392 8492
rect 19524 8440 19576 8492
rect 20168 8483 20220 8492
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 21088 8440 21140 8492
rect 23020 8440 23072 8492
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 9036 8372 9088 8424
rect 11152 8372 11204 8424
rect 13820 8372 13872 8424
rect 15568 8372 15620 8424
rect 18144 8372 18196 8424
rect 8116 8304 8168 8356
rect 8392 8304 8444 8356
rect 2320 8236 2372 8288
rect 2688 8236 2740 8288
rect 4896 8236 4948 8288
rect 7196 8236 7248 8288
rect 11244 8236 11296 8288
rect 12992 8236 13044 8288
rect 13268 8236 13320 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 18696 8236 18748 8288
rect 22284 8372 22336 8424
rect 23940 8415 23992 8424
rect 23940 8381 23949 8415
rect 23949 8381 23983 8415
rect 23983 8381 23992 8415
rect 23940 8372 23992 8381
rect 19708 8304 19760 8356
rect 23480 8304 23532 8356
rect 19984 8236 20036 8288
rect 22928 8236 22980 8288
rect 23204 8236 23256 8288
rect 24308 8279 24360 8288
rect 24308 8245 24317 8279
rect 24317 8245 24351 8279
rect 24351 8245 24360 8279
rect 24308 8236 24360 8245
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 9851 8134 9903 8186
rect 9915 8134 9967 8186
rect 9979 8134 10031 8186
rect 10043 8134 10095 8186
rect 10107 8134 10159 8186
rect 15785 8134 15837 8186
rect 15849 8134 15901 8186
rect 15913 8134 15965 8186
rect 15977 8134 16029 8186
rect 16041 8134 16093 8186
rect 21719 8134 21771 8186
rect 21783 8134 21835 8186
rect 21847 8134 21899 8186
rect 21911 8134 21963 8186
rect 21975 8134 22027 8186
rect 1400 8032 1452 8084
rect 1860 8032 1912 8084
rect 2228 8032 2280 8084
rect 2320 8032 2372 8084
rect 2780 7964 2832 8016
rect 2688 7896 2740 7948
rect 5356 8032 5408 8084
rect 2228 7871 2280 7880
rect 1492 7803 1544 7812
rect 1492 7769 1501 7803
rect 1501 7769 1535 7803
rect 1535 7769 1544 7803
rect 1492 7760 1544 7769
rect 1676 7760 1728 7812
rect 2228 7837 2235 7871
rect 2235 7837 2269 7871
rect 2269 7837 2280 7871
rect 2228 7828 2280 7837
rect 2320 7760 2372 7812
rect 3332 7828 3384 7880
rect 4160 7828 4212 7880
rect 4252 7871 4304 7880
rect 4252 7837 4261 7871
rect 4261 7837 4295 7871
rect 4295 7837 4304 7871
rect 4252 7828 4304 7837
rect 4344 7828 4396 7880
rect 7196 8032 7248 8084
rect 7288 8032 7340 8084
rect 11152 8032 11204 8084
rect 11244 8032 11296 8084
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 7196 7939 7248 7948
rect 7196 7905 7205 7939
rect 7205 7905 7239 7939
rect 7239 7905 7248 7939
rect 7196 7896 7248 7905
rect 9772 7896 9824 7948
rect 12072 8032 12124 8084
rect 13820 8032 13872 8084
rect 16488 8032 16540 8084
rect 16856 8032 16908 8084
rect 18144 8032 18196 8084
rect 18604 8032 18656 8084
rect 20168 8032 20220 8084
rect 23020 8032 23072 8084
rect 6368 7828 6420 7880
rect 7380 7828 7432 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 2412 7692 2464 7744
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 3148 7692 3200 7744
rect 4436 7692 4488 7744
rect 5172 7692 5224 7744
rect 8024 7760 8076 7812
rect 9220 7760 9272 7812
rect 10784 7828 10836 7880
rect 12256 7828 12308 7880
rect 12624 7939 12676 7948
rect 12624 7905 12633 7939
rect 12633 7905 12667 7939
rect 12667 7905 12676 7939
rect 12624 7896 12676 7905
rect 15568 7896 15620 7948
rect 17132 7896 17184 7948
rect 12992 7828 13044 7880
rect 13360 7760 13412 7812
rect 8484 7692 8536 7744
rect 11704 7692 11756 7744
rect 12072 7692 12124 7744
rect 13728 7692 13780 7744
rect 15384 7828 15436 7880
rect 15660 7828 15712 7880
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 18604 7828 18656 7880
rect 21272 7896 21324 7948
rect 19524 7828 19576 7880
rect 19892 7828 19944 7880
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 17776 7760 17828 7812
rect 19984 7760 20036 7812
rect 22560 7871 22612 7880
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 22560 7828 22612 7837
rect 22836 7871 22888 7880
rect 22836 7837 22845 7871
rect 22845 7837 22879 7871
rect 22879 7837 22888 7871
rect 22836 7828 22888 7837
rect 17224 7692 17276 7744
rect 18696 7692 18748 7744
rect 20904 7692 20956 7744
rect 21364 7692 21416 7744
rect 22100 7692 22152 7744
rect 23756 7760 23808 7812
rect 6884 7590 6936 7642
rect 6948 7590 7000 7642
rect 7012 7590 7064 7642
rect 7076 7590 7128 7642
rect 7140 7590 7192 7642
rect 12818 7590 12870 7642
rect 12882 7590 12934 7642
rect 12946 7590 12998 7642
rect 13010 7590 13062 7642
rect 13074 7590 13126 7642
rect 18752 7590 18804 7642
rect 18816 7590 18868 7642
rect 18880 7590 18932 7642
rect 18944 7590 18996 7642
rect 19008 7590 19060 7642
rect 24686 7590 24738 7642
rect 24750 7590 24802 7642
rect 24814 7590 24866 7642
rect 24878 7590 24930 7642
rect 24942 7590 24994 7642
rect 756 7488 808 7540
rect 1124 7488 1176 7540
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 2596 7488 2648 7540
rect 2780 7488 2832 7540
rect 1676 7463 1728 7472
rect 1676 7429 1685 7463
rect 1685 7429 1719 7463
rect 1719 7429 1728 7463
rect 1676 7420 1728 7429
rect 4160 7488 4212 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 8484 7488 8536 7540
rect 18420 7488 18472 7540
rect 19892 7488 19944 7540
rect 20628 7488 20680 7540
rect 480 7352 532 7404
rect 2412 7327 2464 7336
rect 2412 7293 2421 7327
rect 2421 7293 2455 7327
rect 2455 7293 2464 7327
rect 2412 7284 2464 7293
rect 2136 7216 2188 7268
rect 2780 7352 2832 7404
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 5448 7352 5500 7404
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 6184 7352 6236 7404
rect 2964 7284 3016 7336
rect 3792 7284 3844 7336
rect 4436 7284 4488 7336
rect 4620 7284 4672 7336
rect 5080 7284 5132 7336
rect 4988 7259 5040 7268
rect 4988 7225 4997 7259
rect 4997 7225 5031 7259
rect 5031 7225 5040 7259
rect 4988 7216 5040 7225
rect 6092 7216 6144 7268
rect 8852 7352 8904 7404
rect 9220 7352 9272 7404
rect 9588 7352 9640 7404
rect 10968 7352 11020 7404
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 10232 7284 10284 7336
rect 12440 7284 12492 7336
rect 8944 7148 8996 7200
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 9220 7148 9272 7200
rect 11060 7216 11112 7268
rect 12624 7420 12676 7472
rect 13452 7420 13504 7472
rect 13820 7420 13872 7472
rect 14740 7420 14792 7472
rect 13912 7352 13964 7404
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 14648 7352 14700 7404
rect 13452 7284 13504 7336
rect 14372 7284 14424 7336
rect 18788 7352 18840 7404
rect 20260 7352 20312 7404
rect 20444 7395 20496 7404
rect 20444 7361 20478 7395
rect 20478 7361 20496 7395
rect 20444 7352 20496 7361
rect 20720 7352 20772 7404
rect 22560 7488 22612 7540
rect 23480 7488 23532 7540
rect 25136 7488 25188 7540
rect 19340 7284 19392 7336
rect 22652 7352 22704 7404
rect 22192 7284 22244 7336
rect 16304 7216 16356 7268
rect 10324 7148 10376 7200
rect 13268 7148 13320 7200
rect 14464 7148 14516 7200
rect 21272 7216 21324 7268
rect 23756 7420 23808 7472
rect 24308 7420 24360 7472
rect 24216 7352 24268 7404
rect 21180 7148 21232 7200
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 9851 7046 9903 7098
rect 9915 7046 9967 7098
rect 9979 7046 10031 7098
rect 10043 7046 10095 7098
rect 10107 7046 10159 7098
rect 15785 7046 15837 7098
rect 15849 7046 15901 7098
rect 15913 7046 15965 7098
rect 15977 7046 16029 7098
rect 16041 7046 16093 7098
rect 21719 7046 21771 7098
rect 21783 7046 21835 7098
rect 21847 7046 21899 7098
rect 21911 7046 21963 7098
rect 21975 7046 22027 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 3608 6944 3660 6996
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 3332 6740 3384 6792
rect 3608 6740 3660 6792
rect 4344 6876 4396 6928
rect 4068 6740 4120 6792
rect 2780 6604 2832 6656
rect 3424 6604 3476 6656
rect 3700 6604 3752 6656
rect 3884 6604 3936 6656
rect 5540 6987 5592 6996
rect 5540 6953 5549 6987
rect 5549 6953 5583 6987
rect 5583 6953 5592 6987
rect 5540 6944 5592 6953
rect 6644 6944 6696 6996
rect 7840 6944 7892 6996
rect 9036 6876 9088 6928
rect 8668 6808 8720 6860
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 13452 6944 13504 6996
rect 17776 6944 17828 6996
rect 18604 6987 18656 6996
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 15476 6876 15528 6928
rect 19616 6944 19668 6996
rect 20260 6944 20312 6996
rect 21088 6987 21140 6996
rect 21088 6953 21097 6987
rect 21097 6953 21131 6987
rect 21131 6953 21140 6987
rect 21088 6944 21140 6953
rect 21272 6944 21324 6996
rect 20352 6919 20404 6928
rect 20352 6885 20361 6919
rect 20361 6885 20395 6919
rect 20395 6885 20404 6919
rect 20352 6876 20404 6885
rect 20536 6876 20588 6928
rect 8944 6808 8996 6817
rect 10324 6808 10376 6860
rect 15384 6808 15436 6860
rect 17868 6808 17920 6860
rect 5816 6740 5868 6792
rect 9312 6740 9364 6792
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 9956 6783 10008 6792
rect 9956 6749 9990 6783
rect 9990 6749 10008 6783
rect 9956 6740 10008 6749
rect 11704 6740 11756 6792
rect 9036 6672 9088 6724
rect 15476 6740 15528 6792
rect 17776 6740 17828 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 19616 6783 19668 6792
rect 19616 6749 19623 6783
rect 19623 6749 19657 6783
rect 19657 6749 19668 6783
rect 19616 6740 19668 6749
rect 20444 6740 20496 6792
rect 22376 6876 22428 6928
rect 23480 6944 23532 6996
rect 22928 6876 22980 6928
rect 23204 6876 23256 6928
rect 20720 6672 20772 6724
rect 13176 6604 13228 6656
rect 15108 6604 15160 6656
rect 17224 6604 17276 6656
rect 19156 6604 19208 6656
rect 21180 6783 21232 6792
rect 21180 6749 21189 6783
rect 21189 6749 21223 6783
rect 21223 6749 21232 6783
rect 21180 6740 21232 6749
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 23296 6808 23348 6860
rect 21088 6672 21140 6724
rect 22744 6783 22796 6792
rect 22744 6749 22753 6783
rect 22753 6749 22787 6783
rect 22787 6749 22796 6783
rect 22744 6740 22796 6749
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 23480 6783 23532 6792
rect 23480 6749 23489 6783
rect 23489 6749 23523 6783
rect 23523 6749 23532 6783
rect 23480 6740 23532 6749
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 21916 6604 21968 6656
rect 22100 6604 22152 6656
rect 22560 6604 22612 6656
rect 23572 6647 23624 6656
rect 23572 6613 23581 6647
rect 23581 6613 23615 6647
rect 23615 6613 23624 6647
rect 23572 6604 23624 6613
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 1308 6400 1360 6452
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 5632 6400 5684 6452
rect 5724 6400 5776 6452
rect 1216 6332 1268 6384
rect 2964 6332 3016 6384
rect 5448 6332 5500 6384
rect 3148 6196 3200 6248
rect 1308 6128 1360 6180
rect 4712 6264 4764 6316
rect 6276 6264 6328 6316
rect 6460 6264 6512 6316
rect 7380 6307 7432 6316
rect 7380 6273 7414 6307
rect 7414 6273 7432 6307
rect 7380 6264 7432 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 8944 6400 8996 6452
rect 9036 6400 9088 6452
rect 9956 6264 10008 6316
rect 11612 6264 11664 6316
rect 3608 6196 3660 6248
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 8116 6196 8168 6248
rect 9404 6196 9456 6248
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 10232 6196 10284 6248
rect 12532 6400 12584 6452
rect 13268 6400 13320 6452
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 1768 6103 1820 6112
rect 1768 6069 1777 6103
rect 1777 6069 1811 6103
rect 1811 6069 1820 6103
rect 1768 6060 1820 6069
rect 3792 6128 3844 6180
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 7380 6060 7432 6112
rect 12440 6239 12492 6259
rect 12440 6207 12449 6239
rect 12449 6207 12483 6239
rect 12483 6207 12492 6239
rect 13912 6400 13964 6452
rect 15476 6400 15528 6452
rect 16764 6400 16816 6452
rect 17684 6400 17736 6452
rect 17868 6400 17920 6452
rect 18236 6400 18288 6452
rect 19064 6400 19116 6452
rect 21088 6400 21140 6452
rect 17500 6332 17552 6384
rect 19892 6332 19944 6384
rect 13728 6303 13753 6316
rect 13753 6303 13780 6316
rect 13728 6264 13780 6303
rect 15108 6264 15160 6316
rect 15200 6307 15252 6316
rect 15200 6273 15207 6307
rect 15207 6273 15241 6307
rect 15241 6273 15252 6307
rect 15200 6264 15252 6273
rect 16396 6264 16448 6316
rect 18236 6264 18288 6316
rect 20628 6332 20680 6384
rect 22054 6400 22106 6452
rect 22744 6400 22796 6452
rect 24216 6400 24268 6452
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20536 6264 20588 6316
rect 9496 6171 9548 6180
rect 9496 6137 9505 6171
rect 9505 6137 9539 6171
rect 9539 6137 9548 6171
rect 9496 6128 9548 6137
rect 10508 6128 10560 6180
rect 12164 6171 12216 6180
rect 12164 6137 12173 6171
rect 12173 6137 12207 6171
rect 12207 6137 12216 6171
rect 12164 6128 12216 6137
rect 13360 6171 13412 6180
rect 13360 6137 13369 6171
rect 13369 6137 13403 6171
rect 13403 6137 13412 6171
rect 13360 6128 13412 6137
rect 11060 6060 11112 6112
rect 11704 6060 11756 6112
rect 18420 6196 18472 6248
rect 21272 6196 21324 6248
rect 18144 6128 18196 6180
rect 20168 6128 20220 6180
rect 20628 6171 20680 6180
rect 20628 6137 20637 6171
rect 20637 6137 20671 6171
rect 20671 6137 20680 6171
rect 20628 6128 20680 6137
rect 20720 6128 20772 6180
rect 21180 6128 21232 6180
rect 21824 6307 21876 6316
rect 21824 6273 21833 6307
rect 21833 6273 21867 6307
rect 21867 6273 21876 6307
rect 21824 6264 21876 6273
rect 22652 6264 22704 6316
rect 23296 6264 23348 6316
rect 16304 6060 16356 6112
rect 20076 6103 20128 6112
rect 20076 6069 20085 6103
rect 20085 6069 20119 6103
rect 20119 6069 20128 6103
rect 20076 6060 20128 6069
rect 20904 6060 20956 6112
rect 21548 6060 21600 6112
rect 23756 6307 23808 6316
rect 23756 6273 23765 6307
rect 23765 6273 23799 6307
rect 23799 6273 23808 6307
rect 23756 6264 23808 6273
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 24216 6196 24268 6248
rect 23480 6103 23532 6112
rect 23480 6069 23489 6103
rect 23489 6069 23523 6103
rect 23523 6069 23532 6103
rect 23480 6060 23532 6069
rect 24124 6103 24176 6112
rect 24124 6069 24133 6103
rect 24133 6069 24167 6103
rect 24167 6069 24176 6103
rect 24124 6060 24176 6069
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 1400 5856 1452 5908
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 1032 5788 1084 5840
rect 3884 5856 3936 5908
rect 5356 5856 5408 5908
rect 5448 5856 5500 5908
rect 6092 5856 6144 5908
rect 3056 5720 3108 5772
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 4712 5720 4764 5772
rect 2044 5627 2096 5636
rect 2044 5593 2053 5627
rect 2053 5593 2087 5627
rect 2087 5593 2096 5627
rect 2044 5584 2096 5593
rect 3884 5652 3936 5704
rect 5264 5652 5316 5704
rect 5908 5720 5960 5772
rect 7564 5856 7616 5908
rect 9496 5856 9548 5908
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 4344 5516 4396 5568
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 6644 5584 6696 5636
rect 10600 5856 10652 5908
rect 12164 5856 12216 5908
rect 12440 5856 12492 5908
rect 14464 5856 14516 5908
rect 14740 5856 14792 5908
rect 14924 5856 14976 5908
rect 15384 5856 15436 5908
rect 9680 5720 9732 5772
rect 7564 5584 7616 5636
rect 10140 5695 10192 5704
rect 10140 5661 10147 5695
rect 10147 5661 10181 5695
rect 10181 5661 10192 5695
rect 10140 5652 10192 5661
rect 11152 5652 11204 5704
rect 12716 5788 12768 5840
rect 16304 5856 16356 5908
rect 16396 5856 16448 5908
rect 12164 5720 12216 5772
rect 12440 5720 12492 5772
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 15384 5720 15436 5772
rect 16304 5763 16356 5772
rect 16304 5729 16338 5763
rect 16338 5729 16356 5763
rect 16304 5720 16356 5729
rect 17132 5720 17184 5772
rect 14924 5652 14976 5704
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 17500 5695 17552 5704
rect 9956 5584 10008 5636
rect 11428 5584 11480 5636
rect 6368 5516 6420 5568
rect 8024 5516 8076 5568
rect 9680 5516 9732 5568
rect 10140 5516 10192 5568
rect 10968 5516 11020 5568
rect 11060 5516 11112 5568
rect 15384 5584 15436 5636
rect 15200 5516 15252 5568
rect 17500 5661 17507 5695
rect 17507 5661 17541 5695
rect 17541 5661 17552 5695
rect 17500 5652 17552 5661
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 19156 5856 19208 5908
rect 20720 5856 20772 5908
rect 23296 5856 23348 5908
rect 23572 5856 23624 5908
rect 24124 5856 24176 5908
rect 21180 5788 21232 5840
rect 23204 5788 23256 5840
rect 19064 5720 19116 5772
rect 20720 5695 20772 5704
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 21088 5652 21140 5704
rect 21548 5695 21600 5704
rect 21548 5661 21557 5695
rect 21557 5661 21591 5695
rect 21591 5661 21600 5695
rect 21548 5652 21600 5661
rect 23572 5652 23624 5704
rect 23940 5695 23992 5704
rect 23940 5661 23949 5695
rect 23949 5661 23983 5695
rect 23983 5661 23992 5695
rect 23940 5652 23992 5661
rect 19064 5516 19116 5568
rect 19248 5516 19300 5568
rect 19524 5516 19576 5568
rect 21456 5516 21508 5568
rect 23204 5516 23256 5568
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 2964 5312 3016 5364
rect 3056 5312 3108 5364
rect 3332 5312 3384 5364
rect 3976 5312 4028 5364
rect 4712 5312 4764 5364
rect 5816 5312 5868 5364
rect 1124 5176 1176 5228
rect 3608 5244 3660 5296
rect 6460 5244 6512 5296
rect 9220 5244 9272 5296
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 10876 5244 10928 5296
rect 3516 5176 3568 5228
rect 4436 5176 4488 5228
rect 1676 4972 1728 5024
rect 4620 5108 4672 5160
rect 5356 5219 5408 5228
rect 5356 5185 5390 5219
rect 5390 5185 5408 5219
rect 5356 5176 5408 5185
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 7472 5176 7524 5228
rect 7564 5176 7616 5228
rect 12624 5176 12676 5228
rect 4896 5108 4948 5160
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5080 5108 5132 5160
rect 5540 5151 5592 5160
rect 5540 5117 5549 5151
rect 5549 5117 5583 5151
rect 5583 5117 5592 5151
rect 5540 5108 5592 5117
rect 9220 5151 9272 5160
rect 9220 5117 9229 5151
rect 9229 5117 9263 5151
rect 9263 5117 9272 5151
rect 9220 5108 9272 5117
rect 10232 5108 10284 5160
rect 14372 5312 14424 5364
rect 13084 5108 13136 5160
rect 13912 5219 13964 5228
rect 13912 5185 13921 5219
rect 13921 5185 13955 5219
rect 13955 5185 13964 5219
rect 13912 5176 13964 5185
rect 15292 5312 15344 5364
rect 15752 5312 15804 5364
rect 16304 5312 16356 5364
rect 17132 5312 17184 5364
rect 18144 5355 18196 5364
rect 18144 5321 18153 5355
rect 18153 5321 18187 5355
rect 18187 5321 18196 5355
rect 18144 5312 18196 5321
rect 18236 5312 18288 5364
rect 15752 5176 15804 5228
rect 17592 5244 17644 5296
rect 13820 5108 13872 5160
rect 14924 5108 14976 5160
rect 15384 5108 15436 5160
rect 16396 5108 16448 5160
rect 17960 5176 18012 5228
rect 18420 5355 18472 5364
rect 18420 5321 18429 5355
rect 18429 5321 18463 5355
rect 18463 5321 18472 5355
rect 18420 5312 18472 5321
rect 18696 5312 18748 5364
rect 19892 5312 19944 5364
rect 20076 5312 20128 5364
rect 19524 5287 19576 5296
rect 19524 5253 19533 5287
rect 19533 5253 19567 5287
rect 19567 5253 19576 5287
rect 19524 5244 19576 5253
rect 20168 5244 20220 5296
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 18972 5176 19024 5228
rect 19432 5176 19484 5228
rect 7564 5040 7616 5092
rect 8300 5040 8352 5092
rect 9956 5040 10008 5092
rect 11152 5040 11204 5092
rect 13360 5083 13412 5092
rect 13360 5049 13369 5083
rect 13369 5049 13403 5083
rect 13403 5049 13412 5083
rect 13360 5040 13412 5049
rect 2504 4972 2556 5024
rect 3608 4972 3660 5024
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 8668 4972 8720 5024
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 15292 5083 15344 5092
rect 15292 5049 15301 5083
rect 15301 5049 15335 5083
rect 15335 5049 15344 5083
rect 15292 5040 15344 5049
rect 16304 5040 16356 5092
rect 17776 4972 17828 5024
rect 19248 5040 19300 5092
rect 20812 5108 20864 5160
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 21548 5219 21600 5228
rect 21548 5185 21557 5219
rect 21557 5185 21591 5219
rect 21591 5185 21600 5219
rect 21548 5176 21600 5185
rect 22284 5176 22336 5228
rect 24216 5312 24268 5364
rect 24308 5176 24360 5228
rect 22100 5108 22152 5160
rect 20904 5040 20956 5092
rect 21180 5040 21232 5092
rect 21456 5040 21508 5092
rect 22836 5040 22888 5092
rect 24216 5040 24268 5092
rect 24584 5040 24636 5092
rect 20536 4972 20588 5024
rect 20996 4972 21048 5024
rect 25504 4972 25556 5024
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 1492 4811 1544 4820
rect 1492 4777 1501 4811
rect 1501 4777 1535 4811
rect 1535 4777 1544 4811
rect 1492 4768 1544 4777
rect 2412 4768 2464 4820
rect 2320 4632 2372 4684
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 3332 4768 3384 4820
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 3516 4632 3568 4684
rect 5264 4768 5316 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 8852 4768 8904 4820
rect 12348 4768 12400 4820
rect 5356 4700 5408 4752
rect 10232 4700 10284 4752
rect 11152 4700 11204 4752
rect 13360 4768 13412 4820
rect 14096 4768 14148 4820
rect 14464 4768 14516 4820
rect 7840 4632 7892 4684
rect 9864 4632 9916 4684
rect 12164 4632 12216 4684
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 4712 4564 4764 4616
rect 4804 4607 4856 4616
rect 4804 4573 4811 4607
rect 4811 4573 4845 4607
rect 4845 4573 4856 4607
rect 4804 4564 4856 4573
rect 4896 4564 4948 4616
rect 14372 4632 14424 4684
rect 15108 4632 15160 4684
rect 16304 4768 16356 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 19248 4768 19300 4820
rect 19524 4768 19576 4820
rect 21088 4768 21140 4820
rect 21180 4768 21232 4820
rect 21548 4768 21600 4820
rect 18788 4743 18840 4752
rect 18788 4709 18797 4743
rect 18797 4709 18831 4743
rect 18831 4709 18840 4743
rect 18788 4700 18840 4709
rect 18972 4700 19024 4752
rect 20904 4700 20956 4752
rect 20720 4632 20772 4684
rect 21088 4632 21140 4684
rect 10324 4564 10376 4616
rect 10876 4564 10928 4616
rect 12808 4564 12860 4616
rect 14096 4564 14148 4616
rect 14924 4564 14976 4616
rect 8024 4496 8076 4548
rect 14556 4496 14608 4548
rect 16120 4564 16172 4616
rect 18604 4564 18656 4616
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 19432 4564 19484 4616
rect 17868 4496 17920 4548
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20352 4564 20404 4616
rect 20536 4607 20588 4616
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 20812 4607 20864 4616
rect 20812 4573 20821 4607
rect 20821 4573 20855 4607
rect 20855 4573 20864 4607
rect 20812 4564 20864 4573
rect 21456 4632 21508 4684
rect 23296 4768 23348 4820
rect 25780 4768 25832 4820
rect 22192 4632 22244 4684
rect 7748 4428 7800 4480
rect 7840 4428 7892 4480
rect 20168 4428 20220 4480
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 20352 4471 20404 4480
rect 20352 4437 20361 4471
rect 20361 4437 20395 4471
rect 20395 4437 20404 4471
rect 20352 4428 20404 4437
rect 21180 4428 21232 4480
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 22468 4607 22520 4616
rect 22468 4573 22477 4607
rect 22477 4573 22511 4607
rect 22511 4573 22520 4607
rect 22468 4564 22520 4573
rect 23112 4564 23164 4616
rect 23204 4496 23256 4548
rect 23848 4496 23900 4548
rect 22100 4471 22152 4480
rect 22100 4437 22109 4471
rect 22109 4437 22143 4471
rect 22143 4437 22152 4471
rect 22100 4428 22152 4437
rect 23572 4428 23624 4480
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 4068 4224 4120 4276
rect 664 4088 716 4140
rect 1860 4088 1912 4140
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2044 3884 2096 3936
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3516 4088 3568 4140
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 3148 4020 3200 4072
rect 5080 4156 5132 4208
rect 6092 4088 6144 4140
rect 7380 4156 7432 4208
rect 7564 4088 7616 4140
rect 4344 4020 4396 4072
rect 9128 4224 9180 4276
rect 10048 4224 10100 4276
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 10232 4156 10284 4208
rect 10324 4131 10376 4140
rect 8668 4020 8720 4072
rect 2504 3952 2556 4004
rect 4160 3884 4212 3936
rect 10324 4097 10331 4131
rect 10331 4097 10365 4131
rect 10365 4097 10376 4131
rect 10324 4088 10376 4097
rect 10416 4088 10468 4140
rect 12348 4224 12400 4276
rect 13176 4224 13228 4276
rect 14740 4224 14792 4276
rect 15292 4224 15344 4276
rect 16304 4224 16356 4276
rect 19892 4224 19944 4276
rect 20076 4224 20128 4276
rect 20628 4224 20680 4276
rect 20996 4224 21048 4276
rect 21640 4224 21692 4276
rect 11704 4088 11756 4140
rect 12716 4156 12768 4208
rect 14372 4088 14424 4140
rect 16764 4156 16816 4208
rect 23756 4156 23808 4208
rect 24584 4156 24636 4208
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 15568 4020 15620 4072
rect 16212 4020 16264 4072
rect 17960 4020 18012 4072
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 19064 4131 19116 4140
rect 19064 4097 19073 4131
rect 19073 4097 19107 4131
rect 19107 4097 19116 4131
rect 19064 4088 19116 4097
rect 19892 4131 19944 4140
rect 19892 4097 19901 4131
rect 19901 4097 19935 4131
rect 19935 4097 19944 4131
rect 19892 4088 19944 4097
rect 20352 4131 20404 4140
rect 20352 4097 20386 4131
rect 20386 4097 20404 4131
rect 20352 4088 20404 4097
rect 20628 4088 20680 4140
rect 22376 4131 22428 4140
rect 22376 4097 22385 4131
rect 22385 4097 22419 4131
rect 22419 4097 22428 4131
rect 22376 4088 22428 4097
rect 19432 4020 19484 4072
rect 22468 4020 22520 4072
rect 22744 4088 22796 4140
rect 24492 4131 24544 4140
rect 24492 4097 24501 4131
rect 24501 4097 24535 4131
rect 24535 4097 24544 4131
rect 24492 4088 24544 4097
rect 19248 3952 19300 4004
rect 21088 3952 21140 4004
rect 24216 4020 24268 4072
rect 24124 3952 24176 4004
rect 9404 3884 9456 3936
rect 9680 3884 9732 3936
rect 10324 3884 10376 3936
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 18328 3927 18380 3936
rect 18328 3893 18337 3927
rect 18337 3893 18371 3927
rect 18371 3893 18380 3927
rect 18328 3884 18380 3893
rect 18696 3884 18748 3936
rect 19156 3884 19208 3936
rect 19616 3884 19668 3936
rect 25136 3884 25188 3936
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2136 3723 2188 3732
rect 2136 3689 2145 3723
rect 2145 3689 2179 3723
rect 2179 3689 2188 3723
rect 2136 3680 2188 3689
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 4896 3723 4948 3732
rect 4896 3689 4905 3723
rect 4905 3689 4939 3723
rect 4939 3689 4948 3723
rect 4896 3680 4948 3689
rect 3700 3544 3752 3596
rect 6368 3680 6420 3732
rect 9128 3680 9180 3732
rect 9404 3680 9456 3732
rect 7288 3612 7340 3664
rect 7380 3612 7432 3664
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 5448 3476 5500 3528
rect 9036 3544 9088 3596
rect 8852 3476 8904 3528
rect 9496 3544 9548 3596
rect 11060 3680 11112 3732
rect 11152 3680 11204 3732
rect 12072 3680 12124 3732
rect 13912 3680 13964 3732
rect 18420 3680 18472 3732
rect 20812 3680 20864 3732
rect 10048 3544 10100 3596
rect 10508 3544 10560 3596
rect 12532 3544 12584 3596
rect 13176 3544 13228 3596
rect 2044 3451 2096 3460
rect 2044 3417 2053 3451
rect 2053 3417 2087 3451
rect 2087 3417 2096 3451
rect 2044 3408 2096 3417
rect 2320 3340 2372 3392
rect 3792 3408 3844 3460
rect 8300 3408 8352 3460
rect 8668 3408 8720 3460
rect 11520 3519 11572 3528
rect 11520 3485 11529 3519
rect 11529 3485 11563 3519
rect 11563 3485 11572 3519
rect 11520 3476 11572 3485
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 10692 3408 10744 3460
rect 13636 3476 13688 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 14280 3476 14332 3528
rect 14832 3476 14884 3528
rect 16304 3476 16356 3528
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 17316 3476 17368 3528
rect 17960 3519 18012 3528
rect 17960 3485 17969 3519
rect 17969 3485 18003 3519
rect 18003 3485 18012 3519
rect 17960 3476 18012 3485
rect 5172 3340 5224 3392
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 6460 3340 6512 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 12348 3451 12400 3460
rect 12348 3417 12357 3451
rect 12357 3417 12391 3451
rect 12391 3417 12400 3451
rect 12348 3408 12400 3417
rect 12440 3451 12492 3460
rect 12440 3417 12449 3451
rect 12449 3417 12483 3451
rect 12483 3417 12492 3451
rect 12440 3408 12492 3417
rect 12532 3408 12584 3460
rect 12900 3408 12952 3460
rect 17408 3340 17460 3392
rect 17776 3383 17828 3392
rect 17776 3349 17785 3383
rect 17785 3349 17819 3383
rect 17819 3349 17828 3383
rect 17776 3340 17828 3349
rect 18052 3340 18104 3392
rect 18512 3408 18564 3460
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 19892 3476 19944 3528
rect 20720 3476 20772 3528
rect 20996 3544 21048 3596
rect 23756 3612 23808 3664
rect 24216 3612 24268 3664
rect 21456 3476 21508 3528
rect 21640 3476 21692 3528
rect 22928 3519 22980 3528
rect 22928 3485 22935 3519
rect 22935 3485 22969 3519
rect 22969 3485 22980 3519
rect 22928 3476 22980 3485
rect 18788 3340 18840 3392
rect 19984 3408 20036 3460
rect 20628 3408 20680 3460
rect 19248 3340 19300 3392
rect 19340 3340 19392 3392
rect 19708 3340 19760 3392
rect 22468 3340 22520 3392
rect 22928 3340 22980 3392
rect 23756 3340 23808 3392
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 2044 3136 2096 3188
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 4436 3136 4488 3188
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 6276 3136 6328 3188
rect 6644 3136 6696 3188
rect 8300 3136 8352 3188
rect 9680 3136 9732 3188
rect 1032 3000 1084 3052
rect 1768 3000 1820 3052
rect 2320 3068 2372 3120
rect 6460 3068 6512 3120
rect 3148 3000 3200 3052
rect 2688 2932 2740 2984
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 9864 3068 9916 3120
rect 10416 3136 10468 3188
rect 11980 3136 12032 3188
rect 12440 3136 12492 3188
rect 14280 3136 14332 3188
rect 18512 3179 18564 3188
rect 18512 3145 18521 3179
rect 18521 3145 18555 3179
rect 18555 3145 18564 3179
rect 18512 3136 18564 3145
rect 4436 3000 4488 3009
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 7748 3000 7800 3052
rect 6092 2932 6144 2984
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 10324 3111 10376 3120
rect 10324 3077 10333 3111
rect 10333 3077 10367 3111
rect 10367 3077 10376 3111
rect 10324 3068 10376 3077
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11060 3111 11112 3120
rect 11060 3077 11069 3111
rect 11069 3077 11103 3111
rect 11103 3077 11112 3111
rect 11060 3068 11112 3077
rect 12072 3043 12124 3052
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 12624 3068 12676 3120
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 17592 3000 17644 3052
rect 17684 3043 17736 3052
rect 17684 3009 17693 3043
rect 17693 3009 17727 3043
rect 17727 3009 17736 3043
rect 17684 3000 17736 3009
rect 18236 3068 18288 3120
rect 18604 3068 18656 3120
rect 19892 3136 19944 3188
rect 20904 3068 20956 3120
rect 24032 3136 24084 3188
rect 9588 2932 9640 2984
rect 10784 2932 10836 2984
rect 11796 2932 11848 2984
rect 11980 2932 12032 2984
rect 19064 3000 19116 3052
rect 20720 3000 20772 3052
rect 21272 3000 21324 3052
rect 23388 3068 23440 3120
rect 5356 2864 5408 2916
rect 6184 2864 6236 2916
rect 6460 2864 6512 2916
rect 8116 2864 8168 2916
rect 8300 2839 8352 2848
rect 8300 2805 8309 2839
rect 8309 2805 8343 2839
rect 8343 2805 8352 2839
rect 8300 2796 8352 2805
rect 8576 2796 8628 2848
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 13452 2796 13504 2848
rect 15476 2839 15528 2848
rect 15476 2805 15485 2839
rect 15485 2805 15519 2839
rect 15519 2805 15528 2839
rect 15476 2796 15528 2805
rect 17224 2839 17276 2848
rect 17224 2805 17233 2839
rect 17233 2805 17267 2839
rect 17267 2805 17276 2839
rect 17224 2796 17276 2805
rect 17500 2839 17552 2848
rect 17500 2805 17509 2839
rect 17509 2805 17543 2839
rect 17543 2805 17552 2839
rect 17500 2796 17552 2805
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 18972 2864 19024 2916
rect 19616 2932 19668 2984
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 20444 2932 20496 2984
rect 22100 2932 22152 2984
rect 20628 2864 20680 2916
rect 22836 2864 22888 2916
rect 24308 3000 24360 3052
rect 25412 2932 25464 2984
rect 18788 2839 18840 2848
rect 18788 2805 18797 2839
rect 18797 2805 18831 2839
rect 18831 2805 18840 2839
rect 18788 2796 18840 2805
rect 19984 2796 20036 2848
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 388 2592 440 2644
rect 2964 2592 3016 2644
rect 3700 2592 3752 2644
rect 3792 2592 3844 2644
rect 5632 2592 5684 2644
rect 6920 2592 6972 2644
rect 7380 2592 7432 2644
rect 8300 2592 8352 2644
rect 8392 2592 8444 2644
rect 9680 2592 9732 2644
rect 5264 2456 5316 2508
rect 480 2388 532 2440
rect 204 2320 256 2372
rect 1676 2320 1728 2372
rect 3056 2388 3108 2440
rect 3240 2388 3292 2440
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 4988 2431 5040 2440
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 940 2252 992 2304
rect 7472 2456 7524 2508
rect 7748 2456 7800 2508
rect 6460 2388 6512 2440
rect 7656 2388 7708 2440
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8392 2456 8444 2508
rect 8484 2456 8536 2508
rect 9772 2524 9824 2576
rect 10784 2592 10836 2644
rect 11244 2592 11296 2644
rect 13268 2635 13320 2644
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 13544 2592 13596 2644
rect 15384 2592 15436 2644
rect 16120 2592 16172 2644
rect 16672 2635 16724 2644
rect 16672 2601 16681 2635
rect 16681 2601 16715 2635
rect 16715 2601 16724 2635
rect 16672 2592 16724 2601
rect 16764 2635 16816 2644
rect 16764 2601 16773 2635
rect 16773 2601 16807 2635
rect 16807 2601 16816 2635
rect 16764 2592 16816 2601
rect 12164 2524 12216 2576
rect 13912 2524 13964 2576
rect 19432 2592 19484 2644
rect 19524 2592 19576 2644
rect 20076 2592 20128 2644
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 8576 2388 8628 2440
rect 8208 2320 8260 2372
rect 5080 2252 5132 2304
rect 5264 2295 5316 2304
rect 5264 2261 5273 2295
rect 5273 2261 5307 2295
rect 5307 2261 5316 2295
rect 5264 2252 5316 2261
rect 5356 2252 5408 2304
rect 5448 2252 5500 2304
rect 6460 2252 6512 2304
rect 7472 2252 7524 2304
rect 7748 2252 7800 2304
rect 8484 2320 8536 2372
rect 8944 2388 8996 2440
rect 9680 2388 9732 2440
rect 11980 2456 12032 2508
rect 19064 2524 19116 2576
rect 19616 2524 19668 2576
rect 14464 2456 14516 2508
rect 10600 2388 10652 2440
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 13268 2388 13320 2440
rect 13544 2431 13596 2440
rect 13544 2397 13553 2431
rect 13553 2397 13587 2431
rect 13587 2397 13596 2431
rect 13544 2388 13596 2397
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14004 2388 14056 2440
rect 14372 2388 14424 2440
rect 15384 2431 15436 2440
rect 15384 2397 15393 2431
rect 15393 2397 15427 2431
rect 15427 2397 15436 2431
rect 15384 2388 15436 2397
rect 17040 2456 17092 2508
rect 16212 2388 16264 2440
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 8944 2295 8996 2304
rect 8944 2261 8953 2295
rect 8953 2261 8987 2295
rect 8987 2261 8996 2295
rect 8944 2252 8996 2261
rect 12532 2320 12584 2372
rect 15108 2320 15160 2372
rect 18972 2456 19024 2508
rect 21088 2499 21140 2508
rect 21088 2465 21097 2499
rect 21097 2465 21131 2499
rect 21131 2465 21140 2499
rect 21088 2456 21140 2465
rect 17684 2388 17736 2440
rect 17868 2388 17920 2440
rect 19340 2388 19392 2440
rect 9680 2252 9732 2304
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12440 2252 12492 2304
rect 13176 2252 13228 2304
rect 14004 2252 14056 2304
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 17592 2363 17644 2372
rect 17592 2329 17601 2363
rect 17601 2329 17635 2363
rect 17635 2329 17644 2363
rect 17592 2320 17644 2329
rect 18512 2320 18564 2372
rect 17040 2295 17092 2304
rect 17040 2261 17049 2295
rect 17049 2261 17083 2295
rect 17083 2261 17092 2295
rect 17040 2252 17092 2261
rect 17132 2252 17184 2304
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 18420 2252 18472 2304
rect 21180 2388 21232 2440
rect 22100 2592 22152 2644
rect 23204 2635 23256 2644
rect 23204 2601 23213 2635
rect 23213 2601 23247 2635
rect 23247 2601 23256 2635
rect 23204 2592 23256 2601
rect 19524 2320 19576 2372
rect 20168 2363 20220 2372
rect 20168 2329 20177 2363
rect 20177 2329 20211 2363
rect 20211 2329 20220 2363
rect 20168 2320 20220 2329
rect 21732 2431 21784 2440
rect 21732 2397 21741 2431
rect 21741 2397 21775 2431
rect 21775 2397 21784 2431
rect 21732 2388 21784 2397
rect 21916 2388 21968 2440
rect 23572 2524 23624 2576
rect 23940 2592 23992 2644
rect 24216 2456 24268 2508
rect 23572 2431 23624 2440
rect 23572 2397 23581 2431
rect 23581 2397 23615 2431
rect 23615 2397 23624 2431
rect 23572 2388 23624 2397
rect 23756 2388 23808 2440
rect 21640 2252 21692 2304
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 1952 1985 2004 2032
rect 1400 1955 1452 1964
rect 1400 1921 1409 1955
rect 1409 1921 1443 1955
rect 1443 1921 1452 1955
rect 1400 1912 1452 1921
rect 1676 1955 1728 1964
rect 1676 1921 1685 1955
rect 1685 1921 1719 1955
rect 1719 1921 1728 1955
rect 1676 1912 1728 1921
rect 1952 1980 1977 1985
rect 1977 1980 2004 1985
rect 2412 2048 2464 2100
rect 3976 2048 4028 2100
rect 4988 2091 5040 2100
rect 4988 2057 4997 2091
rect 4997 2057 5031 2091
rect 5031 2057 5040 2091
rect 4988 2048 5040 2057
rect 5264 2048 5316 2100
rect 5356 2091 5408 2100
rect 5356 2057 5365 2091
rect 5365 2057 5399 2091
rect 5399 2057 5408 2091
rect 5356 2048 5408 2057
rect 3332 1980 3384 2032
rect 3424 1955 3476 1964
rect 3424 1921 3433 1955
rect 3433 1921 3467 1955
rect 3467 1921 3476 1955
rect 3424 1912 3476 1921
rect 4620 1980 4672 2032
rect 6460 2048 6512 2100
rect 3792 1955 3844 1964
rect 3792 1921 3801 1955
rect 3801 1921 3835 1955
rect 3835 1921 3844 1955
rect 3792 1912 3844 1921
rect 4160 1955 4212 1964
rect 4160 1921 4169 1955
rect 4169 1921 4203 1955
rect 4203 1921 4212 1955
rect 4160 1912 4212 1921
rect 5816 2023 5868 2032
rect 5816 1989 5825 2023
rect 5825 1989 5859 2023
rect 5859 1989 5868 2023
rect 5816 1980 5868 1989
rect 6644 2048 6696 2100
rect 6736 2048 6788 2100
rect 3516 1844 3568 1896
rect 5080 1912 5132 1964
rect 6184 1955 6236 1964
rect 6184 1921 6193 1955
rect 6193 1921 6227 1955
rect 6227 1921 6236 1955
rect 6184 1912 6236 1921
rect 6552 1955 6604 1964
rect 6552 1921 6561 1955
rect 6561 1921 6595 1955
rect 6595 1921 6604 1955
rect 6552 1912 6604 1921
rect 7472 2048 7524 2100
rect 7564 2091 7616 2100
rect 7564 2057 7573 2091
rect 7573 2057 7607 2091
rect 7607 2057 7616 2091
rect 7564 2048 7616 2057
rect 8576 2048 8628 2100
rect 8944 2048 8996 2100
rect 9312 2048 9364 2100
rect 10508 2091 10560 2100
rect 10508 2057 10517 2091
rect 10517 2057 10551 2091
rect 10551 2057 10560 2091
rect 10508 2048 10560 2057
rect 11888 2048 11940 2100
rect 13636 2048 13688 2100
rect 14004 2048 14056 2100
rect 15108 2048 15160 2100
rect 5908 1844 5960 1896
rect 7932 1912 7984 1964
rect 3332 1708 3384 1760
rect 5080 1708 5132 1760
rect 7196 1776 7248 1828
rect 8024 1776 8076 1828
rect 8300 1912 8352 1964
rect 10324 1912 10376 1964
rect 11612 1980 11664 2032
rect 12624 1912 12676 1964
rect 13820 1955 13872 1964
rect 13820 1921 13829 1955
rect 13829 1921 13863 1955
rect 13863 1921 13872 1955
rect 13820 1912 13872 1921
rect 14280 1955 14332 1964
rect 14280 1921 14289 1955
rect 14289 1921 14323 1955
rect 14323 1921 14332 1955
rect 14280 1912 14332 1921
rect 15568 1980 15620 2032
rect 17776 2048 17828 2100
rect 17500 1980 17552 2032
rect 19432 2048 19484 2100
rect 19616 2048 19668 2100
rect 22008 2048 22060 2100
rect 22468 2048 22520 2100
rect 22928 2048 22980 2100
rect 23940 2048 23992 2100
rect 15016 1844 15068 1896
rect 16304 1844 16356 1896
rect 16580 1844 16632 1896
rect 18788 1844 18840 1896
rect 21456 2023 21508 2032
rect 21456 1989 21465 2023
rect 21465 1989 21499 2023
rect 21499 1989 21508 2023
rect 21456 1980 21508 1989
rect 20168 1912 20220 1964
rect 20812 1955 20864 1964
rect 20812 1921 20821 1955
rect 20821 1921 20855 1955
rect 20855 1921 20864 1955
rect 20812 1912 20864 1921
rect 21088 1912 21140 1964
rect 24308 2023 24360 2032
rect 24308 1989 24317 2023
rect 24317 1989 24351 2023
rect 24351 1989 24360 2023
rect 24308 1980 24360 1989
rect 14004 1776 14056 1828
rect 15200 1776 15252 1828
rect 15384 1776 15436 1828
rect 11060 1751 11112 1760
rect 11060 1717 11069 1751
rect 11069 1717 11103 1751
rect 11103 1717 11112 1751
rect 11060 1708 11112 1717
rect 11888 1751 11940 1760
rect 11888 1717 11897 1751
rect 11897 1717 11931 1751
rect 11931 1717 11940 1751
rect 11888 1708 11940 1717
rect 12624 1751 12676 1760
rect 12624 1717 12633 1751
rect 12633 1717 12667 1751
rect 12667 1717 12676 1751
rect 12624 1708 12676 1717
rect 13636 1751 13688 1760
rect 13636 1717 13645 1751
rect 13645 1717 13679 1751
rect 13679 1717 13688 1751
rect 13636 1708 13688 1717
rect 14280 1708 14332 1760
rect 14740 1708 14792 1760
rect 15660 1708 15712 1760
rect 18144 1776 18196 1828
rect 20260 1844 20312 1896
rect 21640 1844 21692 1896
rect 23112 1912 23164 1964
rect 23664 1844 23716 1896
rect 22836 1776 22888 1828
rect 24492 1776 24544 1828
rect 16856 1751 16908 1760
rect 16856 1717 16865 1751
rect 16865 1717 16899 1751
rect 16899 1717 16908 1751
rect 16856 1708 16908 1717
rect 17408 1751 17460 1760
rect 17408 1717 17417 1751
rect 17417 1717 17451 1751
rect 17451 1717 17460 1751
rect 17408 1708 17460 1717
rect 17592 1708 17644 1760
rect 19524 1708 19576 1760
rect 21640 1708 21692 1760
rect 25320 1708 25372 1760
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 2780 1547 2832 1556
rect 2780 1513 2789 1547
rect 2789 1513 2823 1547
rect 2823 1513 2832 1547
rect 2780 1504 2832 1513
rect 4896 1504 4948 1556
rect 6552 1504 6604 1556
rect 9312 1504 9364 1556
rect 10692 1504 10744 1556
rect 3332 1436 3384 1488
rect 8852 1436 8904 1488
rect 572 1368 624 1420
rect 1400 1343 1452 1352
rect 1400 1309 1409 1343
rect 1409 1309 1443 1343
rect 1443 1309 1452 1343
rect 1400 1300 1452 1309
rect 1676 1343 1728 1352
rect 1676 1309 1685 1343
rect 1685 1309 1719 1343
rect 1719 1309 1728 1343
rect 1676 1300 1728 1309
rect 1584 1207 1636 1216
rect 1584 1173 1593 1207
rect 1593 1173 1627 1207
rect 1627 1173 1636 1207
rect 1584 1164 1636 1173
rect 1860 1207 1912 1216
rect 1860 1173 1869 1207
rect 1869 1173 1903 1207
rect 1903 1173 1912 1207
rect 1860 1164 1912 1173
rect 3792 1368 3844 1420
rect 4712 1368 4764 1420
rect 2044 1300 2096 1352
rect 2320 1275 2372 1284
rect 2320 1241 2329 1275
rect 2329 1241 2363 1275
rect 2363 1241 2372 1275
rect 2320 1232 2372 1241
rect 2504 1275 2556 1284
rect 2504 1241 2513 1275
rect 2513 1241 2547 1275
rect 2547 1241 2556 1275
rect 2504 1232 2556 1241
rect 3056 1275 3108 1284
rect 3056 1241 3065 1275
rect 3065 1241 3099 1275
rect 3099 1241 3108 1275
rect 3056 1232 3108 1241
rect 3148 1207 3200 1216
rect 3148 1173 3157 1207
rect 3157 1173 3191 1207
rect 3191 1173 3200 1207
rect 3148 1164 3200 1173
rect 3884 1275 3936 1284
rect 3884 1241 3893 1275
rect 3893 1241 3927 1275
rect 3927 1241 3936 1275
rect 3884 1232 3936 1241
rect 4436 1232 4488 1284
rect 3792 1164 3844 1216
rect 4988 1164 5040 1216
rect 5080 1207 5132 1216
rect 5080 1173 5089 1207
rect 5089 1173 5123 1207
rect 5123 1173 5132 1207
rect 5080 1164 5132 1173
rect 5264 1343 5316 1352
rect 5264 1309 5273 1343
rect 5273 1309 5307 1343
rect 5307 1309 5316 1343
rect 5264 1300 5316 1309
rect 5540 1343 5592 1352
rect 5540 1309 5549 1343
rect 5549 1309 5583 1343
rect 5583 1309 5592 1343
rect 5540 1300 5592 1309
rect 6368 1300 6420 1352
rect 8024 1300 8076 1352
rect 9036 1436 9088 1488
rect 9956 1411 10008 1420
rect 9956 1377 9965 1411
rect 9965 1377 9999 1411
rect 9999 1377 10008 1411
rect 9956 1368 10008 1377
rect 11244 1411 11296 1420
rect 11244 1377 11253 1411
rect 11253 1377 11287 1411
rect 11287 1377 11296 1411
rect 11244 1368 11296 1377
rect 6276 1164 6328 1216
rect 6736 1275 6788 1284
rect 6736 1241 6745 1275
rect 6745 1241 6779 1275
rect 6779 1241 6788 1275
rect 6736 1232 6788 1241
rect 7012 1232 7064 1284
rect 9036 1300 9088 1352
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 6460 1164 6512 1216
rect 7564 1207 7616 1216
rect 7564 1173 7573 1207
rect 7573 1173 7607 1207
rect 7607 1173 7616 1207
rect 7564 1164 7616 1173
rect 7748 1164 7800 1216
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 7932 1164 7984 1173
rect 8300 1207 8352 1216
rect 8300 1173 8309 1207
rect 8309 1173 8343 1207
rect 8343 1173 8352 1207
rect 8300 1164 8352 1173
rect 8668 1207 8720 1216
rect 8668 1173 8677 1207
rect 8677 1173 8711 1207
rect 8711 1173 8720 1207
rect 8668 1164 8720 1173
rect 9220 1232 9272 1284
rect 11336 1232 11388 1284
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 13176 1504 13228 1556
rect 13820 1504 13872 1556
rect 14924 1504 14976 1556
rect 15108 1436 15160 1488
rect 16304 1547 16356 1556
rect 16304 1513 16313 1547
rect 16313 1513 16347 1547
rect 16347 1513 16356 1547
rect 16304 1504 16356 1513
rect 16396 1504 16448 1556
rect 16580 1436 16632 1488
rect 17960 1504 18012 1556
rect 18788 1504 18840 1556
rect 12348 1368 12400 1420
rect 13544 1368 13596 1420
rect 10508 1207 10560 1216
rect 10508 1173 10517 1207
rect 10517 1173 10551 1207
rect 10551 1173 10560 1207
rect 10508 1164 10560 1173
rect 11888 1164 11940 1216
rect 12716 1300 12768 1352
rect 12164 1232 12216 1284
rect 12072 1164 12124 1216
rect 13636 1300 13688 1352
rect 16672 1368 16724 1420
rect 20536 1479 20588 1488
rect 20536 1445 20545 1479
rect 20545 1445 20579 1479
rect 20579 1445 20588 1479
rect 20536 1436 20588 1445
rect 22560 1504 22612 1556
rect 23848 1547 23900 1556
rect 23848 1513 23857 1547
rect 23857 1513 23891 1547
rect 23891 1513 23900 1547
rect 23848 1504 23900 1513
rect 25320 1436 25372 1488
rect 18512 1368 18564 1420
rect 21180 1368 21232 1420
rect 22836 1368 22888 1420
rect 13912 1300 13964 1352
rect 14004 1300 14056 1352
rect 15200 1300 15252 1352
rect 15476 1300 15528 1352
rect 16488 1343 16540 1352
rect 16488 1309 16497 1343
rect 16497 1309 16531 1343
rect 16531 1309 16540 1343
rect 16488 1300 16540 1309
rect 17040 1300 17092 1352
rect 17224 1300 17276 1352
rect 17500 1300 17552 1352
rect 18328 1300 18380 1352
rect 19064 1343 19116 1352
rect 19064 1309 19073 1343
rect 19073 1309 19107 1343
rect 19107 1309 19116 1343
rect 19064 1300 19116 1309
rect 20628 1300 20680 1352
rect 17684 1232 17736 1284
rect 21088 1232 21140 1284
rect 21180 1275 21232 1284
rect 21180 1241 21189 1275
rect 21189 1241 21223 1275
rect 21223 1241 21232 1275
rect 21180 1232 21232 1241
rect 21364 1275 21416 1284
rect 21364 1241 21373 1275
rect 21373 1241 21407 1275
rect 21407 1241 21416 1275
rect 21364 1232 21416 1241
rect 21640 1343 21692 1352
rect 21640 1309 21649 1343
rect 21649 1309 21683 1343
rect 21683 1309 21692 1343
rect 21640 1300 21692 1309
rect 23388 1300 23440 1352
rect 22192 1232 22244 1284
rect 23940 1343 23992 1352
rect 23940 1309 23949 1343
rect 23949 1309 23983 1343
rect 23983 1309 23992 1343
rect 23940 1300 23992 1309
rect 13084 1207 13136 1216
rect 13084 1173 13093 1207
rect 13093 1173 13127 1207
rect 13127 1173 13136 1207
rect 13084 1164 13136 1173
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 14004 1164 14056 1216
rect 23296 1164 23348 1216
rect 23940 1164 23992 1216
rect 24124 1207 24176 1216
rect 24124 1173 24133 1207
rect 24133 1173 24167 1207
rect 24167 1173 24176 1207
rect 24124 1164 24176 1173
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 940 960 992 1012
rect 3884 960 3936 1012
rect 5816 960 5868 1012
rect 6736 960 6788 1012
rect 7932 960 7984 1012
rect 10692 960 10744 1012
rect 11704 960 11756 1012
rect 13360 960 13412 1012
rect 18052 960 18104 1012
rect 20720 960 20772 1012
rect 21180 960 21232 1012
rect 1584 892 1636 944
rect 4344 892 4396 944
rect 5172 892 5224 944
rect 6920 892 6972 944
rect 8024 892 8076 944
rect 8300 892 8352 944
rect 11520 892 11572 944
rect 25596 892 25648 944
rect 3148 824 3200 876
rect 1400 688 1452 740
rect 2412 688 2464 740
rect 8668 824 8720 876
rect 12072 824 12124 876
rect 12440 756 12492 808
rect 11152 688 11204 740
rect 4436 620 4488 672
rect 5540 620 5592 672
rect 6368 620 6420 672
rect 9864 620 9916 672
rect 21088 620 21140 672
rect 22008 620 22060 672
rect 7288 552 7340 604
rect 14372 552 14424 604
rect 4988 484 5040 536
rect 12256 484 12308 536
<< metal2 >>
rect 202 44463 258 44623
rect 478 44463 534 44623
rect 754 44463 810 44623
rect 1030 44463 1086 44623
rect 1306 44463 1362 44623
rect 1582 44463 1638 44623
rect 1858 44463 1914 44623
rect 2134 44463 2190 44623
rect 2410 44463 2466 44623
rect 2686 44463 2742 44623
rect 2962 44463 3018 44623
rect 3238 44463 3294 44623
rect 3514 44463 3570 44623
rect 3790 44463 3846 44623
rect 4066 44463 4122 44623
rect 4342 44463 4398 44623
rect 4618 44463 4674 44623
rect 4894 44463 4950 44623
rect 5170 44463 5226 44623
rect 5446 44463 5502 44623
rect 5722 44463 5778 44623
rect 5998 44463 6054 44623
rect 6274 44463 6330 44623
rect 6550 44463 6606 44623
rect 6826 44463 6882 44623
rect 7102 44463 7158 44623
rect 7378 44463 7434 44623
rect 7654 44463 7710 44623
rect 7930 44463 7986 44623
rect 8206 44463 8262 44623
rect 8482 44463 8538 44623
rect 8758 44463 8814 44623
rect 9034 44463 9090 44623
rect 9310 44463 9366 44623
rect 9586 44463 9642 44623
rect 9862 44463 9918 44623
rect 10138 44463 10194 44623
rect 10414 44463 10470 44623
rect 10690 44463 10746 44623
rect 10966 44463 11022 44623
rect 11242 44463 11298 44623
rect 11518 44463 11574 44623
rect 11794 44463 11850 44623
rect 12070 44463 12126 44623
rect 12346 44463 12402 44623
rect 12622 44463 12678 44623
rect 12898 44463 12954 44623
rect 13174 44463 13230 44623
rect 13450 44463 13506 44623
rect 13726 44463 13782 44623
rect 14002 44463 14058 44623
rect 14278 44463 14334 44623
rect 14554 44463 14610 44623
rect 14830 44463 14886 44623
rect 15106 44463 15162 44623
rect 15382 44463 15438 44623
rect 15658 44463 15714 44623
rect 15934 44463 15990 44623
rect 16210 44463 16266 44623
rect 16486 44463 16542 44623
rect 16762 44463 16818 44623
rect 17038 44463 17094 44623
rect 17314 44463 17370 44623
rect 17590 44463 17646 44623
rect 17866 44463 17922 44623
rect 18142 44463 18198 44623
rect 18418 44463 18474 44623
rect 18602 44568 18658 44577
rect 18602 44503 18658 44512
rect 216 43874 244 44463
rect 216 43846 428 43874
rect 400 43382 428 43846
rect 388 43376 440 43382
rect 388 43318 440 43324
rect 492 42362 520 44463
rect 664 43308 716 43314
rect 664 43250 716 43256
rect 480 42356 532 42362
rect 480 42298 532 42304
rect 478 41576 534 41585
rect 478 41511 534 41520
rect 492 36922 520 41511
rect 572 41472 624 41478
rect 572 41414 624 41420
rect 480 36916 532 36922
rect 480 36858 532 36864
rect 480 36712 532 36718
rect 480 36654 532 36660
rect 388 36100 440 36106
rect 388 36042 440 36048
rect 204 34196 256 34202
rect 204 34138 256 34144
rect 20 27464 72 27470
rect 20 27406 72 27412
rect 32 9654 60 27406
rect 216 22094 244 34138
rect 296 33856 348 33862
rect 296 33798 348 33804
rect 308 24177 336 33798
rect 400 24206 428 36042
rect 492 27169 520 36654
rect 584 33862 612 41414
rect 572 33856 624 33862
rect 572 33798 624 33804
rect 572 30592 624 30598
rect 572 30534 624 30540
rect 584 27554 612 30534
rect 676 30394 704 43250
rect 768 41800 796 44463
rect 1044 42106 1072 44463
rect 1320 42786 1348 44463
rect 1320 42770 1440 42786
rect 1320 42764 1452 42770
rect 1320 42758 1400 42764
rect 1400 42706 1452 42712
rect 1044 42078 1348 42106
rect 1320 42022 1348 42078
rect 1308 42016 1360 42022
rect 1308 41958 1360 41964
rect 940 41812 992 41818
rect 768 41772 940 41800
rect 1596 41800 1624 44463
rect 1872 43450 1900 44463
rect 2148 43602 2176 44463
rect 2148 43574 2268 43602
rect 1860 43444 1912 43450
rect 1860 43386 1912 43392
rect 1768 43104 1820 43110
rect 1768 43046 1820 43052
rect 1676 41812 1728 41818
rect 1596 41772 1676 41800
rect 940 41754 992 41760
rect 1676 41754 1728 41760
rect 1124 41676 1176 41682
rect 1124 41618 1176 41624
rect 756 38276 808 38282
rect 756 38218 808 38224
rect 768 37913 796 38218
rect 754 37904 810 37913
rect 754 37839 810 37848
rect 848 37324 900 37330
rect 848 37266 900 37272
rect 756 35080 808 35086
rect 756 35022 808 35028
rect 768 34649 796 35022
rect 754 34640 810 34649
rect 754 34575 810 34584
rect 756 33992 808 33998
rect 756 33934 808 33940
rect 768 31822 796 33934
rect 756 31816 808 31822
rect 756 31758 808 31764
rect 664 30388 716 30394
rect 664 30330 716 30336
rect 860 30002 888 37266
rect 1032 37256 1084 37262
rect 1032 37198 1084 37204
rect 940 36576 992 36582
rect 1044 36553 1072 37198
rect 940 36518 992 36524
rect 1030 36544 1086 36553
rect 676 29974 888 30002
rect 676 27690 704 29974
rect 952 29832 980 36518
rect 1030 36479 1086 36488
rect 1030 35864 1086 35873
rect 1030 35799 1086 35808
rect 1044 33833 1072 35799
rect 1030 33824 1086 33833
rect 1030 33759 1086 33768
rect 1136 31754 1164 41618
rect 1780 41546 1808 43046
rect 2240 42906 2268 43574
rect 2228 42900 2280 42906
rect 2228 42842 2280 42848
rect 2042 42392 2098 42401
rect 2042 42327 2098 42336
rect 2320 42356 2372 42362
rect 2056 42294 2084 42327
rect 2320 42298 2372 42304
rect 2044 42288 2096 42294
rect 2044 42230 2096 42236
rect 2136 42220 2188 42226
rect 2136 42162 2188 42168
rect 1768 41540 1820 41546
rect 1768 41482 1820 41488
rect 1216 41132 1268 41138
rect 1216 41074 1268 41080
rect 1228 39953 1256 41074
rect 1860 40520 1912 40526
rect 1860 40462 1912 40468
rect 1400 40452 1452 40458
rect 1400 40394 1452 40400
rect 1214 39944 1270 39953
rect 1214 39879 1270 39888
rect 1412 39409 1440 40394
rect 1492 40044 1544 40050
rect 1544 40004 1624 40032
rect 1492 39986 1544 39992
rect 1398 39400 1454 39409
rect 1398 39335 1454 39344
rect 1492 39364 1544 39370
rect 1492 39306 1544 39312
rect 1504 39098 1532 39306
rect 1492 39092 1544 39098
rect 1492 39034 1544 39040
rect 1216 38208 1268 38214
rect 1214 38176 1216 38185
rect 1268 38176 1270 38185
rect 1214 38111 1270 38120
rect 1400 37868 1452 37874
rect 1400 37810 1452 37816
rect 1216 37800 1268 37806
rect 1216 37742 1268 37748
rect 1228 33658 1256 37742
rect 1308 37120 1360 37126
rect 1308 37062 1360 37068
rect 1320 36281 1348 37062
rect 1306 36272 1362 36281
rect 1306 36207 1362 36216
rect 1308 36168 1360 36174
rect 1308 36110 1360 36116
rect 1320 34524 1348 36110
rect 1412 35057 1440 37810
rect 1492 37188 1544 37194
rect 1492 37130 1544 37136
rect 1398 35048 1454 35057
rect 1398 34983 1454 34992
rect 1400 34536 1452 34542
rect 1320 34496 1400 34524
rect 1400 34478 1452 34484
rect 1412 33998 1440 34478
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1308 33924 1360 33930
rect 1308 33866 1360 33872
rect 1216 33652 1268 33658
rect 1216 33594 1268 33600
rect 1320 33561 1348 33866
rect 1306 33552 1362 33561
rect 1306 33487 1362 33496
rect 1400 33448 1452 33454
rect 1400 33390 1452 33396
rect 1412 33046 1440 33390
rect 1400 33040 1452 33046
rect 1504 33017 1532 37130
rect 1596 35465 1624 40004
rect 1768 39976 1820 39982
rect 1768 39918 1820 39924
rect 1674 39400 1730 39409
rect 1674 39335 1676 39344
rect 1728 39335 1730 39344
rect 1676 39306 1728 39312
rect 1780 38758 1808 39918
rect 1768 38752 1820 38758
rect 1768 38694 1820 38700
rect 1780 38350 1808 38694
rect 1768 38344 1820 38350
rect 1768 38286 1820 38292
rect 1780 37806 1808 38286
rect 1676 37800 1728 37806
rect 1676 37742 1728 37748
rect 1768 37800 1820 37806
rect 1768 37742 1820 37748
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1688 34649 1716 37742
rect 1780 35494 1808 37742
rect 1872 36106 1900 40462
rect 1952 39296 2004 39302
rect 1952 39238 2004 39244
rect 1964 39098 1992 39238
rect 1952 39092 2004 39098
rect 1952 39034 2004 39040
rect 2148 37330 2176 42162
rect 2226 41168 2282 41177
rect 2226 41103 2228 41112
rect 2280 41103 2282 41112
rect 2228 41074 2280 41080
rect 2228 40112 2280 40118
rect 2228 40054 2280 40060
rect 2240 39681 2268 40054
rect 2332 40050 2360 42298
rect 2424 41274 2452 44463
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 2516 41818 2544 43250
rect 2700 42786 2728 44463
rect 2976 43450 3004 44463
rect 3252 43602 3280 44463
rect 3252 43574 3372 43602
rect 2964 43444 3016 43450
rect 2964 43386 3016 43392
rect 2964 43240 3016 43246
rect 2964 43182 3016 43188
rect 2700 42770 2820 42786
rect 2700 42764 2832 42770
rect 2700 42758 2780 42764
rect 2780 42706 2832 42712
rect 2596 42628 2648 42634
rect 2596 42570 2648 42576
rect 2608 41818 2636 42570
rect 2780 42220 2832 42226
rect 2780 42162 2832 42168
rect 2792 41818 2820 42162
rect 2504 41812 2556 41818
rect 2504 41754 2556 41760
rect 2596 41812 2648 41818
rect 2596 41754 2648 41760
rect 2780 41812 2832 41818
rect 2780 41754 2832 41760
rect 2700 41682 2912 41698
rect 2700 41676 2924 41682
rect 2700 41670 2872 41676
rect 2700 41478 2728 41670
rect 2872 41618 2924 41624
rect 2688 41472 2740 41478
rect 2872 41472 2924 41478
rect 2688 41414 2740 41420
rect 2870 41440 2872 41449
rect 2924 41440 2926 41449
rect 2870 41375 2926 41384
rect 2412 41268 2464 41274
rect 2412 41210 2464 41216
rect 2780 41268 2832 41274
rect 2780 41210 2832 41216
rect 2792 40730 2820 41210
rect 2872 40928 2924 40934
rect 2872 40870 2924 40876
rect 2780 40724 2832 40730
rect 2780 40666 2832 40672
rect 2780 40452 2832 40458
rect 2780 40394 2832 40400
rect 2320 40044 2372 40050
rect 2320 39986 2372 39992
rect 2320 39840 2372 39846
rect 2320 39782 2372 39788
rect 2226 39672 2282 39681
rect 2226 39607 2282 39616
rect 2332 39370 2360 39782
rect 2688 39500 2740 39506
rect 2688 39442 2740 39448
rect 2320 39364 2372 39370
rect 2320 39306 2372 39312
rect 2596 39364 2648 39370
rect 2596 39306 2648 39312
rect 2228 38276 2280 38282
rect 2228 38218 2280 38224
rect 2240 37777 2268 38218
rect 2226 37768 2282 37777
rect 2226 37703 2282 37712
rect 2136 37324 2188 37330
rect 2136 37266 2188 37272
rect 2228 37188 2280 37194
rect 2228 37130 2280 37136
rect 1860 36100 1912 36106
rect 1860 36042 1912 36048
rect 1860 35692 1912 35698
rect 1860 35634 1912 35640
rect 1768 35488 1820 35494
rect 1768 35430 1820 35436
rect 1674 34640 1730 34649
rect 1674 34575 1730 34584
rect 1768 34400 1820 34406
rect 1768 34342 1820 34348
rect 1780 34202 1808 34342
rect 1768 34196 1820 34202
rect 1768 34138 1820 34144
rect 1768 33856 1820 33862
rect 1768 33798 1820 33804
rect 1400 32982 1452 32988
rect 1490 33008 1546 33017
rect 1490 32943 1546 32952
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1308 32768 1360 32774
rect 1308 32710 1360 32716
rect 1216 32564 1268 32570
rect 1216 32506 1268 32512
rect 1228 32201 1256 32506
rect 1320 32473 1348 32710
rect 1306 32464 1362 32473
rect 1306 32399 1362 32408
rect 1214 32192 1270 32201
rect 1214 32127 1270 32136
rect 1308 31816 1360 31822
rect 1308 31758 1360 31764
rect 768 29804 980 29832
rect 1044 31726 1164 31754
rect 768 28529 796 29804
rect 938 29744 994 29753
rect 938 29679 994 29688
rect 952 29238 980 29679
rect 940 29232 992 29238
rect 940 29174 992 29180
rect 1044 28778 1072 31726
rect 1320 31260 1348 31758
rect 1412 31385 1440 32846
rect 1780 32366 1808 33798
rect 1492 32360 1544 32366
rect 1492 32302 1544 32308
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1768 32360 1820 32366
rect 1768 32302 1820 32308
rect 1504 32026 1532 32302
rect 1492 32020 1544 32026
rect 1492 31962 1544 31968
rect 1596 31498 1624 32302
rect 1872 32298 1900 35634
rect 2044 35624 2096 35630
rect 2042 35592 2044 35601
rect 2096 35592 2098 35601
rect 2042 35527 2098 35536
rect 2136 35556 2188 35562
rect 2136 35498 2188 35504
rect 2044 35488 2096 35494
rect 2044 35430 2096 35436
rect 2056 33538 2084 35430
rect 2148 34746 2176 35498
rect 2136 34740 2188 34746
rect 2136 34682 2188 34688
rect 2240 33697 2268 37130
rect 2320 36576 2372 36582
rect 2320 36518 2372 36524
rect 2332 35086 2360 36518
rect 2412 36100 2464 36106
rect 2412 36042 2464 36048
rect 2320 35080 2372 35086
rect 2320 35022 2372 35028
rect 2424 35034 2452 36042
rect 2504 35080 2556 35086
rect 2424 35028 2504 35034
rect 2424 35022 2556 35028
rect 2424 35006 2544 35022
rect 2424 34610 2452 35006
rect 2608 34898 2636 39306
rect 2700 38894 2728 39442
rect 2792 39001 2820 40394
rect 2884 40186 2912 40870
rect 2976 40186 3004 43182
rect 3344 42906 3372 43574
rect 3332 42900 3384 42906
rect 3332 42842 3384 42848
rect 3240 42628 3292 42634
rect 3240 42570 3292 42576
rect 3056 42560 3108 42566
rect 3056 42502 3108 42508
rect 3148 42560 3200 42566
rect 3148 42502 3200 42508
rect 3068 40730 3096 42502
rect 3160 42362 3188 42502
rect 3252 42362 3280 42570
rect 3148 42356 3200 42362
rect 3148 42298 3200 42304
rect 3240 42356 3292 42362
rect 3240 42298 3292 42304
rect 3332 42220 3384 42226
rect 3332 42162 3384 42168
rect 3344 42022 3372 42162
rect 3528 42158 3556 44463
rect 3804 43704 3832 44463
rect 3712 43676 3832 43704
rect 3608 43648 3660 43654
rect 3608 43590 3660 43596
rect 3516 42152 3568 42158
rect 3422 42120 3478 42129
rect 3516 42094 3568 42100
rect 3422 42055 3478 42064
rect 3332 42016 3384 42022
rect 3332 41958 3384 41964
rect 3436 41818 3464 42055
rect 3424 41812 3476 41818
rect 3424 41754 3476 41760
rect 3344 41670 3464 41698
rect 3148 41608 3200 41614
rect 3148 41550 3200 41556
rect 3160 41478 3188 41550
rect 3148 41472 3200 41478
rect 3148 41414 3200 41420
rect 3240 41132 3292 41138
rect 3240 41074 3292 41080
rect 3056 40724 3108 40730
rect 3056 40666 3108 40672
rect 3056 40452 3108 40458
rect 3056 40394 3108 40400
rect 2872 40180 2924 40186
rect 2872 40122 2924 40128
rect 2964 40180 3016 40186
rect 2964 40122 3016 40128
rect 2872 39908 2924 39914
rect 2872 39850 2924 39856
rect 2778 38992 2834 39001
rect 2884 38962 2912 39850
rect 2964 39296 3016 39302
rect 2964 39238 3016 39244
rect 3068 39250 3096 40394
rect 3252 40089 3280 41074
rect 3238 40080 3294 40089
rect 3148 40044 3200 40050
rect 3238 40015 3294 40024
rect 3148 39986 3200 39992
rect 3160 39642 3188 39986
rect 3240 39976 3292 39982
rect 3240 39918 3292 39924
rect 3148 39636 3200 39642
rect 3148 39578 3200 39584
rect 2778 38927 2834 38936
rect 2872 38956 2924 38962
rect 2872 38898 2924 38904
rect 2688 38888 2740 38894
rect 2688 38830 2740 38836
rect 2884 38282 2912 38898
rect 2976 38826 3004 39238
rect 3068 39222 3188 39250
rect 3056 38956 3108 38962
rect 3056 38898 3108 38904
rect 2964 38820 3016 38826
rect 2964 38762 3016 38768
rect 3068 38457 3096 38898
rect 3054 38448 3110 38457
rect 3054 38383 3110 38392
rect 2872 38276 2924 38282
rect 2872 38218 2924 38224
rect 2778 37224 2834 37233
rect 2778 37159 2780 37168
rect 2832 37159 2834 37168
rect 2872 37188 2924 37194
rect 2780 37130 2832 37136
rect 2872 37130 2924 37136
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2792 36242 2820 36722
rect 2780 36236 2832 36242
rect 2780 36178 2832 36184
rect 2688 36032 2740 36038
rect 2688 35974 2740 35980
rect 2700 35698 2728 35974
rect 2688 35692 2740 35698
rect 2688 35634 2740 35640
rect 2608 34870 2728 34898
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 2412 34604 2464 34610
rect 2412 34546 2464 34552
rect 2226 33688 2282 33697
rect 2226 33623 2282 33632
rect 1964 33510 2084 33538
rect 1860 32292 1912 32298
rect 1860 32234 1912 32240
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1780 31498 1808 31622
rect 1596 31470 1808 31498
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1400 31272 1452 31278
rect 1320 31232 1400 31260
rect 1400 31214 1452 31220
rect 1308 31136 1360 31142
rect 1308 31078 1360 31084
rect 1320 30841 1348 31078
rect 1306 30832 1362 30841
rect 1306 30767 1362 30776
rect 1306 30424 1362 30433
rect 1228 30382 1306 30410
rect 1124 29844 1176 29850
rect 1124 29786 1176 29792
rect 1136 29481 1164 29786
rect 1122 29472 1178 29481
rect 1122 29407 1178 29416
rect 1122 28792 1178 28801
rect 1044 28750 1122 28778
rect 1122 28727 1178 28736
rect 938 28656 994 28665
rect 938 28591 994 28600
rect 848 28552 900 28558
rect 754 28520 810 28529
rect 848 28494 900 28500
rect 754 28455 810 28464
rect 860 28121 888 28494
rect 952 28150 980 28591
rect 940 28144 992 28150
rect 846 28112 902 28121
rect 756 28076 808 28082
rect 940 28086 992 28092
rect 846 28047 902 28056
rect 756 28018 808 28024
rect 768 27849 796 28018
rect 754 27840 810 27849
rect 754 27775 810 27784
rect 1228 27690 1256 30382
rect 1306 30359 1362 30368
rect 1412 29866 1440 31214
rect 1492 30660 1544 30666
rect 1492 30602 1544 30608
rect 1504 30025 1532 30602
rect 1596 30598 1624 31470
rect 1964 30870 1992 33510
rect 2424 33318 2452 34546
rect 2412 33312 2464 33318
rect 2412 33254 2464 33260
rect 2042 32872 2098 32881
rect 2042 32807 2098 32816
rect 1952 30864 2004 30870
rect 1952 30806 2004 30812
rect 1584 30592 1636 30598
rect 1584 30534 1636 30540
rect 1676 30184 1728 30190
rect 1676 30126 1728 30132
rect 1490 30016 1546 30025
rect 1490 29951 1546 29960
rect 1412 29838 1532 29866
rect 1504 29646 1532 29838
rect 1584 29776 1636 29782
rect 1582 29744 1584 29753
rect 1636 29744 1638 29753
rect 1582 29679 1638 29688
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1492 29640 1544 29646
rect 1492 29582 1544 29588
rect 1308 29572 1360 29578
rect 1308 29514 1360 29520
rect 1320 29209 1348 29514
rect 1306 29200 1362 29209
rect 1306 29135 1362 29144
rect 1308 28960 1360 28966
rect 1308 28902 1360 28908
rect 676 27662 888 27690
rect 584 27526 704 27554
rect 478 27160 534 27169
rect 478 27095 534 27104
rect 478 26888 534 26897
rect 478 26823 534 26832
rect 388 24200 440 24206
rect 294 24168 350 24177
rect 388 24142 440 24148
rect 294 24103 350 24112
rect 386 23624 442 23633
rect 386 23559 442 23568
rect 216 22066 336 22094
rect 308 17649 336 22066
rect 294 17640 350 17649
rect 294 17575 350 17584
rect 400 17270 428 23559
rect 388 17264 440 17270
rect 388 17206 440 17212
rect 388 16788 440 16794
rect 388 16730 440 16736
rect 20 9648 72 9654
rect 20 9590 72 9596
rect 400 2650 428 16730
rect 492 16266 520 26823
rect 572 26240 624 26246
rect 572 26182 624 26188
rect 584 16386 612 26182
rect 676 22094 704 27526
rect 756 24812 808 24818
rect 756 24754 808 24760
rect 768 23497 796 24754
rect 860 23905 888 27662
rect 952 27662 1256 27690
rect 846 23896 902 23905
rect 846 23831 902 23840
rect 848 23588 900 23594
rect 848 23530 900 23536
rect 754 23488 810 23497
rect 754 23423 810 23432
rect 860 23050 888 23530
rect 848 23044 900 23050
rect 848 22986 900 22992
rect 860 22642 888 22986
rect 848 22636 900 22642
rect 848 22578 900 22584
rect 676 22066 888 22094
rect 860 21690 888 22066
rect 848 21684 900 21690
rect 848 21626 900 21632
rect 846 20360 902 20369
rect 676 20318 846 20346
rect 676 16402 704 20318
rect 846 20295 902 20304
rect 754 20224 810 20233
rect 754 20159 810 20168
rect 768 19854 796 20159
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 756 19848 808 19854
rect 756 19790 808 19796
rect 860 19378 888 19887
rect 848 19372 900 19378
rect 848 19314 900 19320
rect 952 18426 980 27662
rect 1320 27520 1348 28902
rect 1412 27713 1440 29582
rect 1584 29300 1636 29306
rect 1584 29242 1636 29248
rect 1492 29164 1544 29170
rect 1492 29106 1544 29112
rect 1504 28393 1532 29106
rect 1490 28384 1546 28393
rect 1490 28319 1546 28328
rect 1398 27704 1454 27713
rect 1398 27639 1454 27648
rect 1320 27492 1440 27520
rect 1124 27328 1176 27334
rect 1124 27270 1176 27276
rect 1136 26489 1164 27270
rect 1216 27124 1268 27130
rect 1216 27066 1268 27072
rect 1228 26761 1256 27066
rect 1306 27024 1362 27033
rect 1306 26959 1308 26968
rect 1360 26959 1362 26968
rect 1308 26930 1360 26936
rect 1412 26874 1440 27492
rect 1320 26846 1440 26874
rect 1214 26752 1270 26761
rect 1214 26687 1270 26696
rect 1122 26480 1178 26489
rect 1122 26415 1178 26424
rect 1320 26058 1348 26846
rect 1492 26376 1544 26382
rect 1492 26318 1544 26324
rect 1136 26030 1348 26058
rect 1032 25900 1084 25906
rect 1032 25842 1084 25848
rect 1044 23594 1072 25842
rect 1136 24970 1164 26030
rect 1308 25968 1360 25974
rect 1308 25910 1360 25916
rect 1216 25492 1268 25498
rect 1216 25434 1268 25440
rect 1228 25129 1256 25434
rect 1320 25401 1348 25910
rect 1504 25906 1532 26318
rect 1492 25900 1544 25906
rect 1492 25842 1544 25848
rect 1306 25392 1362 25401
rect 1306 25327 1362 25336
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1214 25120 1270 25129
rect 1214 25055 1270 25064
rect 1136 24942 1256 24970
rect 1124 24744 1176 24750
rect 1124 24686 1176 24692
rect 1136 24585 1164 24686
rect 1122 24576 1178 24585
rect 1122 24511 1178 24520
rect 1032 23588 1084 23594
rect 1032 23530 1084 23536
rect 1032 23112 1084 23118
rect 1032 23054 1084 23060
rect 1122 23080 1178 23089
rect 1044 22953 1072 23054
rect 1122 23015 1178 23024
rect 1030 22944 1086 22953
rect 1030 22879 1086 22888
rect 1032 22024 1084 22030
rect 1032 21966 1084 21972
rect 940 18420 992 18426
rect 940 18362 992 18368
rect 1044 17377 1072 21966
rect 1030 17368 1086 17377
rect 1030 17303 1086 17312
rect 1032 17264 1084 17270
rect 1032 17206 1084 17212
rect 572 16380 624 16386
rect 676 16374 888 16402
rect 572 16322 624 16328
rect 492 16238 704 16266
rect 572 16176 624 16182
rect 572 16118 624 16124
rect 480 10056 532 10062
rect 480 9998 532 10004
rect 492 7410 520 9998
rect 480 7404 532 7410
rect 480 7346 532 7352
rect 388 2644 440 2650
rect 388 2586 440 2592
rect 480 2440 532 2446
rect 480 2382 532 2388
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 160 244 2314
rect 492 160 520 2382
rect 584 1426 612 16118
rect 676 4146 704 16238
rect 756 7540 808 7546
rect 756 7482 808 7488
rect 664 4140 716 4146
rect 664 4082 716 4088
rect 768 2774 796 7482
rect 676 2746 796 2774
rect 676 1873 704 2746
rect 662 1864 718 1873
rect 662 1799 718 1808
rect 860 1465 888 16374
rect 940 14408 992 14414
rect 940 14350 992 14356
rect 952 12306 980 14350
rect 940 12300 992 12306
rect 940 12242 992 12248
rect 940 11008 992 11014
rect 940 10950 992 10956
rect 952 10169 980 10950
rect 938 10160 994 10169
rect 938 10095 994 10104
rect 938 9616 994 9625
rect 938 9551 994 9560
rect 952 9042 980 9551
rect 940 9036 992 9042
rect 940 8978 992 8984
rect 1044 7562 1072 17206
rect 952 7534 1072 7562
rect 1136 7546 1164 23015
rect 1228 22030 1256 24942
rect 1308 24880 1360 24886
rect 1308 24822 1360 24828
rect 1320 23769 1348 24822
rect 1412 24041 1440 25230
rect 1492 24812 1544 24818
rect 1492 24754 1544 24760
rect 1398 24032 1454 24041
rect 1398 23967 1454 23976
rect 1306 23760 1362 23769
rect 1306 23695 1362 23704
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1308 22704 1360 22710
rect 1306 22672 1308 22681
rect 1360 22672 1362 22681
rect 1412 22658 1440 23598
rect 1504 23225 1532 24754
rect 1596 24138 1624 29242
rect 1688 26042 1716 30126
rect 1952 30116 2004 30122
rect 1952 30058 2004 30064
rect 1860 29640 1912 29646
rect 1780 29600 1860 29628
rect 1780 29481 1808 29600
rect 1860 29582 1912 29588
rect 1766 29472 1822 29481
rect 1766 29407 1822 29416
rect 1780 27674 1808 29407
rect 1964 29034 1992 30058
rect 2056 30036 2084 32807
rect 2608 32552 2636 34682
rect 2700 33658 2728 34870
rect 2792 34746 2820 36178
rect 2884 35737 2912 37130
rect 3160 36961 3188 39222
rect 3146 36952 3202 36961
rect 3146 36887 3202 36896
rect 3252 36825 3280 39918
rect 3238 36816 3294 36825
rect 3238 36751 3294 36760
rect 3238 36680 3294 36689
rect 3068 36638 3238 36666
rect 2964 36168 3016 36174
rect 2964 36110 3016 36116
rect 2976 35873 3004 36110
rect 2962 35864 3018 35873
rect 2962 35799 3018 35808
rect 2870 35728 2926 35737
rect 2870 35663 2926 35672
rect 3068 35578 3096 36638
rect 3238 36615 3294 36624
rect 3344 36564 3372 41670
rect 3436 41614 3464 41670
rect 3424 41608 3476 41614
rect 3424 41550 3476 41556
rect 3516 41064 3568 41070
rect 3516 41006 3568 41012
rect 3528 40594 3556 41006
rect 3516 40588 3568 40594
rect 3516 40530 3568 40536
rect 3516 39840 3568 39846
rect 3516 39782 3568 39788
rect 3528 39642 3556 39782
rect 3516 39636 3568 39642
rect 3516 39578 3568 39584
rect 3516 39432 3568 39438
rect 3516 39374 3568 39380
rect 3424 38956 3476 38962
rect 3424 38898 3476 38904
rect 3436 37913 3464 38898
rect 3422 37904 3478 37913
rect 3422 37839 3478 37848
rect 3422 37496 3478 37505
rect 3422 37431 3424 37440
rect 3476 37431 3478 37440
rect 3424 37402 3476 37408
rect 3436 37330 3464 37402
rect 3424 37324 3476 37330
rect 3424 37266 3476 37272
rect 3424 36848 3476 36854
rect 3424 36790 3476 36796
rect 2976 35550 3096 35578
rect 3160 36536 3372 36564
rect 2780 34740 2832 34746
rect 2780 34682 2832 34688
rect 2780 34604 2832 34610
rect 2780 34546 2832 34552
rect 2792 34082 2820 34546
rect 2976 34202 3004 35550
rect 3056 35488 3108 35494
rect 3056 35430 3108 35436
rect 2964 34196 3016 34202
rect 2964 34138 3016 34144
rect 2792 34054 2912 34082
rect 2780 33992 2832 33998
rect 2780 33934 2832 33940
rect 2688 33652 2740 33658
rect 2688 33594 2740 33600
rect 2688 33312 2740 33318
rect 2688 33254 2740 33260
rect 2516 32524 2636 32552
rect 2410 32464 2466 32473
rect 2320 32428 2372 32434
rect 2240 32388 2320 32416
rect 2136 31816 2188 31822
rect 2134 31784 2136 31793
rect 2188 31784 2190 31793
rect 2134 31719 2190 31728
rect 2240 31521 2268 32388
rect 2410 32399 2466 32408
rect 2320 32370 2372 32376
rect 2226 31512 2282 31521
rect 2226 31447 2282 31456
rect 2136 31136 2188 31142
rect 2136 31078 2188 31084
rect 2148 30190 2176 31078
rect 2226 30424 2282 30433
rect 2226 30359 2282 30368
rect 2240 30190 2268 30359
rect 2136 30184 2188 30190
rect 2136 30126 2188 30132
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 2056 30008 2176 30036
rect 2042 29064 2098 29073
rect 1952 29028 2004 29034
rect 2042 28999 2044 29008
rect 1952 28970 2004 28976
rect 2096 28999 2098 29008
rect 2044 28970 2096 28976
rect 1950 28248 2006 28257
rect 1950 28183 2006 28192
rect 1858 28112 1914 28121
rect 1858 28047 1914 28056
rect 1872 27946 1900 28047
rect 1860 27940 1912 27946
rect 1860 27882 1912 27888
rect 1768 27668 1820 27674
rect 1768 27610 1820 27616
rect 1780 26382 1808 27610
rect 1860 27396 1912 27402
rect 1860 27338 1912 27344
rect 1872 26489 1900 27338
rect 1858 26480 1914 26489
rect 1858 26415 1914 26424
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1858 26072 1914 26081
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1780 26030 1858 26058
rect 1780 25906 1808 26030
rect 1964 26058 1992 28183
rect 2044 28144 2096 28150
rect 2044 28086 2096 28092
rect 2056 27062 2084 28086
rect 2044 27056 2096 27062
rect 2044 26998 2096 27004
rect 2042 26344 2098 26353
rect 2042 26279 2098 26288
rect 2056 26246 2084 26279
rect 2044 26240 2096 26246
rect 2044 26182 2096 26188
rect 1964 26030 2084 26058
rect 1858 26007 1914 26016
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1872 25378 1900 25842
rect 1952 25696 2004 25702
rect 1952 25638 2004 25644
rect 1780 25350 1900 25378
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1688 24313 1716 25230
rect 1674 24304 1730 24313
rect 1674 24239 1730 24248
rect 1584 24132 1636 24138
rect 1584 24074 1636 24080
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1412 22630 1532 22658
rect 1306 22607 1362 22616
rect 1400 22500 1452 22506
rect 1400 22442 1452 22448
rect 1216 22024 1268 22030
rect 1216 21966 1268 21972
rect 1216 21888 1268 21894
rect 1216 21830 1268 21836
rect 1306 21856 1362 21865
rect 1228 21593 1256 21830
rect 1306 21791 1362 21800
rect 1320 21622 1348 21791
rect 1308 21616 1360 21622
rect 1214 21584 1270 21593
rect 1308 21558 1360 21564
rect 1412 21554 1440 22442
rect 1504 22409 1532 22630
rect 1490 22400 1546 22409
rect 1490 22335 1546 22344
rect 1780 21962 1808 25350
rect 1858 25256 1914 25265
rect 1858 25191 1914 25200
rect 1872 25158 1900 25191
rect 1860 25152 1912 25158
rect 1860 25094 1912 25100
rect 1858 24304 1914 24313
rect 1858 24239 1914 24248
rect 1768 21956 1820 21962
rect 1768 21898 1820 21904
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1780 21593 1808 21626
rect 1766 21584 1822 21593
rect 1214 21519 1270 21528
rect 1400 21548 1452 21554
rect 1766 21519 1822 21528
rect 1400 21490 1452 21496
rect 1308 21344 1360 21350
rect 1214 21312 1270 21321
rect 1308 21286 1360 21292
rect 1214 21247 1270 21256
rect 1228 21010 1256 21247
rect 1320 21049 1348 21286
rect 1306 21040 1362 21049
rect 1216 21004 1268 21010
rect 1306 20975 1362 20984
rect 1216 20946 1268 20952
rect 1780 20942 1808 21519
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1308 20868 1360 20874
rect 1308 20810 1360 20816
rect 1320 20777 1348 20810
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1412 20505 1440 20878
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1308 19780 1360 19786
rect 1308 19722 1360 19728
rect 1320 19689 1348 19722
rect 1306 19680 1362 19689
rect 1306 19615 1362 19624
rect 1412 18970 1440 20334
rect 1872 20058 1900 24239
rect 1964 24138 1992 25638
rect 2056 24954 2084 26030
rect 2148 25430 2176 30008
rect 2424 29646 2452 32399
rect 2516 31482 2544 32524
rect 2594 32428 2646 32434
rect 2594 32370 2646 32376
rect 2608 32026 2636 32370
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2700 31754 2728 33254
rect 2792 32745 2820 33934
rect 2884 33289 2912 34054
rect 2964 33652 3016 33658
rect 2964 33594 3016 33600
rect 2870 33280 2926 33289
rect 2870 33215 2926 33224
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2608 31726 2728 31754
rect 2504 31476 2556 31482
rect 2504 31418 2556 31424
rect 2412 29640 2464 29646
rect 2412 29582 2464 29588
rect 2228 29096 2280 29102
rect 2228 29038 2280 29044
rect 2240 28626 2268 29038
rect 2228 28620 2280 28626
rect 2228 28562 2280 28568
rect 2240 25922 2268 28562
rect 2424 28490 2452 29582
rect 2516 29170 2544 31418
rect 2608 30734 2636 31726
rect 2792 31113 2820 31758
rect 2976 31754 3004 33594
rect 3068 33590 3096 35430
rect 3056 33584 3108 33590
rect 3056 33526 3108 33532
rect 3068 33017 3096 33526
rect 3054 33008 3110 33017
rect 3054 32943 3110 32952
rect 3056 32224 3108 32230
rect 3056 32166 3108 32172
rect 2884 31726 3004 31754
rect 2778 31104 2834 31113
rect 2778 31039 2834 31048
rect 2596 30728 2648 30734
rect 2594 30696 2596 30705
rect 2648 30696 2650 30705
rect 2594 30631 2650 30640
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2596 30184 2648 30190
rect 2596 30126 2648 30132
rect 2608 29730 2636 30126
rect 2700 29850 2728 30194
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 2792 29730 2820 29786
rect 2608 29702 2820 29730
rect 2504 29164 2556 29170
rect 2504 29106 2556 29112
rect 2516 28665 2544 29106
rect 2884 29050 2912 31726
rect 3068 29850 3096 32166
rect 3160 31482 3188 36536
rect 3436 36394 3464 36790
rect 3344 36366 3464 36394
rect 3238 36272 3294 36281
rect 3238 36207 3294 36216
rect 3252 35290 3280 36207
rect 3240 35284 3292 35290
rect 3240 35226 3292 35232
rect 3240 35080 3292 35086
rect 3240 35022 3292 35028
rect 3252 34762 3280 35022
rect 3344 34950 3372 36366
rect 3424 36032 3476 36038
rect 3422 36000 3424 36009
rect 3476 36000 3478 36009
rect 3422 35935 3478 35944
rect 3528 35834 3556 39374
rect 3620 38706 3648 43590
rect 3712 42752 3740 43676
rect 4080 43602 4108 44463
rect 3804 43574 4108 43602
rect 3804 42906 3832 43574
rect 4356 43450 4384 44463
rect 4344 43444 4396 43450
rect 4344 43386 4396 43392
rect 4344 43308 4396 43314
rect 4396 43268 4568 43296
rect 4344 43250 4396 43256
rect 4252 43240 4304 43246
rect 4252 43182 4304 43188
rect 3917 43004 4225 43013
rect 3917 43002 3923 43004
rect 3979 43002 4003 43004
rect 4059 43002 4083 43004
rect 4139 43002 4163 43004
rect 4219 43002 4225 43004
rect 3979 42950 3981 43002
rect 4161 42950 4163 43002
rect 3917 42948 3923 42950
rect 3979 42948 4003 42950
rect 4059 42948 4083 42950
rect 4139 42948 4163 42950
rect 4219 42948 4225 42950
rect 3917 42939 4225 42948
rect 3792 42900 3844 42906
rect 3792 42842 3844 42848
rect 4264 42786 4292 43182
rect 4436 43104 4488 43110
rect 4436 43046 4488 43052
rect 4172 42758 4292 42786
rect 3712 42724 4016 42752
rect 3884 42628 3936 42634
rect 3884 42570 3936 42576
rect 3700 42220 3752 42226
rect 3700 42162 3752 42168
rect 3712 40390 3740 42162
rect 3896 42106 3924 42570
rect 3988 42344 4016 42724
rect 4172 42566 4200 42758
rect 4252 42696 4304 42702
rect 4252 42638 4304 42644
rect 4160 42560 4212 42566
rect 4160 42502 4212 42508
rect 3988 42316 4108 42344
rect 4080 42226 4108 42316
rect 3976 42220 4028 42226
rect 3976 42162 4028 42168
rect 4068 42220 4120 42226
rect 4068 42162 4120 42168
rect 3988 42129 4016 42162
rect 3804 42078 3924 42106
rect 3974 42120 4030 42129
rect 3804 41800 3832 42078
rect 3974 42055 4030 42064
rect 3917 41916 4225 41925
rect 3917 41914 3923 41916
rect 3979 41914 4003 41916
rect 4059 41914 4083 41916
rect 4139 41914 4163 41916
rect 4219 41914 4225 41916
rect 3979 41862 3981 41914
rect 4161 41862 4163 41914
rect 3917 41860 3923 41862
rect 3979 41860 4003 41862
rect 4059 41860 4083 41862
rect 4139 41860 4163 41862
rect 4219 41860 4225 41862
rect 3917 41851 4225 41860
rect 4264 41818 4292 42638
rect 4448 42022 4476 43046
rect 4540 42344 4568 43268
rect 4632 42566 4660 44463
rect 4712 43172 4764 43178
rect 4712 43114 4764 43120
rect 4724 42702 4752 43114
rect 4908 42770 4936 44463
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 4712 42696 4764 42702
rect 4712 42638 4764 42644
rect 4620 42560 4672 42566
rect 4620 42502 4672 42508
rect 4804 42560 4856 42566
rect 4804 42502 4856 42508
rect 4540 42316 4660 42344
rect 4436 42016 4488 42022
rect 4436 41958 4488 41964
rect 4528 42016 4580 42022
rect 4528 41958 4580 41964
rect 3884 41812 3936 41818
rect 3804 41772 3884 41800
rect 3884 41754 3936 41760
rect 4252 41812 4304 41818
rect 4252 41754 4304 41760
rect 4252 41608 4304 41614
rect 4252 41550 4304 41556
rect 3792 41132 3844 41138
rect 3792 41074 3844 41080
rect 3804 40730 3832 41074
rect 3917 40828 4225 40837
rect 3917 40826 3923 40828
rect 3979 40826 4003 40828
rect 4059 40826 4083 40828
rect 4139 40826 4163 40828
rect 4219 40826 4225 40828
rect 3979 40774 3981 40826
rect 4161 40774 4163 40826
rect 3917 40772 3923 40774
rect 3979 40772 4003 40774
rect 4059 40772 4083 40774
rect 4139 40772 4163 40774
rect 4219 40772 4225 40774
rect 3917 40763 4225 40772
rect 3792 40724 3844 40730
rect 3792 40666 3844 40672
rect 3700 40384 3752 40390
rect 3700 40326 3752 40332
rect 3804 39681 3832 40666
rect 3976 40520 4028 40526
rect 3976 40462 4028 40468
rect 3988 39914 4016 40462
rect 4264 40361 4292 41550
rect 4250 40352 4306 40361
rect 4250 40287 4306 40296
rect 4344 40044 4396 40050
rect 4344 39986 4396 39992
rect 3976 39908 4028 39914
rect 3976 39850 4028 39856
rect 3917 39740 4225 39749
rect 3917 39738 3923 39740
rect 3979 39738 4003 39740
rect 4059 39738 4083 39740
rect 4139 39738 4163 39740
rect 4219 39738 4225 39740
rect 3979 39686 3981 39738
rect 4161 39686 4163 39738
rect 3917 39684 3923 39686
rect 3979 39684 4003 39686
rect 4059 39684 4083 39686
rect 4139 39684 4163 39686
rect 4219 39684 4225 39686
rect 3790 39672 3846 39681
rect 3917 39675 4225 39684
rect 3790 39607 3846 39616
rect 3804 38894 3832 39607
rect 4252 39364 4304 39370
rect 4252 39306 4304 39312
rect 3976 39296 4028 39302
rect 3976 39238 4028 39244
rect 3988 39098 4016 39238
rect 3976 39092 4028 39098
rect 3976 39034 4028 39040
rect 3792 38888 3844 38894
rect 3884 38888 3936 38894
rect 3792 38830 3844 38836
rect 3882 38856 3884 38865
rect 3936 38856 3938 38865
rect 3882 38791 3938 38800
rect 3988 38740 4016 39034
rect 3804 38712 4016 38740
rect 3804 38706 3832 38712
rect 3620 38678 3832 38706
rect 3620 37942 3648 38678
rect 3917 38652 4225 38661
rect 3917 38650 3923 38652
rect 3979 38650 4003 38652
rect 4059 38650 4083 38652
rect 4139 38650 4163 38652
rect 4219 38650 4225 38652
rect 3979 38598 3981 38650
rect 4161 38598 4163 38650
rect 3917 38596 3923 38598
rect 3979 38596 4003 38598
rect 4059 38596 4083 38598
rect 4139 38596 4163 38598
rect 4219 38596 4225 38598
rect 3917 38587 4225 38596
rect 3700 38276 3752 38282
rect 3700 38218 3752 38224
rect 3608 37936 3660 37942
rect 3608 37878 3660 37884
rect 3620 36854 3648 37878
rect 3712 37210 3740 38218
rect 4160 37868 4212 37874
rect 4264 37856 4292 39306
rect 4356 38865 4384 39986
rect 4342 38856 4398 38865
rect 4342 38791 4398 38800
rect 4344 38752 4396 38758
rect 4344 38694 4396 38700
rect 4356 38214 4384 38694
rect 4448 38321 4476 41958
rect 4540 41614 4568 41958
rect 4528 41608 4580 41614
rect 4528 41550 4580 41556
rect 4528 40928 4580 40934
rect 4528 40870 4580 40876
rect 4540 39438 4568 40870
rect 4632 39846 4660 42316
rect 4710 42256 4766 42265
rect 4710 42191 4712 42200
rect 4764 42191 4766 42200
rect 4712 42162 4764 42168
rect 4816 41750 4844 42502
rect 5184 42378 5212 44463
rect 5460 43874 5488 44463
rect 5460 43846 5580 43874
rect 5264 43716 5316 43722
rect 5264 43658 5316 43664
rect 4908 42362 5212 42378
rect 4896 42356 5212 42362
rect 4948 42350 5212 42356
rect 4896 42298 4948 42304
rect 5172 42220 5224 42226
rect 5172 42162 5224 42168
rect 4988 42152 5040 42158
rect 4988 42094 5040 42100
rect 4896 42016 4948 42022
rect 4896 41958 4948 41964
rect 4804 41744 4856 41750
rect 4804 41686 4856 41692
rect 4804 41608 4856 41614
rect 4804 41550 4856 41556
rect 4816 41414 4844 41550
rect 4908 41546 4936 41958
rect 5000 41818 5028 42094
rect 4988 41812 5040 41818
rect 4988 41754 5040 41760
rect 5184 41682 5212 42162
rect 5172 41676 5224 41682
rect 5172 41618 5224 41624
rect 4896 41540 4948 41546
rect 4896 41482 4948 41488
rect 4816 41386 4936 41414
rect 4804 40656 4856 40662
rect 4908 40633 4936 41386
rect 4804 40598 4856 40604
rect 4894 40624 4950 40633
rect 4620 39840 4672 39846
rect 4620 39782 4672 39788
rect 4528 39432 4580 39438
rect 4528 39374 4580 39380
rect 4528 39296 4580 39302
rect 4528 39238 4580 39244
rect 4434 38312 4490 38321
rect 4434 38247 4490 38256
rect 4344 38208 4396 38214
rect 4344 38150 4396 38156
rect 4436 38208 4488 38214
rect 4436 38150 4488 38156
rect 4448 38026 4476 38150
rect 4356 37998 4476 38026
rect 4356 37874 4384 37998
rect 4212 37828 4292 37856
rect 4160 37810 4212 37816
rect 3917 37564 4225 37573
rect 3917 37562 3923 37564
rect 3979 37562 4003 37564
rect 4059 37562 4083 37564
rect 4139 37562 4163 37564
rect 4219 37562 4225 37564
rect 3979 37510 3981 37562
rect 4161 37510 4163 37562
rect 3917 37508 3923 37510
rect 3979 37508 4003 37510
rect 4059 37508 4083 37510
rect 4139 37508 4163 37510
rect 4219 37508 4225 37510
rect 3917 37499 4225 37508
rect 3884 37460 3936 37466
rect 3884 37402 3936 37408
rect 3712 37182 3832 37210
rect 3700 37120 3752 37126
rect 3700 37062 3752 37068
rect 3712 36922 3740 37062
rect 3700 36916 3752 36922
rect 3700 36858 3752 36864
rect 3608 36848 3660 36854
rect 3608 36790 3660 36796
rect 3804 36258 3832 37182
rect 3896 37097 3924 37402
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 3882 37088 3938 37097
rect 3882 37023 3938 37032
rect 4080 36689 4108 37130
rect 4264 36854 4292 37828
rect 4344 37868 4396 37874
rect 4344 37810 4396 37816
rect 4252 36848 4304 36854
rect 4252 36790 4304 36796
rect 4066 36680 4122 36689
rect 4066 36615 4122 36624
rect 3917 36476 4225 36485
rect 3917 36474 3923 36476
rect 3979 36474 4003 36476
rect 4059 36474 4083 36476
rect 4139 36474 4163 36476
rect 4219 36474 4225 36476
rect 3979 36422 3981 36474
rect 4161 36422 4163 36474
rect 3917 36420 3923 36422
rect 3979 36420 4003 36422
rect 4059 36420 4083 36422
rect 4139 36420 4163 36422
rect 4219 36420 4225 36422
rect 3917 36411 4225 36420
rect 3712 36230 3832 36258
rect 3884 36304 3936 36310
rect 3884 36246 3936 36252
rect 3712 35986 3740 36230
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3620 35958 3740 35986
rect 3516 35828 3568 35834
rect 3516 35770 3568 35776
rect 3620 35714 3648 35958
rect 3698 35864 3754 35873
rect 3698 35799 3754 35808
rect 3424 35692 3476 35698
rect 3424 35634 3476 35640
rect 3528 35686 3648 35714
rect 3332 34944 3384 34950
rect 3332 34886 3384 34892
rect 3330 34776 3386 34785
rect 3252 34734 3330 34762
rect 3330 34711 3386 34720
rect 3344 34610 3372 34711
rect 3332 34604 3384 34610
rect 3332 34546 3384 34552
rect 3240 33516 3292 33522
rect 3240 33458 3292 33464
rect 3252 32026 3280 33458
rect 3344 32978 3372 34546
rect 3436 34105 3464 35634
rect 3422 34096 3478 34105
rect 3422 34031 3478 34040
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3436 33114 3464 33458
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 3332 32972 3384 32978
rect 3332 32914 3384 32920
rect 3332 32428 3384 32434
rect 3528 32416 3556 35686
rect 3608 35624 3660 35630
rect 3608 35566 3660 35572
rect 3620 34678 3648 35566
rect 3608 34672 3660 34678
rect 3608 34614 3660 34620
rect 3606 32600 3662 32609
rect 3606 32535 3662 32544
rect 3332 32370 3384 32376
rect 3436 32388 3556 32416
rect 3240 32020 3292 32026
rect 3240 31962 3292 31968
rect 3344 31929 3372 32370
rect 3330 31920 3386 31929
rect 3330 31855 3386 31864
rect 3240 31816 3292 31822
rect 3240 31758 3292 31764
rect 3148 31476 3200 31482
rect 3148 31418 3200 31424
rect 3056 29844 3108 29850
rect 2792 29022 2912 29050
rect 2976 29804 3056 29832
rect 2596 28960 2648 28966
rect 2596 28902 2648 28908
rect 2502 28656 2558 28665
rect 2502 28591 2558 28600
rect 2412 28484 2464 28490
rect 2412 28426 2464 28432
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2332 27577 2360 28018
rect 2424 27985 2452 28426
rect 2410 27976 2466 27985
rect 2410 27911 2466 27920
rect 2318 27568 2374 27577
rect 2318 27503 2374 27512
rect 2504 27328 2556 27334
rect 2608 27305 2636 28902
rect 2792 28762 2820 29022
rect 2976 28994 3004 29804
rect 3056 29786 3108 29792
rect 3146 29200 3202 29209
rect 3146 29135 3202 29144
rect 2884 28966 3004 28994
rect 2780 28756 2832 28762
rect 2780 28698 2832 28704
rect 2792 28150 2820 28698
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2686 27976 2742 27985
rect 2686 27911 2688 27920
rect 2740 27911 2742 27920
rect 2688 27882 2740 27888
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2688 27396 2740 27402
rect 2688 27338 2740 27344
rect 2504 27270 2556 27276
rect 2594 27296 2650 27305
rect 2320 26988 2372 26994
rect 2320 26930 2372 26936
rect 2412 26988 2464 26994
rect 2412 26930 2464 26936
rect 2332 26450 2360 26930
rect 2424 26586 2452 26930
rect 2516 26926 2544 27270
rect 2594 27231 2650 27240
rect 2504 26920 2556 26926
rect 2504 26862 2556 26868
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 2608 26330 2636 27231
rect 2700 27062 2728 27338
rect 2688 27056 2740 27062
rect 2688 26998 2740 27004
rect 2516 26302 2636 26330
rect 2240 25894 2360 25922
rect 2228 25764 2280 25770
rect 2228 25706 2280 25712
rect 2240 25498 2268 25706
rect 2228 25492 2280 25498
rect 2228 25434 2280 25440
rect 2136 25424 2188 25430
rect 2136 25366 2188 25372
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 2044 24948 2096 24954
rect 2044 24890 2096 24896
rect 2148 24857 2176 25230
rect 2134 24848 2190 24857
rect 2134 24783 2190 24792
rect 2332 24290 2360 25894
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2240 24262 2360 24290
rect 1952 24132 2004 24138
rect 1952 24074 2004 24080
rect 2240 23730 2268 24262
rect 2320 24132 2372 24138
rect 2320 24074 2372 24080
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2056 23322 2084 23666
rect 2228 23588 2280 23594
rect 2228 23530 2280 23536
rect 2240 23322 2268 23530
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 2228 23316 2280 23322
rect 2228 23258 2280 23264
rect 2056 22094 2084 23258
rect 2332 22522 2360 24074
rect 2424 23866 2452 24550
rect 2412 23860 2464 23866
rect 2412 23802 2464 23808
rect 2516 23594 2544 26302
rect 2596 26240 2648 26246
rect 2594 26208 2596 26217
rect 2792 26234 2820 27814
rect 2648 26208 2650 26217
rect 2594 26143 2650 26152
rect 2700 26206 2820 26234
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2608 25702 2636 25978
rect 2700 25906 2728 26206
rect 2688 25900 2740 25906
rect 2688 25842 2740 25848
rect 2596 25696 2648 25702
rect 2596 25638 2648 25644
rect 2686 25528 2742 25537
rect 2686 25463 2742 25472
rect 2700 25294 2728 25463
rect 2688 25288 2740 25294
rect 2688 25230 2740 25236
rect 2778 24984 2834 24993
rect 2778 24919 2834 24928
rect 2884 24936 2912 28966
rect 3054 28792 3110 28801
rect 3054 28727 3110 28736
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2976 28218 3004 28494
rect 2964 28212 3016 28218
rect 2964 28154 3016 28160
rect 3068 27062 3096 28727
rect 3160 27146 3188 29135
rect 3252 29050 3280 31758
rect 3332 31272 3384 31278
rect 3332 31214 3384 31220
rect 3344 30938 3372 31214
rect 3332 30932 3384 30938
rect 3332 30874 3384 30880
rect 3436 30682 3464 32388
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3528 31890 3556 31962
rect 3516 31884 3568 31890
rect 3516 31826 3568 31832
rect 3344 30654 3464 30682
rect 3344 30138 3372 30654
rect 3422 30560 3478 30569
rect 3422 30495 3478 30504
rect 3436 30258 3464 30495
rect 3424 30252 3476 30258
rect 3424 30194 3476 30200
rect 3422 30152 3478 30161
rect 3344 30110 3422 30138
rect 3422 30087 3478 30096
rect 3332 29572 3384 29578
rect 3332 29514 3384 29520
rect 3344 29238 3372 29514
rect 3332 29232 3384 29238
rect 3332 29174 3384 29180
rect 3252 29022 3464 29050
rect 3240 28960 3292 28966
rect 3240 28902 3292 28908
rect 3252 28014 3280 28902
rect 3332 28416 3384 28422
rect 3332 28358 3384 28364
rect 3344 28218 3372 28358
rect 3332 28212 3384 28218
rect 3332 28154 3384 28160
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 3160 27118 3280 27146
rect 3056 27056 3108 27062
rect 3056 26998 3108 27004
rect 3148 27056 3200 27062
rect 3148 26998 3200 27004
rect 2964 26988 3016 26994
rect 2964 26930 3016 26936
rect 2976 26518 3004 26930
rect 2964 26512 3016 26518
rect 2964 26454 3016 26460
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 2976 25401 3004 26318
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 2962 25392 3018 25401
rect 2962 25327 3018 25336
rect 3068 24954 3096 25638
rect 2964 24948 3016 24954
rect 2792 24818 2820 24919
rect 2884 24908 2964 24936
rect 2964 24890 3016 24896
rect 3056 24948 3108 24954
rect 3056 24890 3108 24896
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2608 24682 2820 24698
rect 2596 24676 2820 24682
rect 2648 24670 2820 24676
rect 2596 24618 2648 24624
rect 2792 24410 2820 24670
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2976 24274 3004 24890
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2504 23588 2556 23594
rect 2504 23530 2556 23536
rect 2608 23322 2636 24210
rect 3068 24154 3096 24890
rect 3160 24857 3188 26998
rect 3252 26586 3280 27118
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3240 26580 3292 26586
rect 3240 26522 3292 26528
rect 3252 26382 3280 26522
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3344 25906 3372 26930
rect 3332 25900 3384 25906
rect 3252 25860 3332 25888
rect 3252 25498 3280 25860
rect 3332 25842 3384 25848
rect 3332 25696 3384 25702
rect 3332 25638 3384 25644
rect 3240 25492 3292 25498
rect 3240 25434 3292 25440
rect 3146 24848 3202 24857
rect 3146 24783 3202 24792
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 2976 24126 3096 24154
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2870 24032 2926 24041
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2504 23044 2556 23050
rect 2504 22986 2556 22992
rect 2516 22953 2544 22986
rect 2502 22944 2558 22953
rect 2502 22879 2558 22888
rect 2700 22778 2728 24006
rect 2870 23967 2926 23976
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2884 22642 2912 23967
rect 2872 22636 2924 22642
rect 2872 22578 2924 22584
rect 2332 22494 2544 22522
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2056 22066 2176 22094
rect 2044 21956 2096 21962
rect 2044 21898 2096 21904
rect 2056 20641 2084 21898
rect 2148 20806 2176 22066
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 21690 2360 22034
rect 2424 22030 2452 22374
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2516 21690 2544 22494
rect 2596 22500 2648 22506
rect 2596 22442 2648 22448
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2608 21554 2636 22442
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2596 21548 2648 21554
rect 2596 21490 2648 21496
rect 2318 21040 2374 21049
rect 2318 20975 2374 20984
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2042 20632 2098 20641
rect 2042 20567 2098 20576
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 1860 20052 1912 20058
rect 1860 19994 1912 20000
rect 2056 19854 2084 20402
rect 2148 19922 2176 20742
rect 2226 19952 2282 19961
rect 2136 19916 2188 19922
rect 2226 19887 2282 19896
rect 2136 19858 2188 19864
rect 2044 19848 2096 19854
rect 1582 19816 1638 19825
rect 2044 19790 2096 19796
rect 1582 19751 1638 19760
rect 1596 19514 1624 19751
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1766 19408 1822 19417
rect 1766 19343 1822 19352
rect 1860 19372 1912 19378
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1398 18864 1454 18873
rect 1398 18799 1454 18808
rect 1584 18828 1636 18834
rect 1308 18692 1360 18698
rect 1308 18634 1360 18640
rect 1216 18352 1268 18358
rect 1320 18329 1348 18634
rect 1216 18294 1268 18300
rect 1306 18320 1362 18329
rect 1228 18057 1256 18294
rect 1306 18255 1362 18264
rect 1214 18048 1270 18057
rect 1214 17983 1270 17992
rect 1412 17678 1440 18799
rect 1584 18770 1636 18776
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 18193 1532 18226
rect 1596 18222 1624 18770
rect 1674 18592 1730 18601
rect 1674 18527 1730 18536
rect 1584 18216 1636 18222
rect 1490 18184 1546 18193
rect 1584 18158 1636 18164
rect 1490 18119 1546 18128
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1504 17354 1532 18022
rect 1596 17921 1624 18022
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1688 17762 1716 18527
rect 1412 17326 1532 17354
rect 1596 17734 1716 17762
rect 1412 15450 1440 17326
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1320 15422 1440 15450
rect 1320 15162 1348 15422
rect 1398 15328 1454 15337
rect 1398 15263 1454 15272
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 1306 13696 1362 13705
rect 1306 13631 1362 13640
rect 1216 13524 1268 13530
rect 1216 13466 1268 13472
rect 1228 13161 1256 13466
rect 1320 13462 1348 13631
rect 1308 13456 1360 13462
rect 1308 13398 1360 13404
rect 1412 13394 1440 15263
rect 1504 13870 1532 17167
rect 1596 16590 1624 17734
rect 1780 17660 1808 19343
rect 1860 19314 1912 19320
rect 1872 18601 1900 19314
rect 1858 18592 1914 18601
rect 1858 18527 1914 18536
rect 1872 18290 1900 18527
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1688 17632 1808 17660
rect 1688 16658 1716 17632
rect 1766 17504 1822 17513
rect 1766 17439 1822 17448
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1780 15706 1808 17439
rect 1872 16114 1900 17818
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1584 15632 1636 15638
rect 1584 15574 1636 15580
rect 1596 14006 1624 15574
rect 1872 15570 1900 16050
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 1964 15502 1992 19450
rect 2056 19378 2084 19790
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 2148 17882 2176 19858
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2056 16969 2084 17070
rect 2148 17066 2176 17614
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2042 16960 2098 16969
rect 2042 16895 2098 16904
rect 2042 16824 2098 16833
rect 2042 16759 2098 16768
rect 2056 16182 2084 16759
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 2148 15706 2176 17002
rect 2240 16658 2268 19887
rect 2332 18766 2360 20975
rect 2778 20496 2834 20505
rect 2596 20460 2648 20466
rect 2778 20431 2834 20440
rect 2596 20402 2648 20408
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2332 18290 2360 18702
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2424 17134 2452 20198
rect 2608 19122 2636 20402
rect 2516 19094 2636 19122
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2318 16960 2374 16969
rect 2516 16946 2544 19094
rect 2700 17882 2728 19110
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2792 17678 2820 20431
rect 2884 19825 2912 21830
rect 2976 21078 3004 24126
rect 3252 23322 3280 24754
rect 3344 23730 3372 25638
rect 3436 23746 3464 29022
rect 3528 28422 3556 31826
rect 3620 29850 3648 32535
rect 3712 32502 3740 35799
rect 3804 35193 3832 36110
rect 3896 35630 3924 36246
rect 4068 36100 4120 36106
rect 4068 36042 4120 36048
rect 4080 36009 4108 36042
rect 4066 36000 4122 36009
rect 4066 35935 4122 35944
rect 3884 35624 3936 35630
rect 3884 35566 3936 35572
rect 3917 35388 4225 35397
rect 3917 35386 3923 35388
rect 3979 35386 4003 35388
rect 4059 35386 4083 35388
rect 4139 35386 4163 35388
rect 4219 35386 4225 35388
rect 3979 35334 3981 35386
rect 4161 35334 4163 35386
rect 3917 35332 3923 35334
rect 3979 35332 4003 35334
rect 4059 35332 4083 35334
rect 4139 35332 4163 35334
rect 4219 35332 4225 35334
rect 3917 35323 4225 35332
rect 3790 35184 3846 35193
rect 3790 35119 3846 35128
rect 4264 35086 4292 36790
rect 4356 36786 4384 37810
rect 4344 36780 4396 36786
rect 4344 36722 4396 36728
rect 4540 35766 4568 39238
rect 4632 38457 4660 39782
rect 4816 39506 4844 40598
rect 4894 40559 4950 40568
rect 5080 40384 5132 40390
rect 5080 40326 5132 40332
rect 4804 39500 4856 39506
rect 4804 39442 4856 39448
rect 4712 39364 4764 39370
rect 4712 39306 4764 39312
rect 4618 38448 4674 38457
rect 4618 38383 4674 38392
rect 4724 38214 4752 39306
rect 4988 39296 5040 39302
rect 4988 39238 5040 39244
rect 5000 38826 5028 39238
rect 4988 38820 5040 38826
rect 4988 38762 5040 38768
rect 4712 38208 4764 38214
rect 4712 38150 4764 38156
rect 4804 38208 4856 38214
rect 4804 38150 4856 38156
rect 4896 38208 4948 38214
rect 4896 38150 4948 38156
rect 4816 38010 4844 38150
rect 4804 38004 4856 38010
rect 4804 37946 4856 37952
rect 4712 37868 4764 37874
rect 4712 37810 4764 37816
rect 4724 36786 4752 37810
rect 4804 37188 4856 37194
rect 4804 37130 4856 37136
rect 4816 36854 4844 37130
rect 4908 37126 4936 38150
rect 5000 38010 5028 38762
rect 4988 38004 5040 38010
rect 4988 37946 5040 37952
rect 4988 37868 5040 37874
rect 4988 37810 5040 37816
rect 5000 37466 5028 37810
rect 4988 37460 5040 37466
rect 4988 37402 5040 37408
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 4896 37120 4948 37126
rect 4896 37062 4948 37068
rect 4804 36848 4856 36854
rect 4804 36790 4856 36796
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 4712 36780 4764 36786
rect 4712 36722 4764 36728
rect 4528 35760 4580 35766
rect 4528 35702 4580 35708
rect 4528 35624 4580 35630
rect 4526 35592 4528 35601
rect 4580 35592 4582 35601
rect 4526 35527 4582 35536
rect 4252 35080 4304 35086
rect 4252 35022 4304 35028
rect 4344 35012 4396 35018
rect 4344 34954 4396 34960
rect 3792 34944 3844 34950
rect 3792 34886 3844 34892
rect 3804 34082 3832 34886
rect 4356 34746 4384 34954
rect 4436 34944 4488 34950
rect 4436 34886 4488 34892
rect 4344 34740 4396 34746
rect 4344 34682 4396 34688
rect 3976 34672 4028 34678
rect 3976 34614 4028 34620
rect 3988 34388 4016 34614
rect 4160 34604 4212 34610
rect 4160 34546 4212 34552
rect 4066 34504 4122 34513
rect 4172 34490 4200 34546
rect 4122 34462 4200 34490
rect 4066 34439 4122 34448
rect 3988 34360 4292 34388
rect 3917 34300 4225 34309
rect 3917 34298 3923 34300
rect 3979 34298 4003 34300
rect 4059 34298 4083 34300
rect 4139 34298 4163 34300
rect 4219 34298 4225 34300
rect 3979 34246 3981 34298
rect 4161 34246 4163 34298
rect 3917 34244 3923 34246
rect 3979 34244 4003 34246
rect 4059 34244 4083 34246
rect 4139 34244 4163 34246
rect 4219 34244 4225 34246
rect 3917 34235 4225 34244
rect 3804 34054 3924 34082
rect 3792 33652 3844 33658
rect 3792 33594 3844 33600
rect 3804 33522 3832 33594
rect 3792 33516 3844 33522
rect 3792 33458 3844 33464
rect 3896 33402 3924 34054
rect 4066 33960 4122 33969
rect 4066 33895 4068 33904
rect 4120 33895 4122 33904
rect 4068 33866 4120 33872
rect 3804 33374 3924 33402
rect 3700 32496 3752 32502
rect 3700 32438 3752 32444
rect 3804 32314 3832 33374
rect 3917 33212 4225 33221
rect 3917 33210 3923 33212
rect 3979 33210 4003 33212
rect 4059 33210 4083 33212
rect 4139 33210 4163 33212
rect 4219 33210 4225 33212
rect 3979 33158 3981 33210
rect 4161 33158 4163 33210
rect 3917 33156 3923 33158
rect 3979 33156 4003 33158
rect 4059 33156 4083 33158
rect 4139 33156 4163 33158
rect 4219 33156 4225 33158
rect 3917 33147 4225 33156
rect 4160 32972 4212 32978
rect 4160 32914 4212 32920
rect 4172 32434 4200 32914
rect 4160 32428 4212 32434
rect 4160 32370 4212 32376
rect 4068 32360 4120 32366
rect 3712 32286 3832 32314
rect 4066 32328 4068 32337
rect 4120 32328 4122 32337
rect 3712 31328 3740 32286
rect 4066 32263 4122 32272
rect 4080 32230 4108 32263
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 3917 32124 4225 32133
rect 3917 32122 3923 32124
rect 3979 32122 4003 32124
rect 4059 32122 4083 32124
rect 4139 32122 4163 32124
rect 4219 32122 4225 32124
rect 3979 32070 3981 32122
rect 4161 32070 4163 32122
rect 3917 32068 3923 32070
rect 3979 32068 4003 32070
rect 4059 32068 4083 32070
rect 4139 32068 4163 32070
rect 4219 32068 4225 32070
rect 3917 32059 4225 32068
rect 4264 32008 4292 34360
rect 4342 33416 4398 33425
rect 4342 33351 4344 33360
rect 4396 33351 4398 33360
rect 4344 33322 4396 33328
rect 4172 31980 4292 32008
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3804 31657 3832 31758
rect 3790 31648 3846 31657
rect 3790 31583 3846 31592
rect 4172 31521 4200 31980
rect 4448 31754 4476 34886
rect 4540 33590 4568 35527
rect 4632 35018 4660 36722
rect 4724 36038 4752 36722
rect 4896 36712 4948 36718
rect 4896 36654 4948 36660
rect 4908 36310 4936 36654
rect 4896 36304 4948 36310
rect 4896 36246 4948 36252
rect 4804 36168 4856 36174
rect 4804 36110 4856 36116
rect 4712 36032 4764 36038
rect 4712 35974 4764 35980
rect 4712 35556 4764 35562
rect 4712 35498 4764 35504
rect 4620 35012 4672 35018
rect 4620 34954 4672 34960
rect 4632 34746 4660 34954
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 4528 33584 4580 33590
rect 4528 33526 4580 33532
rect 4620 33516 4672 33522
rect 4620 33458 4672 33464
rect 4528 32836 4580 32842
rect 4528 32778 4580 32784
rect 4540 32745 4568 32778
rect 4526 32736 4582 32745
rect 4526 32671 4582 32680
rect 4540 32570 4568 32671
rect 4528 32564 4580 32570
rect 4528 32506 4580 32512
rect 4632 32434 4660 33458
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4264 31726 4476 31754
rect 4158 31512 4214 31521
rect 4158 31447 4214 31456
rect 4160 31408 4212 31414
rect 4158 31376 4160 31385
rect 4212 31376 4214 31385
rect 3712 31300 3832 31328
rect 4158 31311 4214 31320
rect 3700 31204 3752 31210
rect 3700 31146 3752 31152
rect 3712 30394 3740 31146
rect 3804 30920 3832 31300
rect 3917 31036 4225 31045
rect 3917 31034 3923 31036
rect 3979 31034 4003 31036
rect 4059 31034 4083 31036
rect 4139 31034 4163 31036
rect 4219 31034 4225 31036
rect 3979 30982 3981 31034
rect 4161 30982 4163 31034
rect 3917 30980 3923 30982
rect 3979 30980 4003 30982
rect 4059 30980 4083 30982
rect 4139 30980 4163 30982
rect 4219 30980 4225 30982
rect 3917 30971 4225 30980
rect 4264 30920 4292 31726
rect 4724 31668 4752 35498
rect 3804 30892 3924 30920
rect 3792 30728 3844 30734
rect 3792 30670 3844 30676
rect 3700 30388 3752 30394
rect 3700 30330 3752 30336
rect 3804 30297 3832 30670
rect 3790 30288 3846 30297
rect 3790 30223 3846 30232
rect 3896 30138 3924 30892
rect 3712 30110 3924 30138
rect 4080 30892 4292 30920
rect 4356 31640 4752 31668
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 3620 29345 3648 29582
rect 3606 29336 3662 29345
rect 3606 29271 3662 29280
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3620 28937 3648 29106
rect 3606 28928 3662 28937
rect 3606 28863 3662 28872
rect 3608 28552 3660 28558
rect 3608 28494 3660 28500
rect 3516 28416 3568 28422
rect 3516 28358 3568 28364
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 3528 26586 3556 28018
rect 3620 26994 3648 28494
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 3516 26580 3568 26586
rect 3516 26522 3568 26528
rect 3608 26512 3660 26518
rect 3608 26454 3660 26460
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 3528 25945 3556 26318
rect 3514 25936 3570 25945
rect 3514 25871 3570 25880
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3528 24886 3556 25094
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3528 23866 3556 24686
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3332 23724 3384 23730
rect 3436 23718 3556 23746
rect 3332 23666 3384 23672
rect 3240 23316 3292 23322
rect 3240 23258 3292 23264
rect 3054 23216 3110 23225
rect 3054 23151 3110 23160
rect 3068 22234 3096 23151
rect 3344 23118 3372 23666
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3238 22128 3294 22137
rect 3238 22063 3294 22072
rect 3252 22030 3280 22063
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3160 21894 3188 21966
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 2964 21072 3016 21078
rect 2964 21014 3016 21020
rect 3344 20874 3372 22918
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3148 20392 3200 20398
rect 3436 20380 3464 23598
rect 3528 22778 3556 23718
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3620 22234 3648 26454
rect 3712 24721 3740 30110
rect 4080 30036 4108 30892
rect 4160 30728 4212 30734
rect 4160 30670 4212 30676
rect 4172 30190 4200 30670
rect 4252 30660 4304 30666
rect 4252 30602 4304 30608
rect 4264 30433 4292 30602
rect 4250 30424 4306 30433
rect 4250 30359 4306 30368
rect 4160 30184 4212 30190
rect 4212 30144 4292 30172
rect 4160 30126 4212 30132
rect 3804 30008 4108 30036
rect 3804 28218 3832 30008
rect 3917 29948 4225 29957
rect 3917 29946 3923 29948
rect 3979 29946 4003 29948
rect 4059 29946 4083 29948
rect 4139 29946 4163 29948
rect 4219 29946 4225 29948
rect 3979 29894 3981 29946
rect 4161 29894 4163 29946
rect 3917 29892 3923 29894
rect 3979 29892 4003 29894
rect 4059 29892 4083 29894
rect 4139 29892 4163 29894
rect 4219 29892 4225 29894
rect 3917 29883 4225 29892
rect 3882 29744 3938 29753
rect 3882 29679 3938 29688
rect 3896 28994 3924 29679
rect 4264 29170 4292 30144
rect 4252 29164 4304 29170
rect 4252 29106 4304 29112
rect 3896 28966 4292 28994
rect 3917 28860 4225 28869
rect 3917 28858 3923 28860
rect 3979 28858 4003 28860
rect 4059 28858 4083 28860
rect 4139 28858 4163 28860
rect 4219 28858 4225 28860
rect 3979 28806 3981 28858
rect 4161 28806 4163 28858
rect 3917 28804 3923 28806
rect 3979 28804 4003 28806
rect 4059 28804 4083 28806
rect 4139 28804 4163 28806
rect 4219 28804 4225 28806
rect 3917 28795 4225 28804
rect 3882 28248 3938 28257
rect 3792 28212 3844 28218
rect 3882 28183 3884 28192
rect 3792 28154 3844 28160
rect 3936 28183 3938 28192
rect 3884 28154 3936 28160
rect 3804 27674 3832 28154
rect 3917 27772 4225 27781
rect 3917 27770 3923 27772
rect 3979 27770 4003 27772
rect 4059 27770 4083 27772
rect 4139 27770 4163 27772
rect 4219 27770 4225 27772
rect 3979 27718 3981 27770
rect 4161 27718 4163 27770
rect 3917 27716 3923 27718
rect 3979 27716 4003 27718
rect 4059 27716 4083 27718
rect 4139 27716 4163 27718
rect 4219 27716 4225 27718
rect 3917 27707 4225 27716
rect 3792 27668 3844 27674
rect 3792 27610 3844 27616
rect 3792 27328 3844 27334
rect 3792 27270 3844 27276
rect 3804 25158 3832 27270
rect 3917 26684 4225 26693
rect 3917 26682 3923 26684
rect 3979 26682 4003 26684
rect 4059 26682 4083 26684
rect 4139 26682 4163 26684
rect 4219 26682 4225 26684
rect 3979 26630 3981 26682
rect 4161 26630 4163 26682
rect 3917 26628 3923 26630
rect 3979 26628 4003 26630
rect 4059 26628 4083 26630
rect 4139 26628 4163 26630
rect 4219 26628 4225 26630
rect 3917 26619 4225 26628
rect 4068 26376 4120 26382
rect 4068 26318 4120 26324
rect 3976 25968 4028 25974
rect 3974 25936 3976 25945
rect 4028 25936 4030 25945
rect 3974 25871 4030 25880
rect 4080 25809 4108 26318
rect 4066 25800 4122 25809
rect 4066 25735 4122 25744
rect 4264 25702 4292 28966
rect 4356 28422 4384 31640
rect 4618 31512 4674 31521
rect 4540 31470 4618 31498
rect 4540 30734 4568 31470
rect 4618 31447 4674 31456
rect 4620 31408 4672 31414
rect 4620 31350 4672 31356
rect 4632 30938 4660 31350
rect 4620 30932 4672 30938
rect 4620 30874 4672 30880
rect 4528 30728 4580 30734
rect 4448 30688 4528 30716
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4356 28150 4384 28358
rect 4344 28144 4396 28150
rect 4344 28086 4396 28092
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 3917 25596 4225 25605
rect 3917 25594 3923 25596
rect 3979 25594 4003 25596
rect 4059 25594 4083 25596
rect 4139 25594 4163 25596
rect 4219 25594 4225 25596
rect 3979 25542 3981 25594
rect 4161 25542 4163 25594
rect 3917 25540 3923 25542
rect 3979 25540 4003 25542
rect 4059 25540 4083 25542
rect 4139 25540 4163 25542
rect 4219 25540 4225 25542
rect 3917 25531 4225 25540
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3988 24818 4016 25094
rect 3792 24812 3844 24818
rect 3792 24754 3844 24760
rect 3976 24812 4028 24818
rect 3976 24754 4028 24760
rect 3698 24712 3754 24721
rect 3698 24647 3754 24656
rect 3804 23848 3832 24754
rect 4080 24750 4108 25230
rect 4160 25152 4212 25158
rect 4160 25094 4212 25100
rect 4172 24954 4200 25094
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4158 24848 4214 24857
rect 4158 24783 4214 24792
rect 4068 24744 4120 24750
rect 4068 24686 4120 24692
rect 4172 24682 4200 24783
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 4252 24676 4304 24682
rect 4252 24618 4304 24624
rect 3917 24508 4225 24517
rect 3917 24506 3923 24508
rect 3979 24506 4003 24508
rect 4059 24506 4083 24508
rect 4139 24506 4163 24508
rect 4219 24506 4225 24508
rect 3979 24454 3981 24506
rect 4161 24454 4163 24506
rect 3917 24452 3923 24454
rect 3979 24452 4003 24454
rect 4059 24452 4083 24454
rect 4139 24452 4163 24454
rect 4219 24452 4225 24454
rect 3917 24443 4225 24452
rect 4264 24274 4292 24618
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4066 23896 4122 23905
rect 3804 23820 3924 23848
rect 4066 23831 4068 23840
rect 3792 23724 3844 23730
rect 3896 23712 3924 23820
rect 4120 23831 4122 23840
rect 4068 23802 4120 23808
rect 3976 23724 4028 23730
rect 3896 23684 3976 23712
rect 3792 23666 3844 23672
rect 3976 23666 4028 23672
rect 3700 23588 3752 23594
rect 3700 23530 3752 23536
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3712 22094 3740 23530
rect 3804 23225 3832 23666
rect 3917 23420 4225 23429
rect 3917 23418 3923 23420
rect 3979 23418 4003 23420
rect 4059 23418 4083 23420
rect 4139 23418 4163 23420
rect 4219 23418 4225 23420
rect 3979 23366 3981 23418
rect 4161 23366 4163 23418
rect 3917 23364 3923 23366
rect 3979 23364 4003 23366
rect 4059 23364 4083 23366
rect 4139 23364 4163 23366
rect 4219 23364 4225 23366
rect 3917 23355 4225 23364
rect 3790 23216 3846 23225
rect 3790 23151 3846 23160
rect 4160 23112 4212 23118
rect 4080 23060 4160 23066
rect 4080 23054 4212 23060
rect 4080 23038 4200 23054
rect 4080 22506 4108 23038
rect 4252 22976 4304 22982
rect 4252 22918 4304 22924
rect 4068 22500 4120 22506
rect 4068 22442 4120 22448
rect 3917 22332 4225 22341
rect 3917 22330 3923 22332
rect 3979 22330 4003 22332
rect 4059 22330 4083 22332
rect 4139 22330 4163 22332
rect 4219 22330 4225 22332
rect 3979 22278 3981 22330
rect 4161 22278 4163 22330
rect 3917 22276 3923 22278
rect 3979 22276 4003 22278
rect 4059 22276 4083 22278
rect 4139 22276 4163 22278
rect 4219 22276 4225 22278
rect 3917 22267 4225 22276
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3200 20352 3464 20380
rect 3620 22066 3740 22094
rect 3148 20334 3200 20340
rect 2870 19816 2926 19825
rect 2870 19751 2926 19760
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2596 17128 2648 17134
rect 2700 17116 2728 17614
rect 2648 17088 2728 17116
rect 2596 17070 2648 17076
rect 2700 16998 2728 17088
rect 2374 16918 2544 16946
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2318 16895 2374 16904
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2410 16552 2466 16561
rect 2228 16516 2280 16522
rect 2410 16487 2466 16496
rect 2228 16458 2280 16464
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 2240 15162 2268 16458
rect 2424 15502 2452 16487
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2332 15065 2360 15302
rect 2318 15056 2374 15065
rect 1768 15020 1820 15026
rect 2318 14991 2374 15000
rect 1768 14962 1820 14968
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 1674 13968 1730 13977
rect 1780 13954 1808 14962
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 1860 14408 1912 14414
rect 1858 14376 1860 14385
rect 1952 14408 2004 14414
rect 1912 14376 1914 14385
rect 2004 14368 2084 14396
rect 1952 14350 2004 14356
rect 1858 14311 1914 14320
rect 1780 13926 1900 13954
rect 1674 13903 1730 13912
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1504 13326 1532 13631
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1214 13152 1270 13161
rect 1214 13087 1270 13096
rect 1582 12608 1638 12617
rect 1582 12543 1638 12552
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1412 10554 1440 11999
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1504 10742 1532 11494
rect 1596 10810 1624 12543
rect 1688 11286 1716 13903
rect 1766 13832 1822 13841
rect 1766 13767 1822 13776
rect 1780 12986 1808 13767
rect 1872 13025 1900 13926
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1858 13016 1914 13025
rect 1768 12980 1820 12986
rect 1858 12951 1914 12960
rect 1768 12922 1820 12928
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 11694 1808 12718
rect 1964 12102 1992 13670
rect 2056 12306 2084 14368
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2148 13394 2176 13874
rect 2332 13734 2360 14758
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2134 12880 2190 12889
rect 2134 12815 2190 12824
rect 2228 12844 2280 12850
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2056 11830 2084 12242
rect 2044 11824 2096 11830
rect 2044 11766 2096 11772
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1492 10736 1544 10742
rect 1492 10678 1544 10684
rect 1780 10606 1808 11630
rect 1950 11520 2006 11529
rect 1950 11455 2006 11464
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1768 10600 1820 10606
rect 1320 9586 1348 10542
rect 1412 10526 1532 10554
rect 1768 10542 1820 10548
rect 1398 9888 1454 9897
rect 1398 9823 1454 9832
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1214 9072 1270 9081
rect 1214 9007 1270 9016
rect 1228 8634 1256 9007
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 1320 8537 1348 9114
rect 1306 8528 1362 8537
rect 1306 8463 1362 8472
rect 1412 8090 1440 9823
rect 1504 9110 1532 10526
rect 1674 10432 1730 10441
rect 1674 10367 1730 10376
rect 1582 9616 1638 9625
rect 1582 9551 1584 9560
rect 1636 9551 1638 9560
rect 1584 9522 1636 9528
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1504 8566 1532 8871
rect 1492 8560 1544 8566
rect 1492 8502 1544 8508
rect 1596 8344 1624 9386
rect 1688 8566 1716 10367
rect 1872 8906 1900 11222
rect 1964 10690 1992 11455
rect 2148 11354 2176 12815
rect 2228 12786 2280 12792
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2044 11076 2096 11082
rect 2240 11064 2268 12786
rect 2332 12782 2360 13670
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2424 11898 2452 12242
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2516 11150 2544 14214
rect 2608 13258 2636 16934
rect 2700 14414 2728 16934
rect 2792 16114 2820 17614
rect 2884 17202 2912 18566
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2976 17678 3004 18022
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2870 16688 2926 16697
rect 3160 16658 3188 20334
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 20058 3556 20266
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3344 19145 3372 19314
rect 3330 19136 3386 19145
rect 3330 19071 3386 19080
rect 3620 17785 3648 22066
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3712 20448 3740 21286
rect 3804 20754 3832 22170
rect 4158 21992 4214 22001
rect 3976 21956 4028 21962
rect 4158 21927 4214 21936
rect 3976 21898 4028 21904
rect 3988 21622 4016 21898
rect 4172 21690 4200 21927
rect 4160 21684 4212 21690
rect 4160 21626 4212 21632
rect 3976 21616 4028 21622
rect 3976 21558 4028 21564
rect 3917 21244 4225 21253
rect 3917 21242 3923 21244
rect 3979 21242 4003 21244
rect 4059 21242 4083 21244
rect 4139 21242 4163 21244
rect 4219 21242 4225 21244
rect 3979 21190 3981 21242
rect 4161 21190 4163 21242
rect 3917 21188 3923 21190
rect 3979 21188 4003 21190
rect 4059 21188 4083 21190
rect 4139 21188 4163 21190
rect 4219 21188 4225 21190
rect 3917 21179 4225 21188
rect 3974 21040 4030 21049
rect 3974 20975 4030 20984
rect 3988 20942 4016 20975
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4068 20800 4120 20806
rect 3804 20726 4016 20754
rect 4068 20742 4120 20748
rect 3988 20602 4016 20726
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3882 20496 3938 20505
rect 3792 20460 3844 20466
rect 3712 20420 3792 20448
rect 4080 20466 4108 20742
rect 3882 20431 3884 20440
rect 3792 20402 3844 20408
rect 3936 20431 3938 20440
rect 4068 20460 4120 20466
rect 3884 20402 3936 20408
rect 4068 20402 4120 20408
rect 3804 19378 3832 20402
rect 3917 20156 4225 20165
rect 3917 20154 3923 20156
rect 3979 20154 4003 20156
rect 4059 20154 4083 20156
rect 4139 20154 4163 20156
rect 4219 20154 4225 20156
rect 3979 20102 3981 20154
rect 4161 20102 4163 20154
rect 3917 20100 3923 20102
rect 3979 20100 4003 20102
rect 4059 20100 4083 20102
rect 4139 20100 4163 20102
rect 4219 20100 4225 20102
rect 3917 20091 4225 20100
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3790 19272 3846 19281
rect 3790 19207 3846 19216
rect 3606 17776 3662 17785
rect 3804 17746 3832 19207
rect 3917 19068 4225 19077
rect 3917 19066 3923 19068
rect 3979 19066 4003 19068
rect 4059 19066 4083 19068
rect 4139 19066 4163 19068
rect 4219 19066 4225 19068
rect 3979 19014 3981 19066
rect 4161 19014 4163 19066
rect 3917 19012 3923 19014
rect 3979 19012 4003 19014
rect 4059 19012 4083 19014
rect 4139 19012 4163 19014
rect 4219 19012 4225 19014
rect 3917 19003 4225 19012
rect 3974 18864 4030 18873
rect 3974 18799 4030 18808
rect 3988 18766 4016 18799
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 18442 4108 18566
rect 4158 18456 4214 18465
rect 4080 18414 4158 18442
rect 4080 18358 4108 18414
rect 4158 18391 4214 18400
rect 4068 18352 4120 18358
rect 4068 18294 4120 18300
rect 4158 18320 4214 18329
rect 4158 18255 4160 18264
rect 4212 18255 4214 18264
rect 4160 18226 4212 18232
rect 3917 17980 4225 17989
rect 3917 17978 3923 17980
rect 3979 17978 4003 17980
rect 4059 17978 4083 17980
rect 4139 17978 4163 17980
rect 4219 17978 4225 17980
rect 3979 17926 3981 17978
rect 4161 17926 4163 17978
rect 3917 17924 3923 17926
rect 3979 17924 4003 17926
rect 4059 17924 4083 17926
rect 4139 17924 4163 17926
rect 4219 17924 4225 17926
rect 3917 17915 4225 17924
rect 3606 17711 3662 17720
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3252 16726 3280 17478
rect 3436 17354 3464 17478
rect 3344 17338 3464 17354
rect 3332 17332 3464 17338
rect 3384 17326 3464 17332
rect 3332 17274 3384 17280
rect 3424 17264 3476 17270
rect 3424 17206 3476 17212
rect 3240 16720 3292 16726
rect 3240 16662 3292 16668
rect 2870 16623 2926 16632
rect 3148 16652 3200 16658
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2884 15706 2912 16623
rect 3148 16594 3200 16600
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 3068 16153 3096 16390
rect 3330 16280 3386 16289
rect 3330 16215 3386 16224
rect 3344 16182 3372 16215
rect 3332 16176 3384 16182
rect 3054 16144 3110 16153
rect 3332 16118 3384 16124
rect 3054 16079 3110 16088
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2792 14890 2820 15642
rect 3054 15600 3110 15609
rect 3054 15535 3110 15544
rect 3068 15162 3096 15535
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3252 15094 3280 15302
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2872 14816 2924 14822
rect 2778 14784 2834 14793
rect 2872 14758 2924 14764
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 2778 14719 2834 14728
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2700 12238 2728 14350
rect 2792 13190 2820 14719
rect 2884 14618 2912 14758
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2780 12300 2832 12306
rect 2884 12288 2912 14418
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 14074 3004 14350
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3148 13252 3200 13258
rect 3148 13194 3200 13200
rect 2832 12260 2912 12288
rect 2780 12242 2832 12248
rect 2688 12232 2740 12238
rect 2884 12209 2912 12260
rect 2688 12174 2740 12180
rect 2870 12200 2926 12209
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 2596 11076 2648 11082
rect 2240 11036 2360 11064
rect 2044 11018 2096 11024
rect 2056 10810 2084 11018
rect 2226 10976 2282 10985
rect 2226 10911 2282 10920
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 1964 10662 2084 10690
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 8974 1992 10406
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1766 8800 1822 8809
rect 2056 8786 2084 10662
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10266 2176 10610
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2134 10160 2190 10169
rect 2134 10095 2136 10104
rect 2188 10095 2190 10104
rect 2136 10066 2188 10072
rect 1766 8735 1822 8744
rect 1872 8758 2084 8786
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1504 8316 1624 8344
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1504 7936 1532 8316
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1320 7908 1532 7936
rect 1124 7540 1176 7546
rect 952 2310 980 7534
rect 1124 7482 1176 7488
rect 1320 6984 1348 7908
rect 1492 7812 1544 7818
rect 1492 7754 1544 7760
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1136 6956 1348 6984
rect 1030 6624 1086 6633
rect 1030 6559 1086 6568
rect 1044 5846 1072 6559
rect 1032 5840 1084 5846
rect 1032 5782 1084 5788
rect 1136 5234 1164 6956
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6390 1256 6831
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1216 6384 1268 6390
rect 1320 6361 1348 6394
rect 1216 6326 1268 6332
rect 1306 6352 1362 6361
rect 1306 6287 1362 6296
rect 1308 6180 1360 6186
rect 1308 6122 1360 6128
rect 1320 5817 1348 6122
rect 1412 5914 1440 7647
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1306 5808 1362 5817
rect 1306 5743 1362 5752
rect 1124 5228 1176 5234
rect 1124 5170 1176 5176
rect 1504 4826 1532 7754
rect 1596 7002 1624 8191
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7478 1716 7754
rect 1780 7546 1808 8735
rect 1872 8498 1900 8758
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1766 7440 1822 7449
rect 1766 7375 1822 7384
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1780 6118 1808 7375
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1596 3738 1624 5607
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1032 3052 1084 3058
rect 1032 2994 1084 3000
rect 940 2304 992 2310
rect 940 2246 992 2252
rect 846 1456 902 1465
rect 572 1420 624 1426
rect 846 1391 902 1400
rect 572 1362 624 1368
rect 940 1012 992 1018
rect 940 954 992 960
rect 202 0 258 160
rect 478 0 534 160
rect 754 82 810 160
rect 952 82 980 954
rect 1044 160 1072 2994
rect 1688 2378 1716 4966
rect 1872 4298 1900 8026
rect 2148 7274 2176 10066
rect 2240 9110 2268 10911
rect 2332 9761 2360 11036
rect 2596 11018 2648 11024
rect 2608 10180 2636 11018
rect 2514 10152 2636 10180
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2318 9752 2374 9761
rect 2424 9722 2452 10066
rect 2514 9908 2542 10152
rect 2700 10130 2728 12174
rect 2870 12135 2926 12144
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3068 11665 3096 11766
rect 3054 11656 3110 11665
rect 3054 11591 3110 11600
rect 3056 11348 3108 11354
rect 3056 11290 3108 11296
rect 2964 10464 3016 10470
rect 2884 10424 2964 10452
rect 2884 10248 2912 10424
rect 2964 10406 3016 10412
rect 3068 10305 3096 11290
rect 3160 10554 3188 13194
rect 3252 12850 3280 14758
rect 3330 14512 3386 14521
rect 3330 14447 3386 14456
rect 3344 14074 3372 14447
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3344 13326 3372 13670
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3252 12481 3280 12650
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3238 12472 3294 12481
rect 3238 12407 3294 12416
rect 3344 12306 3372 12582
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 3436 11880 3464 17206
rect 3528 16794 3556 17546
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 15910 3556 16526
rect 3620 16046 3648 17614
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3620 14498 3648 15982
rect 3712 15638 3740 17002
rect 3804 16794 3832 17138
rect 3917 16892 4225 16901
rect 3917 16890 3923 16892
rect 3979 16890 4003 16892
rect 4059 16890 4083 16892
rect 4139 16890 4163 16892
rect 4219 16890 4225 16892
rect 3979 16838 3981 16890
rect 4161 16838 4163 16890
rect 3917 16836 3923 16838
rect 3979 16836 4003 16838
rect 4059 16836 4083 16838
rect 4139 16836 4163 16838
rect 4219 16836 4225 16838
rect 3917 16827 4225 16836
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3976 16448 4028 16454
rect 3974 16416 3976 16425
rect 4028 16416 4030 16425
rect 3974 16351 4030 16360
rect 3917 15804 4225 15813
rect 3917 15802 3923 15804
rect 3979 15802 4003 15804
rect 4059 15802 4083 15804
rect 4139 15802 4163 15804
rect 4219 15802 4225 15804
rect 3979 15750 3981 15802
rect 4161 15750 4163 15802
rect 3917 15748 3923 15750
rect 3979 15748 4003 15750
rect 4059 15748 4083 15750
rect 4139 15748 4163 15750
rect 4219 15748 4225 15750
rect 3917 15739 4225 15748
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3974 15600 4030 15609
rect 4158 15600 4214 15609
rect 3974 15535 4030 15544
rect 4080 15558 4158 15586
rect 3700 15496 3752 15502
rect 3700 15438 3752 15444
rect 3712 14929 3740 15438
rect 3988 15162 4016 15535
rect 4080 15502 4108 15558
rect 4158 15535 4214 15544
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 15162 4200 15438
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4264 15026 4292 22918
rect 4356 21350 4384 26386
rect 4448 25906 4476 30688
rect 4528 30670 4580 30676
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4528 30592 4580 30598
rect 4528 30534 4580 30540
rect 4540 28150 4568 30534
rect 4528 28144 4580 28150
rect 4528 28086 4580 28092
rect 4540 27334 4568 28086
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4528 26988 4580 26994
rect 4528 26930 4580 26936
rect 4540 26518 4568 26930
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4436 25900 4488 25906
rect 4436 25842 4488 25848
rect 4436 25696 4488 25702
rect 4436 25638 4488 25644
rect 4448 25294 4476 25638
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4540 24818 4568 25230
rect 4632 25226 4660 30670
rect 4712 30320 4764 30326
rect 4712 30262 4764 30268
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4528 24812 4580 24818
rect 4528 24754 4580 24760
rect 4436 24744 4488 24750
rect 4436 24686 4488 24692
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4342 21040 4398 21049
rect 4342 20975 4398 20984
rect 4356 20058 4384 20975
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4356 17134 4384 18226
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4356 16096 4384 17070
rect 4448 16776 4476 24686
rect 4540 21418 4568 24754
rect 4632 24138 4660 25162
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4620 21888 4672 21894
rect 4618 21856 4620 21865
rect 4672 21856 4674 21865
rect 4618 21791 4674 21800
rect 4724 21672 4752 30262
rect 4816 28150 4844 36110
rect 4908 34785 4936 36246
rect 4894 34776 4950 34785
rect 4894 34711 4950 34720
rect 4896 33924 4948 33930
rect 4896 33866 4948 33872
rect 4908 33522 4936 33866
rect 4896 33516 4948 33522
rect 4896 33458 4948 33464
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4908 32434 4936 32710
rect 4896 32428 4948 32434
rect 4896 32370 4948 32376
rect 4908 31906 4936 32370
rect 5000 32366 5028 37198
rect 4988 32360 5040 32366
rect 4988 32302 5040 32308
rect 5092 32026 5120 40326
rect 5172 40180 5224 40186
rect 5172 40122 5224 40128
rect 5184 39386 5212 40122
rect 5276 39506 5304 43658
rect 5552 43450 5580 43846
rect 5540 43444 5592 43450
rect 5540 43386 5592 43392
rect 5448 43308 5500 43314
rect 5448 43250 5500 43256
rect 5540 43308 5592 43314
rect 5540 43250 5592 43256
rect 5460 42294 5488 43250
rect 5448 42288 5500 42294
rect 5448 42230 5500 42236
rect 5552 41818 5580 43250
rect 5736 42566 5764 44463
rect 6012 43602 6040 44463
rect 6012 43574 6132 43602
rect 6104 42906 6132 43574
rect 6288 43450 6316 44463
rect 6276 43444 6328 43450
rect 6276 43386 6328 43392
rect 6564 43330 6592 44463
rect 6840 43874 6868 44463
rect 6656 43846 6868 43874
rect 7116 43874 7144 44463
rect 7392 44010 7420 44463
rect 7392 43982 7512 44010
rect 7116 43846 7420 43874
rect 6656 43450 6684 43846
rect 6884 43548 7192 43557
rect 6884 43546 6890 43548
rect 6946 43546 6970 43548
rect 7026 43546 7050 43548
rect 7106 43546 7130 43548
rect 7186 43546 7192 43548
rect 6946 43494 6948 43546
rect 7128 43494 7130 43546
rect 6884 43492 6890 43494
rect 6946 43492 6970 43494
rect 7026 43492 7050 43494
rect 7106 43492 7130 43494
rect 7186 43492 7192 43494
rect 6884 43483 7192 43492
rect 6644 43444 6696 43450
rect 6644 43386 6696 43392
rect 6276 43308 6328 43314
rect 6564 43302 6868 43330
rect 6276 43250 6328 43256
rect 6092 42900 6144 42906
rect 6092 42842 6144 42848
rect 6000 42628 6052 42634
rect 6000 42570 6052 42576
rect 5724 42560 5776 42566
rect 5724 42502 5776 42508
rect 5908 42560 5960 42566
rect 5908 42502 5960 42508
rect 5814 42392 5870 42401
rect 5920 42362 5948 42502
rect 5814 42327 5870 42336
rect 5908 42356 5960 42362
rect 5828 42294 5856 42327
rect 5908 42298 5960 42304
rect 5816 42288 5868 42294
rect 5816 42230 5868 42236
rect 5816 42084 5868 42090
rect 5816 42026 5868 42032
rect 5540 41812 5592 41818
rect 5540 41754 5592 41760
rect 5828 41614 5856 42026
rect 6012 41818 6040 42570
rect 6288 42362 6316 43250
rect 6840 42906 6868 43302
rect 7288 43308 7340 43314
rect 7288 43250 7340 43256
rect 6828 42900 6880 42906
rect 6828 42842 6880 42848
rect 7300 42786 7328 43250
rect 7392 42906 7420 43846
rect 7380 42900 7432 42906
rect 7380 42842 7432 42848
rect 7300 42758 7420 42786
rect 6736 42628 6788 42634
rect 6736 42570 6788 42576
rect 7288 42628 7340 42634
rect 7288 42570 7340 42576
rect 6276 42356 6328 42362
rect 6276 42298 6328 42304
rect 6276 42152 6328 42158
rect 6276 42094 6328 42100
rect 6288 41857 6316 42094
rect 6274 41848 6330 41857
rect 6000 41812 6052 41818
rect 6748 41818 6776 42570
rect 6884 42460 7192 42469
rect 6884 42458 6890 42460
rect 6946 42458 6970 42460
rect 7026 42458 7050 42460
rect 7106 42458 7130 42460
rect 7186 42458 7192 42460
rect 6946 42406 6948 42458
rect 7128 42406 7130 42458
rect 6884 42404 6890 42406
rect 6946 42404 6970 42406
rect 7026 42404 7050 42406
rect 7106 42404 7130 42406
rect 7186 42404 7192 42406
rect 6884 42395 7192 42404
rect 7196 42356 7248 42362
rect 7196 42298 7248 42304
rect 6920 42152 6972 42158
rect 6920 42094 6972 42100
rect 7102 42120 7158 42129
rect 6274 41783 6330 41792
rect 6736 41812 6788 41818
rect 6000 41754 6052 41760
rect 6736 41754 6788 41760
rect 5356 41608 5408 41614
rect 5356 41550 5408 41556
rect 5816 41608 5868 41614
rect 5816 41550 5868 41556
rect 5368 40225 5396 41550
rect 6092 41472 6144 41478
rect 6932 41460 6960 42094
rect 7102 42055 7158 42064
rect 7116 42022 7144 42055
rect 7104 42016 7156 42022
rect 7104 41958 7156 41964
rect 7208 41478 7236 42298
rect 7300 41818 7328 42570
rect 7392 42362 7420 42758
rect 7484 42566 7512 43982
rect 7668 43450 7696 44463
rect 7944 43450 7972 44463
rect 7656 43444 7708 43450
rect 7656 43386 7708 43392
rect 7932 43444 7984 43450
rect 7932 43386 7984 43392
rect 8116 43240 8168 43246
rect 8116 43182 8168 43188
rect 7748 42696 7800 42702
rect 7748 42638 7800 42644
rect 7472 42560 7524 42566
rect 7472 42502 7524 42508
rect 7380 42356 7432 42362
rect 7380 42298 7432 42304
rect 7472 42220 7524 42226
rect 7472 42162 7524 42168
rect 7656 42220 7708 42226
rect 7656 42162 7708 42168
rect 7380 42016 7432 42022
rect 7380 41958 7432 41964
rect 7392 41818 7420 41958
rect 7484 41857 7512 42162
rect 7564 42084 7616 42090
rect 7564 42026 7616 42032
rect 7470 41848 7526 41857
rect 7288 41812 7340 41818
rect 7288 41754 7340 41760
rect 7380 41812 7432 41818
rect 7470 41783 7526 41792
rect 7380 41754 7432 41760
rect 7576 41682 7604 42026
rect 7564 41676 7616 41682
rect 7564 41618 7616 41624
rect 6092 41414 6144 41420
rect 6748 41432 6960 41460
rect 7196 41472 7248 41478
rect 5540 41200 5592 41206
rect 5540 41142 5592 41148
rect 5552 40594 5580 41142
rect 6000 40928 6052 40934
rect 6000 40870 6052 40876
rect 5630 40624 5686 40633
rect 5540 40588 5592 40594
rect 5592 40568 5630 40576
rect 5592 40559 5686 40568
rect 5592 40548 5672 40559
rect 5540 40530 5592 40536
rect 5448 40520 5500 40526
rect 5448 40462 5500 40468
rect 5354 40216 5410 40225
rect 5460 40186 5488 40462
rect 5354 40151 5410 40160
rect 5448 40180 5500 40186
rect 5448 40122 5500 40128
rect 5552 40118 5580 40530
rect 5540 40112 5592 40118
rect 5540 40054 5592 40060
rect 5264 39500 5316 39506
rect 5264 39442 5316 39448
rect 5184 39358 5304 39386
rect 5172 39296 5224 39302
rect 5172 39238 5224 39244
rect 5184 38350 5212 39238
rect 5172 38344 5224 38350
rect 5172 38286 5224 38292
rect 5184 36174 5212 38286
rect 5276 36825 5304 39358
rect 5552 38654 5580 40054
rect 5908 39840 5960 39846
rect 5908 39782 5960 39788
rect 5920 39642 5948 39782
rect 5908 39636 5960 39642
rect 5908 39578 5960 39584
rect 5552 38626 5764 38654
rect 5356 38548 5408 38554
rect 5356 38490 5408 38496
rect 5368 38350 5396 38490
rect 5356 38344 5408 38350
rect 5356 38286 5408 38292
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 5448 38276 5500 38282
rect 5448 38218 5500 38224
rect 5356 37868 5408 37874
rect 5356 37810 5408 37816
rect 5368 37505 5396 37810
rect 5354 37496 5410 37505
rect 5354 37431 5410 37440
rect 5460 37262 5488 38218
rect 5552 37369 5580 38286
rect 5736 37874 5764 38626
rect 6012 38486 6040 40870
rect 6000 38480 6052 38486
rect 6000 38422 6052 38428
rect 5724 37868 5776 37874
rect 5724 37810 5776 37816
rect 6000 37664 6052 37670
rect 6000 37606 6052 37612
rect 5538 37360 5594 37369
rect 5538 37295 5594 37304
rect 5448 37256 5500 37262
rect 5448 37198 5500 37204
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5262 36816 5318 36825
rect 5262 36751 5318 36760
rect 5172 36168 5224 36174
rect 5448 36168 5500 36174
rect 5172 36110 5224 36116
rect 5446 36136 5448 36145
rect 5500 36136 5502 36145
rect 5446 36071 5502 36080
rect 5172 36032 5224 36038
rect 5172 35974 5224 35980
rect 5354 36000 5410 36009
rect 5184 34950 5212 35974
rect 5354 35935 5410 35944
rect 5264 35624 5316 35630
rect 5264 35566 5316 35572
rect 5276 35154 5304 35566
rect 5264 35148 5316 35154
rect 5264 35090 5316 35096
rect 5276 35018 5304 35090
rect 5264 35012 5316 35018
rect 5264 34954 5316 34960
rect 5172 34944 5224 34950
rect 5172 34886 5224 34892
rect 5170 34640 5226 34649
rect 5226 34598 5304 34626
rect 5170 34575 5226 34584
rect 5172 34400 5224 34406
rect 5172 34342 5224 34348
rect 5184 33658 5212 34342
rect 5276 33998 5304 34598
rect 5368 34513 5396 35935
rect 5448 35624 5500 35630
rect 5448 35566 5500 35572
rect 5354 34504 5410 34513
rect 5354 34439 5410 34448
rect 5264 33992 5316 33998
rect 5264 33934 5316 33940
rect 5172 33652 5224 33658
rect 5172 33594 5224 33600
rect 5368 33590 5396 34439
rect 5356 33584 5408 33590
rect 5356 33526 5408 33532
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 5356 33312 5408 33318
rect 5356 33254 5408 33260
rect 5184 32570 5212 33254
rect 5262 33008 5318 33017
rect 5262 32943 5318 32952
rect 5276 32910 5304 32943
rect 5368 32910 5396 33254
rect 5460 32910 5488 35566
rect 5552 35290 5580 37130
rect 5724 37120 5776 37126
rect 5724 37062 5776 37068
rect 5632 36576 5684 36582
rect 5632 36518 5684 36524
rect 5644 36038 5672 36518
rect 5736 36310 5764 37062
rect 5816 36848 5868 36854
rect 5816 36790 5868 36796
rect 5724 36304 5776 36310
rect 5724 36246 5776 36252
rect 5632 36032 5684 36038
rect 5632 35974 5684 35980
rect 5540 35284 5592 35290
rect 5540 35226 5592 35232
rect 5540 34604 5592 34610
rect 5540 34546 5592 34552
rect 5552 34202 5580 34546
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5552 32978 5580 33798
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5264 32904 5316 32910
rect 5264 32846 5316 32852
rect 5356 32904 5408 32910
rect 5356 32846 5408 32852
rect 5448 32904 5500 32910
rect 5448 32846 5500 32852
rect 5460 32722 5488 32846
rect 5276 32694 5488 32722
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5172 32360 5224 32366
rect 5172 32302 5224 32308
rect 5080 32020 5132 32026
rect 5080 31962 5132 31968
rect 4908 31878 5120 31906
rect 4896 31816 4948 31822
rect 4948 31776 5028 31804
rect 4896 31758 4948 31764
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4908 30841 4936 31282
rect 5000 31249 5028 31776
rect 4986 31240 5042 31249
rect 4986 31175 5042 31184
rect 4894 30832 4950 30841
rect 4894 30767 4950 30776
rect 5092 30734 5120 31878
rect 5080 30728 5132 30734
rect 5080 30670 5132 30676
rect 5184 30274 5212 32302
rect 5276 30598 5304 32694
rect 5644 32586 5672 35974
rect 5736 35494 5764 36246
rect 5724 35488 5776 35494
rect 5724 35430 5776 35436
rect 5724 35080 5776 35086
rect 5724 35022 5776 35028
rect 5356 32564 5408 32570
rect 5356 32506 5408 32512
rect 5460 32558 5672 32586
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 4908 30246 5212 30274
rect 5262 30288 5318 30297
rect 4908 28744 4936 30246
rect 5262 30223 5318 30232
rect 5080 30184 5132 30190
rect 5080 30126 5132 30132
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 5000 29209 5028 29446
rect 5092 29288 5120 30126
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5184 29714 5212 29990
rect 5172 29708 5224 29714
rect 5172 29650 5224 29656
rect 5276 29578 5304 30223
rect 5368 30036 5396 32506
rect 5460 30190 5488 32558
rect 5630 32328 5686 32337
rect 5630 32263 5686 32272
rect 5540 31816 5592 31822
rect 5540 31758 5592 31764
rect 5552 30190 5580 31758
rect 5644 31482 5672 32263
rect 5736 32230 5764 35022
rect 5828 34950 5856 36790
rect 6012 36394 6040 37606
rect 6104 36553 6132 41414
rect 6748 41256 6776 41432
rect 7196 41414 7248 41420
rect 7668 41414 7696 42162
rect 7760 41818 7788 42638
rect 7840 42152 7892 42158
rect 7840 42094 7892 42100
rect 7748 41812 7800 41818
rect 7748 41754 7800 41760
rect 7484 41386 7696 41414
rect 6884 41372 7192 41381
rect 6884 41370 6890 41372
rect 6946 41370 6970 41372
rect 7026 41370 7050 41372
rect 7106 41370 7130 41372
rect 7186 41370 7192 41372
rect 6946 41318 6948 41370
rect 7128 41318 7130 41370
rect 6884 41316 6890 41318
rect 6946 41316 6970 41318
rect 7026 41316 7050 41318
rect 7106 41316 7130 41318
rect 7186 41316 7192 41318
rect 6884 41307 7192 41316
rect 6748 41228 6960 41256
rect 6932 41002 6960 41228
rect 6920 40996 6972 41002
rect 6920 40938 6972 40944
rect 7484 40934 7512 41386
rect 7852 41274 7880 42094
rect 7932 42016 7984 42022
rect 7932 41958 7984 41964
rect 8024 42016 8076 42022
rect 8024 41958 8076 41964
rect 7944 41818 7972 41958
rect 7932 41812 7984 41818
rect 7932 41754 7984 41760
rect 8036 41414 8064 41958
rect 8128 41818 8156 43182
rect 8220 42362 8248 44463
rect 8496 43450 8524 44463
rect 8484 43444 8536 43450
rect 8484 43386 8536 43392
rect 8392 42832 8444 42838
rect 8392 42774 8444 42780
rect 8208 42356 8260 42362
rect 8208 42298 8260 42304
rect 8208 42220 8260 42226
rect 8208 42162 8260 42168
rect 8220 41857 8248 42162
rect 8206 41848 8262 41857
rect 8116 41812 8168 41818
rect 8404 41818 8432 42774
rect 8772 42770 8800 44463
rect 9048 43450 9076 44463
rect 9036 43444 9088 43450
rect 9036 43386 9088 43392
rect 8944 43376 8996 43382
rect 8944 43318 8996 43324
rect 8760 42764 8812 42770
rect 8760 42706 8812 42712
rect 8850 42664 8906 42673
rect 8760 42628 8812 42634
rect 8850 42599 8906 42608
rect 8760 42570 8812 42576
rect 8668 42560 8720 42566
rect 8668 42502 8720 42508
rect 8576 42288 8628 42294
rect 8576 42230 8628 42236
rect 8206 41783 8262 41792
rect 8392 41812 8444 41818
rect 8116 41754 8168 41760
rect 8392 41754 8444 41760
rect 8588 41698 8616 42230
rect 7944 41386 8064 41414
rect 8128 41670 8616 41698
rect 8680 41698 8708 42502
rect 8772 42158 8800 42570
rect 8864 42226 8892 42599
rect 8852 42220 8904 42226
rect 8852 42162 8904 42168
rect 8760 42152 8812 42158
rect 8760 42094 8812 42100
rect 8852 42016 8904 42022
rect 8852 41958 8904 41964
rect 8864 41818 8892 41958
rect 8956 41818 8984 43318
rect 9324 42770 9352 44463
rect 9600 43450 9628 44463
rect 9876 43450 9904 44463
rect 9588 43444 9640 43450
rect 9588 43386 9640 43392
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9404 43376 9456 43382
rect 9404 43318 9456 43324
rect 9312 42764 9364 42770
rect 9312 42706 9364 42712
rect 9128 42696 9180 42702
rect 9128 42638 9180 42644
rect 9140 42294 9168 42638
rect 9312 42560 9364 42566
rect 9312 42502 9364 42508
rect 9128 42288 9180 42294
rect 9128 42230 9180 42236
rect 9036 42220 9088 42226
rect 9036 42162 9088 42168
rect 9048 41818 9076 42162
rect 8852 41812 8904 41818
rect 8852 41754 8904 41760
rect 8944 41812 8996 41818
rect 8944 41754 8996 41760
rect 9036 41812 9088 41818
rect 9036 41754 9088 41760
rect 9324 41698 9352 42502
rect 8680 41670 8892 41698
rect 7564 41268 7616 41274
rect 7564 41210 7616 41216
rect 7840 41268 7892 41274
rect 7840 41210 7892 41216
rect 7380 40928 7432 40934
rect 7380 40870 7432 40876
rect 7472 40928 7524 40934
rect 7472 40870 7524 40876
rect 7286 40488 7342 40497
rect 6736 40452 6788 40458
rect 7286 40423 7342 40432
rect 6736 40394 6788 40400
rect 6644 40384 6696 40390
rect 6644 40326 6696 40332
rect 6460 40044 6512 40050
rect 6460 39986 6512 39992
rect 6472 39438 6500 39986
rect 6656 39438 6684 40326
rect 6748 39642 6776 40394
rect 6884 40284 7192 40293
rect 6884 40282 6890 40284
rect 6946 40282 6970 40284
rect 7026 40282 7050 40284
rect 7106 40282 7130 40284
rect 7186 40282 7192 40284
rect 6946 40230 6948 40282
rect 7128 40230 7130 40282
rect 6884 40228 6890 40230
rect 6946 40228 6970 40230
rect 7026 40228 7050 40230
rect 7106 40228 7130 40230
rect 7186 40228 7192 40230
rect 6884 40219 7192 40228
rect 7300 40186 7328 40423
rect 7288 40180 7340 40186
rect 7288 40122 7340 40128
rect 6736 39636 6788 39642
rect 6736 39578 6788 39584
rect 6460 39432 6512 39438
rect 6460 39374 6512 39380
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 6276 38344 6328 38350
rect 6276 38286 6328 38292
rect 6184 37800 6236 37806
rect 6184 37742 6236 37748
rect 6196 37466 6224 37742
rect 6288 37738 6316 38286
rect 6368 37800 6420 37806
rect 6368 37742 6420 37748
rect 6276 37732 6328 37738
rect 6276 37674 6328 37680
rect 6184 37460 6236 37466
rect 6184 37402 6236 37408
rect 6090 36544 6146 36553
rect 6090 36479 6146 36488
rect 6012 36366 6132 36394
rect 6104 36174 6132 36366
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 6092 36168 6144 36174
rect 6092 36110 6144 36116
rect 6276 36168 6328 36174
rect 6276 36110 6328 36116
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 5816 34944 5868 34950
rect 5816 34886 5868 34892
rect 5920 34542 5948 35430
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5724 32224 5776 32230
rect 5724 32166 5776 32172
rect 5828 31890 5856 32846
rect 5816 31884 5868 31890
rect 5816 31826 5868 31832
rect 5724 31748 5776 31754
rect 5724 31690 5776 31696
rect 5736 31482 5764 31690
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5724 31476 5776 31482
rect 5724 31418 5776 31424
rect 5632 31340 5684 31346
rect 5632 31282 5684 31288
rect 5448 30184 5500 30190
rect 5448 30126 5500 30132
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 5368 30008 5488 30036
rect 5264 29572 5316 29578
rect 5264 29514 5316 29520
rect 5356 29572 5408 29578
rect 5356 29514 5408 29520
rect 5368 29306 5396 29514
rect 5356 29300 5408 29306
rect 5092 29260 5212 29288
rect 4986 29200 5042 29209
rect 4986 29135 5042 29144
rect 5080 29164 5132 29170
rect 5080 29106 5132 29112
rect 5092 29073 5120 29106
rect 5078 29064 5134 29073
rect 5078 28999 5134 29008
rect 4908 28716 5120 28744
rect 5092 28558 5120 28716
rect 4896 28552 4948 28558
rect 4894 28520 4896 28529
rect 5080 28552 5132 28558
rect 4948 28520 4950 28529
rect 5080 28494 5132 28500
rect 4894 28455 4950 28464
rect 4896 28416 4948 28422
rect 4896 28358 4948 28364
rect 4804 28144 4856 28150
rect 4804 28086 4856 28092
rect 4816 24274 4844 28086
rect 4908 28014 4936 28358
rect 4896 28008 4948 28014
rect 4896 27950 4948 27956
rect 4986 27840 5042 27849
rect 4986 27775 5042 27784
rect 5000 27470 5028 27775
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4896 26988 4948 26994
rect 5092 26976 5120 28494
rect 4948 26948 5120 26976
rect 4896 26930 4948 26936
rect 4908 26382 4936 26930
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4908 24154 4936 25638
rect 4632 21644 4752 21672
rect 4816 24126 4936 24154
rect 4528 21412 4580 21418
rect 4528 21354 4580 21360
rect 4540 18970 4568 21354
rect 4632 21026 4660 21644
rect 4710 21040 4766 21049
rect 4632 20998 4710 21026
rect 4710 20975 4766 20984
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4724 19514 4752 20198
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4632 19378 4660 19450
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4540 17338 4568 18702
rect 4632 17542 4660 18838
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4816 18714 4844 24126
rect 4896 22976 4948 22982
rect 4896 22918 4948 22924
rect 4908 22438 4936 22918
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4908 21554 4936 22374
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 4896 20528 4948 20534
rect 4896 20470 4948 20476
rect 4908 19378 4936 20470
rect 5000 19786 5028 26182
rect 5184 24993 5212 29260
rect 5356 29242 5408 29248
rect 5356 28484 5408 28490
rect 5356 28426 5408 28432
rect 5368 28082 5396 28426
rect 5356 28076 5408 28082
rect 5356 28018 5408 28024
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 5170 24984 5226 24993
rect 5170 24919 5226 24928
rect 5080 24268 5132 24274
rect 5080 24210 5132 24216
rect 5092 24018 5120 24210
rect 5184 24138 5212 24919
rect 5276 24818 5304 27610
rect 5356 27056 5408 27062
rect 5356 26998 5408 27004
rect 5368 26790 5396 26998
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5356 25968 5408 25974
rect 5356 25910 5408 25916
rect 5368 25276 5396 25910
rect 5460 25498 5488 30008
rect 5540 28144 5592 28150
rect 5540 28086 5592 28092
rect 5552 26926 5580 28086
rect 5540 26920 5592 26926
rect 5540 26862 5592 26868
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5448 25492 5500 25498
rect 5448 25434 5500 25440
rect 5448 25288 5500 25294
rect 5368 25248 5448 25276
rect 5448 25230 5500 25236
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5276 24290 5304 24754
rect 5276 24262 5396 24290
rect 5172 24132 5224 24138
rect 5172 24074 5224 24080
rect 5092 23990 5304 24018
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22098 5212 22374
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5080 21956 5132 21962
rect 5132 21916 5212 21944
rect 5080 21898 5132 21904
rect 5184 21690 5212 21916
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5092 20942 5120 21626
rect 5080 20936 5132 20942
rect 5080 20878 5132 20884
rect 4988 19780 5040 19786
rect 4988 19722 5040 19728
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4724 18358 4752 18702
rect 4816 18686 4936 18714
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4712 18352 4764 18358
rect 4712 18294 4764 18300
rect 4816 17882 4844 18566
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4816 17202 4844 17478
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4908 16946 4936 18686
rect 5000 18222 5028 19722
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 17678 5028 18022
rect 5078 17776 5134 17785
rect 5078 17711 5134 17720
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4908 16918 5028 16946
rect 4448 16748 4844 16776
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 4436 16108 4488 16114
rect 4356 16068 4436 16096
rect 4356 15094 4384 16068
rect 4436 16050 4488 16056
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 3698 14920 3754 14929
rect 3698 14855 3754 14864
rect 3804 14618 3832 14962
rect 3917 14716 4225 14725
rect 3917 14714 3923 14716
rect 3979 14714 4003 14716
rect 4059 14714 4083 14716
rect 4139 14714 4163 14716
rect 4219 14714 4225 14716
rect 3979 14662 3981 14714
rect 4161 14662 4163 14714
rect 3917 14660 3923 14662
rect 3979 14660 4003 14662
rect 4059 14660 4083 14662
rect 4139 14660 4163 14662
rect 4219 14660 4225 14662
rect 3917 14651 4225 14660
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 4356 14550 4384 15030
rect 4344 14544 4396 14550
rect 4250 14512 4306 14521
rect 3620 14470 3832 14498
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3344 11852 3464 11880
rect 3238 11792 3294 11801
rect 3238 11727 3294 11736
rect 3252 11286 3280 11727
rect 3344 11642 3372 11852
rect 3422 11792 3478 11801
rect 3422 11727 3424 11736
rect 3476 11727 3478 11736
rect 3424 11698 3476 11704
rect 3344 11614 3464 11642
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3332 11144 3384 11150
rect 3330 11112 3332 11121
rect 3384 11112 3386 11121
rect 3330 11047 3386 11056
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3160 10526 3280 10554
rect 2838 10220 2912 10248
rect 3054 10296 3110 10305
rect 3054 10231 3110 10240
rect 2838 10146 2866 10220
rect 2688 10124 2740 10130
rect 2838 10118 3004 10146
rect 2688 10066 2740 10072
rect 2976 10062 3004 10118
rect 2872 10056 2924 10062
rect 2870 10024 2872 10033
rect 2964 10056 3016 10062
rect 2924 10024 2926 10033
rect 2964 9998 3016 10004
rect 2870 9959 2926 9968
rect 2514 9880 2636 9908
rect 2318 9687 2374 9696
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2318 9344 2374 9353
rect 2318 9279 2374 9288
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 2240 8090 2268 8434
rect 2332 8430 2360 9279
rect 2608 9058 2636 9880
rect 2884 9846 3188 9874
rect 2686 9752 2742 9761
rect 2686 9687 2742 9696
rect 2516 9030 2636 9058
rect 2700 9058 2728 9687
rect 2778 9480 2834 9489
rect 2778 9415 2780 9424
rect 2832 9415 2834 9424
rect 2780 9386 2832 9392
rect 2700 9030 2820 9058
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 8090 2360 8230
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2228 7880 2280 7886
rect 2226 7848 2228 7857
rect 2280 7848 2282 7857
rect 2226 7783 2282 7792
rect 2320 7812 2372 7818
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2134 7168 2190 7177
rect 2134 7103 2190 7112
rect 2148 5914 2176 7103
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2044 5636 2096 5642
rect 2044 5578 2096 5584
rect 1950 5400 2006 5409
rect 1950 5335 2006 5344
rect 1780 4270 1900 4298
rect 1780 3058 1808 4270
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1872 2417 1900 4082
rect 1964 4078 1992 5335
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 2056 3942 2084 5578
rect 2134 4992 2190 5001
rect 2134 4927 2190 4936
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2148 3738 2176 4927
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2056 3194 2084 3402
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2240 2774 2268 7783
rect 2320 7754 2372 7760
rect 2332 6866 2360 7754
rect 2424 7750 2452 8842
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2424 5930 2452 7278
rect 2516 7154 2544 9030
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2608 7546 2636 8842
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2700 7954 2728 8230
rect 2792 8022 2820 9030
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2792 7410 2820 7482
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2516 7126 2728 7154
rect 2594 6624 2650 6633
rect 2594 6559 2650 6568
rect 2332 5902 2452 5930
rect 2332 4690 2360 5902
rect 2608 5114 2636 6559
rect 2424 5086 2636 5114
rect 2424 4826 2452 5086
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2332 4185 2360 4626
rect 2318 4176 2374 4185
rect 2318 4111 2374 4120
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3126 2360 3334
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 1964 2746 2268 2774
rect 1858 2408 1914 2417
rect 1676 2372 1728 2378
rect 1858 2343 1914 2352
rect 1676 2314 1728 2320
rect 1688 1970 1716 2314
rect 1964 2038 1992 2746
rect 2424 2106 2452 4626
rect 2516 4010 2544 4966
rect 2608 4146 2636 5086
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2700 3738 2728 7126
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2884 6610 2912 9846
rect 3160 9761 3188 9846
rect 2962 9752 3018 9761
rect 2962 9687 3018 9696
rect 3146 9752 3202 9761
rect 3146 9687 3202 9696
rect 2976 8922 3004 9687
rect 3148 9648 3200 9654
rect 3148 9590 3200 9596
rect 3160 9450 3188 9590
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9178 3096 9318
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3054 8936 3110 8945
rect 2976 8894 3054 8922
rect 3054 8871 3110 8880
rect 3160 7834 3188 9386
rect 3252 9178 3280 10526
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3344 8480 3372 10950
rect 3436 8974 3464 11614
rect 3528 9654 3556 14214
rect 3698 12880 3754 12889
rect 3608 12844 3660 12850
rect 3698 12815 3754 12824
rect 3608 12786 3660 12792
rect 3620 12442 3648 12786
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3620 10062 3648 12378
rect 3712 12238 3740 12815
rect 3804 12782 3832 14470
rect 4344 14486 4396 14492
rect 4250 14447 4306 14456
rect 4264 14414 4292 14447
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4342 13968 4398 13977
rect 4342 13903 4344 13912
rect 4396 13903 4398 13912
rect 4344 13874 4396 13880
rect 4436 13728 4488 13734
rect 4356 13688 4436 13716
rect 3917 13628 4225 13637
rect 3917 13626 3923 13628
rect 3979 13626 4003 13628
rect 4059 13626 4083 13628
rect 4139 13626 4163 13628
rect 4219 13626 4225 13628
rect 3979 13574 3981 13626
rect 4161 13574 4163 13626
rect 3917 13572 3923 13574
rect 3979 13572 4003 13574
rect 4059 13572 4083 13574
rect 4139 13572 4163 13574
rect 4219 13572 4225 13574
rect 3917 13563 4225 13572
rect 4066 13424 4122 13433
rect 4122 13382 4292 13410
rect 4066 13359 4122 13368
rect 3976 13320 4028 13326
rect 3896 13297 3976 13308
rect 3882 13288 3976 13297
rect 3938 13280 3976 13288
rect 3976 13262 4028 13268
rect 3882 13223 3938 13232
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 3804 12434 3832 12582
rect 3917 12540 4225 12549
rect 3917 12538 3923 12540
rect 3979 12538 4003 12540
rect 4059 12538 4083 12540
rect 4139 12538 4163 12540
rect 4219 12538 4225 12540
rect 3979 12486 3981 12538
rect 4161 12486 4163 12538
rect 3917 12484 3923 12486
rect 3979 12484 4003 12486
rect 4059 12484 4083 12486
rect 4139 12484 4163 12486
rect 4219 12484 4225 12486
rect 3917 12475 4225 12484
rect 4264 12442 4292 13382
rect 4252 12436 4304 12442
rect 3804 12406 3924 12434
rect 3790 12336 3846 12345
rect 3790 12271 3846 12280
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3804 12102 3832 12271
rect 3792 12096 3844 12102
rect 3698 12064 3754 12073
rect 3792 12038 3844 12044
rect 3698 11999 3754 12008
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3606 9752 3662 9761
rect 3606 9687 3662 9696
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3620 9500 3648 9687
rect 3528 9472 3648 9500
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3528 8786 3556 9472
rect 3068 7806 3188 7834
rect 3252 8452 3372 8480
rect 3436 8758 3556 8786
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7342 3004 7686
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2962 6624 3018 6633
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2412 2100 2464 2106
rect 2412 2042 2464 2048
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 1400 1964 1452 1970
rect 1320 1924 1400 1952
rect 1320 160 1348 1924
rect 1400 1906 1452 1912
rect 1676 1964 1728 1970
rect 1676 1906 1728 1912
rect 1400 1352 1452 1358
rect 1400 1294 1452 1300
rect 1676 1352 1728 1358
rect 2044 1352 2096 1358
rect 1676 1294 1728 1300
rect 1858 1320 1914 1329
rect 1412 746 1440 1294
rect 1584 1216 1636 1222
rect 1584 1158 1636 1164
rect 1596 950 1624 1158
rect 1584 944 1636 950
rect 1584 886 1636 892
rect 1400 740 1452 746
rect 1400 682 1452 688
rect 754 54 980 82
rect 754 0 810 54
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 82 1638 160
rect 1688 82 1716 1294
rect 2044 1294 2096 1300
rect 2502 1320 2558 1329
rect 1858 1255 1914 1264
rect 1872 1222 1900 1255
rect 1860 1216 1912 1222
rect 1860 1158 1912 1164
rect 1582 54 1716 82
rect 1858 82 1914 160
rect 2056 82 2084 1294
rect 2320 1284 2372 1290
rect 2502 1255 2504 1264
rect 2320 1226 2372 1232
rect 2556 1255 2558 1264
rect 2504 1226 2556 1232
rect 1858 54 2084 82
rect 2134 82 2190 160
rect 2332 82 2360 1226
rect 2412 740 2464 746
rect 2412 682 2464 688
rect 2424 160 2452 682
rect 2700 160 2728 2926
rect 2792 1562 2820 6598
rect 2884 6582 2962 6610
rect 2962 6559 3018 6568
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 2976 6390 3004 6423
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2962 6216 3018 6225
rect 2962 6151 3018 6160
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5273 2912 5510
rect 2976 5370 3004 6151
rect 3068 5778 3096 7806
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 6254 3188 7686
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2870 5264 2926 5273
rect 2870 5199 2926 5208
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2976 2650 3004 4558
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3068 2446 3096 5306
rect 3146 4176 3202 4185
rect 3146 4111 3202 4120
rect 3160 4078 3188 4111
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3146 3088 3202 3097
rect 3252 3074 3280 8452
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3344 7993 3372 8298
rect 3330 7984 3386 7993
rect 3330 7919 3386 7928
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3344 7410 3372 7822
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3344 5370 3372 6734
rect 3436 6662 3464 8758
rect 3712 8616 3740 11999
rect 3896 11914 3924 12406
rect 4252 12378 4304 12384
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3974 12064 4030 12073
rect 3974 11999 4030 12008
rect 3804 11886 3924 11914
rect 3804 11218 3832 11886
rect 3988 11830 4016 11999
rect 4172 11898 4200 12174
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3917 11452 4225 11461
rect 3917 11450 3923 11452
rect 3979 11450 4003 11452
rect 4059 11450 4083 11452
rect 4139 11450 4163 11452
rect 4219 11450 4225 11452
rect 3979 11398 3981 11450
rect 4161 11398 4163 11450
rect 3917 11396 3923 11398
rect 3979 11396 4003 11398
rect 4059 11396 4083 11398
rect 4139 11396 4163 11398
rect 4219 11396 4225 11398
rect 3917 11387 4225 11396
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3896 11257 3924 11290
rect 3882 11248 3938 11257
rect 3792 11212 3844 11218
rect 3882 11183 3938 11192
rect 3976 11212 4028 11218
rect 3792 11154 3844 11160
rect 3976 11154 4028 11160
rect 3988 11098 4016 11154
rect 3528 8588 3740 8616
rect 3804 11070 4016 11098
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3344 4146 3372 4762
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3330 4040 3386 4049
rect 3436 4026 3464 5743
rect 3528 5234 3556 8588
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 7002 3648 7346
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3606 6896 3662 6905
rect 3606 6831 3662 6840
rect 3620 6798 3648 6831
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3712 6662 3740 8434
rect 3804 7342 3832 11070
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10713 4016 10950
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 4068 10600 4120 10606
rect 4066 10568 4068 10577
rect 4120 10568 4122 10577
rect 4066 10503 4122 10512
rect 3917 10364 4225 10373
rect 3917 10362 3923 10364
rect 3979 10362 4003 10364
rect 4059 10362 4083 10364
rect 4139 10362 4163 10364
rect 4219 10362 4225 10364
rect 3979 10310 3981 10362
rect 4161 10310 4163 10362
rect 3917 10308 3923 10310
rect 3979 10308 4003 10310
rect 4059 10308 4083 10310
rect 4139 10308 4163 10310
rect 4219 10308 4225 10310
rect 3917 10299 4225 10308
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3974 10160 4030 10169
rect 3974 10095 3976 10104
rect 4028 10095 4030 10104
rect 3976 10066 4028 10072
rect 4080 10033 4108 10202
rect 4158 10160 4214 10169
rect 4158 10095 4214 10104
rect 4066 10024 4122 10033
rect 4066 9959 4122 9968
rect 4172 9722 4200 10095
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 3917 9276 4225 9285
rect 3917 9274 3923 9276
rect 3979 9274 4003 9276
rect 4059 9274 4083 9276
rect 4139 9274 4163 9276
rect 4219 9274 4225 9276
rect 3979 9222 3981 9274
rect 4161 9222 4163 9274
rect 3917 9220 3923 9222
rect 3979 9220 4003 9222
rect 4059 9220 4083 9222
rect 4139 9220 4163 9222
rect 4219 9220 4225 9222
rect 3917 9211 4225 9220
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 4264 7886 4292 12242
rect 4356 11150 4384 13688
rect 4436 13670 4488 13676
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4448 12782 4476 13126
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 4448 11558 4476 12310
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4540 11218 4568 16594
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4632 16046 4660 16458
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4712 16040 4764 16046
rect 4816 16028 4844 16748
rect 5000 16454 5028 16918
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4896 16040 4948 16046
rect 4816 16000 4896 16028
rect 4712 15982 4764 15988
rect 4896 15982 4948 15988
rect 4632 12866 4660 15982
rect 4724 15706 4752 15982
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 5092 15586 5120 17711
rect 5172 17264 5224 17270
rect 5172 17206 5224 17212
rect 5184 15688 5212 17206
rect 5276 16522 5304 23990
rect 5368 23662 5396 24262
rect 5460 23662 5488 25230
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5448 22704 5500 22710
rect 5448 22646 5500 22652
rect 5460 22030 5488 22646
rect 5448 22024 5500 22030
rect 5368 21984 5448 22012
rect 5368 19786 5396 21984
rect 5448 21966 5500 21972
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5446 18592 5502 18601
rect 5446 18527 5502 18536
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5368 16182 5396 16526
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 5184 15660 5304 15688
rect 5092 15558 5212 15586
rect 5078 15192 5134 15201
rect 5078 15127 5134 15136
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4724 13938 4752 14758
rect 4816 14414 4844 14758
rect 5000 14414 5028 14962
rect 4804 14408 4856 14414
rect 4802 14376 4804 14385
rect 4988 14408 5040 14414
rect 4856 14376 4858 14385
rect 4988 14350 5040 14356
rect 4802 14311 4858 14320
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 14074 4844 14214
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4632 12838 4752 12866
rect 4724 12782 4752 12838
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4620 12776 4672 12782
rect 4724 12776 4789 12782
rect 4724 12736 4737 12776
rect 4620 12718 4672 12724
rect 4737 12718 4789 12724
rect 4632 12594 4660 12718
rect 4802 12608 4858 12617
rect 4632 12566 4802 12594
rect 4802 12543 4858 12552
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4342 10976 4398 10985
rect 4342 10911 4398 10920
rect 4356 10810 4384 10911
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4356 10674 4384 10746
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4448 10282 4476 11018
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4356 10254 4476 10282
rect 4356 9489 4384 10254
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4448 9722 4476 10066
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4342 9480 4398 9489
rect 4342 9415 4398 9424
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3792 7336 3844 7342
rect 4356 7313 4384 7822
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7342 4476 7686
rect 4436 7336 4488 7342
rect 3792 7278 3844 7284
rect 4342 7304 4398 7313
rect 4436 7278 4488 7284
rect 4342 7239 4398 7248
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 4356 6934 4384 7239
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6440 3924 6598
rect 3712 6412 3924 6440
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5302 3648 6190
rect 3608 5296 3660 5302
rect 3608 5238 3660 5244
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 4146 3556 4626
rect 3620 4146 3648 4966
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3436 3998 3648 4026
rect 3330 3975 3386 3984
rect 3344 3194 3372 3975
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3252 3046 3556 3074
rect 3146 3023 3148 3032
rect 3200 3023 3202 3032
rect 3148 2994 3200 3000
rect 3160 2774 3188 2994
rect 3160 2746 3372 2774
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 2780 1556 2832 1562
rect 2780 1498 2832 1504
rect 3056 1284 3108 1290
rect 3056 1226 3108 1232
rect 2134 54 2360 82
rect 1582 0 1638 54
rect 1858 0 1914 54
rect 2134 0 2190 54
rect 2410 0 2466 160
rect 2686 0 2742 160
rect 2962 82 3018 160
rect 3068 82 3096 1226
rect 3148 1216 3200 1222
rect 3148 1158 3200 1164
rect 3160 882 3188 1158
rect 3148 876 3200 882
rect 3148 818 3200 824
rect 3252 160 3280 2382
rect 3344 2038 3372 2746
rect 3332 2032 3384 2038
rect 3332 1974 3384 1980
rect 3424 1964 3476 1970
rect 3424 1906 3476 1912
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 3344 1494 3372 1702
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 2962 54 3096 82
rect 2962 0 3018 54
rect 3238 0 3294 160
rect 3436 82 3464 1906
rect 3528 1902 3556 3046
rect 3620 2774 3648 3998
rect 3712 3602 3740 6412
rect 3976 6248 4028 6254
rect 4080 6236 4108 6734
rect 4028 6208 4108 6236
rect 3976 6190 4028 6196
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3804 4826 3832 6122
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3896 5710 3924 5850
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3988 5370 4016 5714
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4250 5128 4306 5137
rect 4250 5063 4306 5072
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3976 4616 4028 4622
rect 3974 4584 3976 4593
rect 4028 4584 4030 4593
rect 3974 4519 4030 4528
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 4080 4282 4108 4422
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4264 4026 4292 5063
rect 4356 4078 4384 5510
rect 4448 5234 4476 7278
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4540 4842 4568 10746
rect 4632 7342 4660 12271
rect 4724 9586 4752 12378
rect 4804 12232 4856 12238
rect 4802 12200 4804 12209
rect 4856 12200 4858 12209
rect 4802 12135 4858 12144
rect 4816 10130 4844 12135
rect 4908 11898 4936 12786
rect 5000 12345 5028 14350
rect 5092 13938 5120 15127
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5092 13841 5120 13874
rect 5078 13832 5134 13841
rect 5078 13767 5134 13776
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4986 12336 5042 12345
rect 4986 12271 5042 12280
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4896 11688 4948 11694
rect 4894 11656 4896 11665
rect 4948 11656 4950 11665
rect 4894 11591 4950 11600
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4908 9926 4936 11591
rect 5000 10606 5028 12174
rect 4988 10600 5040 10606
rect 4988 10542 5040 10548
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 10130 5028 10406
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4896 9920 4948 9926
rect 5092 9897 5120 13398
rect 5184 11257 5212 15558
rect 5276 15502 5304 15660
rect 5460 15570 5488 18527
rect 5552 18086 5580 26318
rect 5644 24154 5672 31282
rect 5828 30802 5856 31826
rect 5816 30796 5868 30802
rect 5816 30738 5868 30744
rect 5814 30424 5870 30433
rect 5814 30359 5870 30368
rect 5724 29572 5776 29578
rect 5724 29514 5776 29520
rect 5736 28422 5764 29514
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 5828 26858 5856 30359
rect 5920 30326 5948 34478
rect 6012 31634 6040 36110
rect 6104 35766 6132 36110
rect 6092 35760 6144 35766
rect 6092 35702 6144 35708
rect 6104 32434 6132 35702
rect 6288 35630 6316 36110
rect 6276 35624 6328 35630
rect 6276 35566 6328 35572
rect 6288 35290 6316 35566
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 6276 35284 6328 35290
rect 6276 35226 6328 35232
rect 6196 34542 6224 35226
rect 6380 35136 6408 37742
rect 6288 35108 6408 35136
rect 6184 34536 6236 34542
rect 6184 34478 6236 34484
rect 6196 34241 6224 34478
rect 6182 34232 6238 34241
rect 6182 34167 6238 34176
rect 6196 33930 6224 34167
rect 6184 33924 6236 33930
rect 6184 33866 6236 33872
rect 6196 32978 6224 33866
rect 6184 32972 6236 32978
rect 6184 32914 6236 32920
rect 6184 32768 6236 32774
rect 6184 32710 6236 32716
rect 6196 32570 6224 32710
rect 6184 32564 6236 32570
rect 6184 32506 6236 32512
rect 6092 32428 6144 32434
rect 6092 32370 6144 32376
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6012 31606 6132 31634
rect 6000 31408 6052 31414
rect 6000 31350 6052 31356
rect 5908 30320 5960 30326
rect 5908 30262 5960 30268
rect 5908 30184 5960 30190
rect 5908 30126 5960 30132
rect 5816 26852 5868 26858
rect 5816 26794 5868 26800
rect 5816 25696 5868 25702
rect 5920 25684 5948 30126
rect 6012 30122 6040 31350
rect 6104 31142 6132 31606
rect 6196 31346 6224 32370
rect 6184 31340 6236 31346
rect 6184 31282 6236 31288
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 6104 30938 6132 31078
rect 6092 30932 6144 30938
rect 6092 30874 6144 30880
rect 6104 30569 6132 30874
rect 6090 30560 6146 30569
rect 6090 30495 6146 30504
rect 6000 30116 6052 30122
rect 6000 30058 6052 30064
rect 6196 29850 6224 31282
rect 6184 29844 6236 29850
rect 6184 29786 6236 29792
rect 6092 29708 6144 29714
rect 6012 29668 6092 29696
rect 6012 25974 6040 29668
rect 6092 29650 6144 29656
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 6104 29345 6132 29446
rect 6090 29336 6146 29345
rect 6090 29271 6092 29280
rect 6144 29271 6146 29280
rect 6092 29242 6144 29248
rect 6092 28008 6144 28014
rect 6092 27950 6144 27956
rect 6104 27849 6132 27950
rect 6090 27840 6146 27849
rect 6090 27775 6146 27784
rect 6090 27568 6146 27577
rect 6090 27503 6146 27512
rect 6104 27470 6132 27503
rect 6092 27464 6144 27470
rect 6092 27406 6144 27412
rect 6090 26616 6146 26625
rect 6090 26551 6146 26560
rect 6104 26450 6132 26551
rect 6092 26444 6144 26450
rect 6092 26386 6144 26392
rect 6000 25968 6052 25974
rect 6000 25910 6052 25916
rect 6012 25809 6040 25910
rect 5998 25800 6054 25809
rect 5998 25735 6054 25744
rect 6104 25702 6132 26386
rect 6196 26246 6224 29786
rect 6184 26240 6236 26246
rect 6184 26182 6236 26188
rect 6092 25696 6144 25702
rect 5920 25656 6040 25684
rect 5816 25638 5868 25644
rect 5724 24608 5776 24614
rect 5828 24596 5856 25638
rect 5776 24568 5856 24596
rect 5724 24550 5776 24556
rect 5828 24342 5856 24568
rect 5908 24608 5960 24614
rect 5908 24550 5960 24556
rect 5920 24410 5948 24550
rect 5908 24404 5960 24410
rect 5908 24346 5960 24352
rect 5816 24336 5868 24342
rect 5816 24278 5868 24284
rect 5908 24268 5960 24274
rect 5908 24210 5960 24216
rect 5644 24126 5764 24154
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5644 21865 5672 21898
rect 5630 21856 5686 21865
rect 5630 21791 5686 21800
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5644 19854 5672 20878
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5630 18456 5686 18465
rect 5630 18391 5632 18400
rect 5684 18391 5686 18400
rect 5632 18362 5684 18368
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5264 15088 5316 15094
rect 5264 15030 5316 15036
rect 5170 11248 5226 11257
rect 5170 11183 5226 11192
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10130 5212 10542
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 4896 9862 4948 9868
rect 5078 9888 5134 9897
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4632 5273 4660 7278
rect 4724 6322 4752 9522
rect 4908 9518 4936 9862
rect 5078 9823 5134 9832
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 8294 4936 9454
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5184 7750 5212 10066
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 5000 6458 5028 7210
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4724 5370 4752 5714
rect 4988 5568 5040 5574
rect 4802 5536 4858 5545
rect 4988 5510 5040 5516
rect 4802 5471 4858 5480
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4618 5264 4674 5273
rect 4618 5199 4674 5208
rect 4632 5166 4660 5199
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4448 4814 4568 4842
rect 4172 3998 4292 4026
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4172 3942 4200 3998
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3620 2746 3740 2774
rect 3712 2650 3740 2746
rect 3804 2650 3832 3402
rect 4448 3194 4476 4814
rect 4526 4720 4582 4729
rect 4526 4655 4582 4664
rect 4540 3194 4568 4655
rect 4724 4622 4752 5306
rect 4816 4622 4844 5471
rect 5000 5166 5028 5510
rect 5092 5166 5120 7278
rect 5170 6216 5226 6225
rect 5170 6151 5226 6160
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4908 4622 4936 5102
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4894 4448 4950 4457
rect 4894 4383 4950 4392
rect 4908 3738 4936 4383
rect 5092 4214 5120 5102
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2774 4476 2994
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 4356 2746 4476 2774
rect 5092 2774 5120 3470
rect 5184 3398 5212 6151
rect 5276 5710 5304 15030
rect 5460 14822 5488 15506
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5368 14550 5396 14758
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5552 13326 5580 17478
rect 5644 16969 5672 18226
rect 5630 16960 5686 16969
rect 5630 16895 5686 16904
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5368 12442 5396 13126
rect 5446 12608 5502 12617
rect 5446 12543 5502 12552
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5356 8084 5408 8090
rect 5460 8072 5488 12543
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 11898 5580 12242
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5644 10810 5672 16895
rect 5736 13462 5764 24126
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5828 21350 5856 21966
rect 5920 21894 5948 24210
rect 6012 23118 6040 25656
rect 6092 25638 6144 25644
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 6104 23769 6132 25094
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6196 24410 6224 24550
rect 6184 24404 6236 24410
rect 6184 24346 6236 24352
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 6288 24154 6316 35108
rect 6472 34066 6500 39374
rect 7288 39296 7340 39302
rect 7288 39238 7340 39244
rect 6884 39196 7192 39205
rect 6884 39194 6890 39196
rect 6946 39194 6970 39196
rect 7026 39194 7050 39196
rect 7106 39194 7130 39196
rect 7186 39194 7192 39196
rect 6946 39142 6948 39194
rect 7128 39142 7130 39194
rect 6884 39140 6890 39142
rect 6946 39140 6970 39142
rect 7026 39140 7050 39142
rect 7106 39140 7130 39142
rect 7186 39140 7192 39142
rect 6884 39131 7192 39140
rect 7300 39098 7328 39238
rect 7392 39098 7420 40870
rect 7288 39092 7340 39098
rect 7288 39034 7340 39040
rect 7380 39092 7432 39098
rect 7380 39034 7432 39040
rect 6736 38956 6788 38962
rect 6736 38898 6788 38904
rect 7380 38956 7432 38962
rect 7380 38898 7432 38904
rect 6552 38344 6604 38350
rect 6552 38286 6604 38292
rect 6564 38010 6592 38286
rect 6552 38004 6604 38010
rect 6552 37946 6604 37952
rect 6748 37874 6776 38898
rect 6884 38108 7192 38117
rect 6884 38106 6890 38108
rect 6946 38106 6970 38108
rect 7026 38106 7050 38108
rect 7106 38106 7130 38108
rect 7186 38106 7192 38108
rect 6946 38054 6948 38106
rect 7128 38054 7130 38106
rect 6884 38052 6890 38054
rect 6946 38052 6970 38054
rect 7026 38052 7050 38054
rect 7106 38052 7130 38054
rect 7186 38052 7192 38054
rect 6884 38043 7192 38052
rect 6552 37868 6604 37874
rect 6552 37810 6604 37816
rect 6736 37868 6788 37874
rect 6736 37810 6788 37816
rect 6564 37754 6592 37810
rect 7104 37800 7156 37806
rect 6564 37748 7104 37754
rect 6564 37742 7156 37748
rect 6564 37726 7144 37742
rect 6564 37097 6592 37726
rect 6642 37632 6698 37641
rect 6642 37567 6698 37576
rect 6550 37088 6606 37097
rect 6550 37023 6606 37032
rect 6656 34728 6684 37567
rect 7288 37324 7340 37330
rect 7288 37266 7340 37272
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6748 36582 6776 37062
rect 6884 37020 7192 37029
rect 6884 37018 6890 37020
rect 6946 37018 6970 37020
rect 7026 37018 7050 37020
rect 7106 37018 7130 37020
rect 7186 37018 7192 37020
rect 6946 36966 6948 37018
rect 7128 36966 7130 37018
rect 6884 36964 6890 36966
rect 6946 36964 6970 36966
rect 7026 36964 7050 36966
rect 7106 36964 7130 36966
rect 7186 36964 7192 36966
rect 6884 36955 7192 36964
rect 7300 36786 7328 37266
rect 7392 36904 7420 38898
rect 7484 37466 7512 40870
rect 7576 39545 7604 41210
rect 7944 41138 7972 41386
rect 8024 41268 8076 41274
rect 8024 41210 8076 41216
rect 7932 41132 7984 41138
rect 7932 41074 7984 41080
rect 7748 40928 7800 40934
rect 7748 40870 7800 40876
rect 7840 40928 7892 40934
rect 7840 40870 7892 40876
rect 7656 40452 7708 40458
rect 7656 40394 7708 40400
rect 7668 40186 7696 40394
rect 7656 40180 7708 40186
rect 7656 40122 7708 40128
rect 7760 40089 7788 40870
rect 7852 40526 7880 40870
rect 8036 40730 8064 41210
rect 8024 40724 8076 40730
rect 8024 40666 8076 40672
rect 7840 40520 7892 40526
rect 7840 40462 7892 40468
rect 7746 40080 7802 40089
rect 7746 40015 7802 40024
rect 7852 39828 7880 40462
rect 7932 40384 7984 40390
rect 7932 40326 7984 40332
rect 8024 40384 8076 40390
rect 8024 40326 8076 40332
rect 7944 39982 7972 40326
rect 8036 40118 8064 40326
rect 8024 40112 8076 40118
rect 8024 40054 8076 40060
rect 7932 39976 7984 39982
rect 7932 39918 7984 39924
rect 7852 39800 7972 39828
rect 7748 39636 7800 39642
rect 7748 39578 7800 39584
rect 7562 39536 7618 39545
rect 7562 39471 7618 39480
rect 7564 39432 7616 39438
rect 7564 39374 7616 39380
rect 7576 39302 7604 39374
rect 7564 39296 7616 39302
rect 7564 39238 7616 39244
rect 7576 37806 7604 39238
rect 7656 39092 7708 39098
rect 7656 39034 7708 39040
rect 7564 37800 7616 37806
rect 7564 37742 7616 37748
rect 7472 37460 7524 37466
rect 7472 37402 7524 37408
rect 7564 37392 7616 37398
rect 7564 37334 7616 37340
rect 7392 36876 7512 36904
rect 6920 36780 6972 36786
rect 6920 36722 6972 36728
rect 7288 36780 7340 36786
rect 7288 36722 7340 36728
rect 7380 36780 7432 36786
rect 7380 36722 7432 36728
rect 6736 36576 6788 36582
rect 6736 36518 6788 36524
rect 6564 34700 6684 34728
rect 6460 34060 6512 34066
rect 6460 34002 6512 34008
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6380 33114 6408 33934
rect 6460 33856 6512 33862
rect 6460 33798 6512 33804
rect 6368 33108 6420 33114
rect 6368 33050 6420 33056
rect 6366 33008 6422 33017
rect 6366 32943 6422 32952
rect 6380 31226 6408 32943
rect 6472 32434 6500 33798
rect 6460 32428 6512 32434
rect 6460 32370 6512 32376
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6472 31521 6500 31758
rect 6458 31512 6514 31521
rect 6458 31447 6514 31456
rect 6380 31198 6500 31226
rect 6368 30796 6420 30802
rect 6368 30738 6420 30744
rect 6380 30122 6408 30738
rect 6472 30297 6500 31198
rect 6564 30734 6592 34700
rect 6644 34604 6696 34610
rect 6644 34546 6696 34552
rect 6656 31754 6684 34546
rect 6748 32502 6776 36518
rect 6932 36378 6960 36722
rect 7288 36644 7340 36650
rect 7288 36586 7340 36592
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 7300 36310 7328 36586
rect 7288 36304 7340 36310
rect 7288 36246 7340 36252
rect 7392 36242 7420 36722
rect 7380 36236 7432 36242
rect 7380 36178 7432 36184
rect 7288 36168 7340 36174
rect 7288 36110 7340 36116
rect 6884 35932 7192 35941
rect 6884 35930 6890 35932
rect 6946 35930 6970 35932
rect 7026 35930 7050 35932
rect 7106 35930 7130 35932
rect 7186 35930 7192 35932
rect 6946 35878 6948 35930
rect 7128 35878 7130 35930
rect 6884 35876 6890 35878
rect 6946 35876 6970 35878
rect 7026 35876 7050 35878
rect 7106 35876 7130 35878
rect 7186 35876 7192 35878
rect 6884 35867 7192 35876
rect 7300 35834 7328 36110
rect 7288 35828 7340 35834
rect 7288 35770 7340 35776
rect 7484 35494 7512 36876
rect 7576 36038 7604 37334
rect 7668 36961 7696 39034
rect 7760 39030 7788 39578
rect 7748 39024 7800 39030
rect 7748 38966 7800 38972
rect 7760 38826 7788 38966
rect 7944 38894 7972 39800
rect 7932 38888 7984 38894
rect 7932 38830 7984 38836
rect 7748 38820 7800 38826
rect 7748 38762 7800 38768
rect 7654 36952 7710 36961
rect 7654 36887 7710 36896
rect 7656 36780 7708 36786
rect 7656 36722 7708 36728
rect 7668 36689 7696 36722
rect 7654 36680 7710 36689
rect 7944 36666 7972 38830
rect 8128 37126 8156 41670
rect 8576 41608 8628 41614
rect 8576 41550 8628 41556
rect 8588 41414 8616 41550
rect 8588 41386 8800 41414
rect 8576 41064 8628 41070
rect 8576 41006 8628 41012
rect 8392 40384 8444 40390
rect 8392 40326 8444 40332
rect 8208 40112 8260 40118
rect 8208 40054 8260 40060
rect 8220 38593 8248 40054
rect 8404 39642 8432 40326
rect 8392 39636 8444 39642
rect 8392 39578 8444 39584
rect 8588 39438 8616 41006
rect 8576 39432 8628 39438
rect 8576 39374 8628 39380
rect 8484 39024 8536 39030
rect 8484 38966 8536 38972
rect 8206 38584 8262 38593
rect 8206 38519 8262 38528
rect 8496 38350 8524 38966
rect 8588 38758 8616 39374
rect 8576 38752 8628 38758
rect 8576 38694 8628 38700
rect 8484 38344 8536 38350
rect 8484 38286 8536 38292
rect 8576 37936 8628 37942
rect 8576 37878 8628 37884
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8116 37120 8168 37126
rect 8116 37062 8168 37068
rect 8496 36922 8524 37198
rect 8588 36922 8616 37878
rect 8668 37256 8720 37262
rect 8668 37198 8720 37204
rect 8484 36916 8536 36922
rect 8484 36858 8536 36864
rect 8576 36916 8628 36922
rect 8576 36858 8628 36864
rect 7654 36615 7710 36624
rect 7852 36638 7972 36666
rect 8484 36712 8536 36718
rect 8484 36654 8536 36660
rect 7564 36032 7616 36038
rect 7564 35974 7616 35980
rect 7472 35488 7524 35494
rect 7524 35448 7696 35476
rect 7472 35430 7524 35436
rect 7288 35148 7340 35154
rect 7288 35090 7340 35096
rect 6884 34844 7192 34853
rect 6884 34842 6890 34844
rect 6946 34842 6970 34844
rect 7026 34842 7050 34844
rect 7106 34842 7130 34844
rect 7186 34842 7192 34844
rect 6946 34790 6948 34842
rect 7128 34790 7130 34842
rect 6884 34788 6890 34790
rect 6946 34788 6970 34790
rect 7026 34788 7050 34790
rect 7106 34788 7130 34790
rect 7186 34788 7192 34790
rect 6884 34779 7192 34788
rect 6826 34096 6882 34105
rect 6826 34031 6828 34040
rect 6880 34031 6882 34040
rect 6828 34002 6880 34008
rect 6884 33756 7192 33765
rect 6884 33754 6890 33756
rect 6946 33754 6970 33756
rect 7026 33754 7050 33756
rect 7106 33754 7130 33756
rect 7186 33754 7192 33756
rect 6946 33702 6948 33754
rect 7128 33702 7130 33754
rect 6884 33700 6890 33702
rect 6946 33700 6970 33702
rect 7026 33700 7050 33702
rect 7106 33700 7130 33702
rect 7186 33700 7192 33702
rect 6884 33691 7192 33700
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 6920 33448 6972 33454
rect 6920 33390 6972 33396
rect 7116 33402 7144 33594
rect 7300 33522 7328 35090
rect 7564 35012 7616 35018
rect 7564 34954 7616 34960
rect 7380 34400 7432 34406
rect 7380 34342 7432 34348
rect 7392 34134 7420 34342
rect 7380 34128 7432 34134
rect 7380 34070 7432 34076
rect 7288 33516 7340 33522
rect 7288 33458 7340 33464
rect 7196 33448 7248 33454
rect 7116 33396 7196 33402
rect 7248 33396 7328 33402
rect 6932 32881 6960 33390
rect 7116 33374 7328 33396
rect 7392 33386 7420 34070
rect 7470 33552 7526 33561
rect 7470 33487 7526 33496
rect 6918 32872 6974 32881
rect 6918 32807 6974 32816
rect 7300 32745 7328 33374
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7484 32910 7512 33487
rect 7472 32904 7524 32910
rect 7472 32846 7524 32852
rect 7576 32756 7604 34954
rect 7668 32881 7696 35448
rect 7852 33561 7880 36638
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 8300 36168 8352 36174
rect 8300 36110 8352 36116
rect 8116 36032 8168 36038
rect 8116 35974 8168 35980
rect 7932 35216 7984 35222
rect 7932 35158 7984 35164
rect 7838 33552 7894 33561
rect 7838 33487 7894 33496
rect 7654 32872 7710 32881
rect 7654 32807 7710 32816
rect 7286 32736 7342 32745
rect 6884 32668 7192 32677
rect 7286 32671 7342 32680
rect 7392 32728 7604 32756
rect 6884 32666 6890 32668
rect 6946 32666 6970 32668
rect 7026 32666 7050 32668
rect 7106 32666 7130 32668
rect 7186 32666 7192 32668
rect 6946 32614 6948 32666
rect 7128 32614 7130 32666
rect 6884 32612 6890 32614
rect 6946 32612 6970 32614
rect 7026 32612 7050 32614
rect 7106 32612 7130 32614
rect 7186 32612 7192 32614
rect 6884 32603 7192 32612
rect 6736 32496 6788 32502
rect 6736 32438 6788 32444
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6840 31754 6868 31894
rect 6644 31748 6696 31754
rect 6644 31690 6696 31696
rect 6748 31726 6868 31754
rect 6642 31648 6698 31657
rect 6642 31583 6698 31592
rect 6656 31346 6684 31583
rect 6644 31340 6696 31346
rect 6644 31282 6696 31288
rect 6748 31278 6776 31726
rect 6884 31580 7192 31589
rect 6884 31578 6890 31580
rect 6946 31578 6970 31580
rect 7026 31578 7050 31580
rect 7106 31578 7130 31580
rect 7186 31578 7192 31580
rect 6946 31526 6948 31578
rect 7128 31526 7130 31578
rect 6884 31524 6890 31526
rect 6946 31524 6970 31526
rect 7026 31524 7050 31526
rect 7106 31524 7130 31526
rect 7186 31524 7192 31526
rect 6884 31515 7192 31524
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 6736 31272 6788 31278
rect 6736 31214 6788 31220
rect 7116 30938 7144 31282
rect 6644 30932 6696 30938
rect 6644 30874 6696 30880
rect 7104 30932 7156 30938
rect 7104 30874 7156 30880
rect 6552 30728 6604 30734
rect 6552 30670 6604 30676
rect 6458 30288 6514 30297
rect 6458 30223 6514 30232
rect 6368 30116 6420 30122
rect 6368 30058 6420 30064
rect 6460 30116 6512 30122
rect 6460 30058 6512 30064
rect 6380 28014 6408 30058
rect 6472 29481 6500 30058
rect 6564 30025 6592 30670
rect 6550 30016 6606 30025
rect 6550 29951 6606 29960
rect 6458 29472 6514 29481
rect 6458 29407 6514 29416
rect 6472 29102 6500 29407
rect 6460 29096 6512 29102
rect 6460 29038 6512 29044
rect 6368 28008 6420 28014
rect 6368 27950 6420 27956
rect 6656 27402 6684 30874
rect 7288 30660 7340 30666
rect 7288 30602 7340 30608
rect 6884 30492 7192 30501
rect 6884 30490 6890 30492
rect 6946 30490 6970 30492
rect 7026 30490 7050 30492
rect 7106 30490 7130 30492
rect 7186 30490 7192 30492
rect 6946 30438 6948 30490
rect 7128 30438 7130 30490
rect 6884 30436 6890 30438
rect 6946 30436 6970 30438
rect 7026 30436 7050 30438
rect 7106 30436 7130 30438
rect 7186 30436 7192 30438
rect 6884 30427 7192 30436
rect 6828 30320 6880 30326
rect 6734 30288 6790 30297
rect 6828 30262 6880 30268
rect 6734 30223 6790 30232
rect 6748 30190 6776 30223
rect 6736 30184 6788 30190
rect 6736 30126 6788 30132
rect 6840 29628 6868 30262
rect 7300 30138 7328 30602
rect 7116 30110 7328 30138
rect 7116 29782 7144 30110
rect 7104 29776 7156 29782
rect 7104 29718 7156 29724
rect 6920 29640 6972 29646
rect 6748 29600 6920 29628
rect 6748 28098 6776 29600
rect 6920 29582 6972 29588
rect 7288 29640 7340 29646
rect 7288 29582 7340 29588
rect 7300 29492 7328 29582
rect 6822 29481 7328 29492
rect 6822 29472 7342 29481
rect 6822 29464 7286 29472
rect 6822 29288 6850 29464
rect 6884 29404 7192 29413
rect 7286 29407 7342 29416
rect 6884 29402 6890 29404
rect 6946 29402 6970 29404
rect 7026 29402 7050 29404
rect 7106 29402 7130 29404
rect 7186 29402 7192 29404
rect 6946 29350 6948 29402
rect 7128 29350 7130 29402
rect 6884 29348 6890 29350
rect 6946 29348 6970 29350
rect 7026 29348 7050 29350
rect 7106 29348 7130 29350
rect 7186 29348 7192 29350
rect 6884 29339 7192 29348
rect 6822 29260 7052 29288
rect 7024 28994 7052 29260
rect 7288 29096 7340 29102
rect 7288 29038 7340 29044
rect 7024 28966 7236 28994
rect 7208 28801 7236 28966
rect 7194 28792 7250 28801
rect 7194 28727 7250 28736
rect 7300 28626 7328 29038
rect 7288 28620 7340 28626
rect 7288 28562 7340 28568
rect 6884 28316 7192 28325
rect 6884 28314 6890 28316
rect 6946 28314 6970 28316
rect 7026 28314 7050 28316
rect 7106 28314 7130 28316
rect 7186 28314 7192 28316
rect 6946 28262 6948 28314
rect 7128 28262 7130 28314
rect 6884 28260 6890 28262
rect 6946 28260 6970 28262
rect 7026 28260 7050 28262
rect 7106 28260 7130 28262
rect 7186 28260 7192 28262
rect 6884 28251 7192 28260
rect 6748 28070 6868 28098
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 6748 27470 6776 27814
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6552 27396 6604 27402
rect 6552 27338 6604 27344
rect 6644 27396 6696 27402
rect 6644 27338 6696 27344
rect 6460 27328 6512 27334
rect 6366 27296 6422 27305
rect 6422 27276 6460 27282
rect 6422 27270 6512 27276
rect 6422 27254 6500 27270
rect 6366 27231 6422 27240
rect 6564 27130 6592 27338
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6564 25362 6592 26386
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 6380 24750 6408 25094
rect 6460 24812 6512 24818
rect 6460 24754 6512 24760
rect 6368 24744 6420 24750
rect 6368 24686 6420 24692
rect 6380 24274 6408 24686
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6196 24070 6224 24142
rect 6288 24126 6408 24154
rect 6184 24064 6236 24070
rect 6236 24024 6316 24052
rect 6184 24006 6236 24012
rect 6090 23760 6146 23769
rect 6090 23695 6146 23704
rect 6000 23112 6052 23118
rect 6000 23054 6052 23060
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6092 22772 6144 22778
rect 6092 22714 6144 22720
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5908 21548 5960 21554
rect 5908 21490 5960 21496
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5920 20942 5948 21490
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5828 19922 5856 20198
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5828 19514 5856 19722
rect 5816 19508 5868 19514
rect 5816 19450 5868 19456
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5828 14414 5856 19110
rect 5920 18902 5948 20198
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 6012 18737 6040 22102
rect 6104 21554 6132 22714
rect 6196 22574 6224 23054
rect 6184 22568 6236 22574
rect 6184 22510 6236 22516
rect 6196 22098 6224 22510
rect 6184 22092 6236 22098
rect 6184 22034 6236 22040
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 6196 21690 6224 21830
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 5998 18728 6054 18737
rect 5998 18663 6054 18672
rect 6104 18601 6132 20742
rect 6090 18592 6146 18601
rect 6090 18527 6146 18536
rect 5906 17368 5962 17377
rect 5906 17303 5962 17312
rect 5920 16658 5948 17303
rect 6196 17134 6224 21626
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6196 16998 6224 17070
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 6288 16538 6316 24024
rect 6380 20806 6408 24126
rect 6472 23594 6500 24754
rect 6460 23588 6512 23594
rect 6460 23530 6512 23536
rect 6564 23118 6592 25298
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6656 22964 6684 27338
rect 6840 27316 6868 28070
rect 6748 27288 6868 27316
rect 7288 27328 7340 27334
rect 6748 23526 6776 27288
rect 7288 27270 7340 27276
rect 6884 27228 7192 27237
rect 6884 27226 6890 27228
rect 6946 27226 6970 27228
rect 7026 27226 7050 27228
rect 7106 27226 7130 27228
rect 7186 27226 7192 27228
rect 6946 27174 6948 27226
rect 7128 27174 7130 27226
rect 6884 27172 6890 27174
rect 6946 27172 6970 27174
rect 7026 27172 7050 27174
rect 7106 27172 7130 27174
rect 7186 27172 7192 27174
rect 6884 27163 7192 27172
rect 6826 26480 6882 26489
rect 6826 26415 6882 26424
rect 6840 26382 6868 26415
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6884 26140 7192 26149
rect 6884 26138 6890 26140
rect 6946 26138 6970 26140
rect 7026 26138 7050 26140
rect 7106 26138 7130 26140
rect 7186 26138 7192 26140
rect 6946 26086 6948 26138
rect 7128 26086 7130 26138
rect 6884 26084 6890 26086
rect 6946 26084 6970 26086
rect 7026 26084 7050 26086
rect 7106 26084 7130 26086
rect 7186 26084 7192 26086
rect 6884 26075 7192 26084
rect 7300 25974 7328 27270
rect 7104 25968 7156 25974
rect 7104 25910 7156 25916
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7116 25702 7144 25910
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 6918 25392 6974 25401
rect 6918 25327 6974 25336
rect 7286 25392 7342 25401
rect 7286 25327 7288 25336
rect 6932 25294 6960 25327
rect 7340 25327 7342 25336
rect 7288 25298 7340 25304
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6884 25052 7192 25061
rect 6884 25050 6890 25052
rect 6946 25050 6970 25052
rect 7026 25050 7050 25052
rect 7106 25050 7130 25052
rect 7186 25050 7192 25052
rect 6946 24998 6948 25050
rect 7128 24998 7130 25050
rect 6884 24996 6890 24998
rect 6946 24996 6970 24998
rect 7026 24996 7050 24998
rect 7106 24996 7130 24998
rect 7186 24996 7192 24998
rect 6884 24987 7192 24996
rect 6884 23964 7192 23973
rect 6884 23962 6890 23964
rect 6946 23962 6970 23964
rect 7026 23962 7050 23964
rect 7106 23962 7130 23964
rect 7186 23962 7192 23964
rect 6946 23910 6948 23962
rect 7128 23910 7130 23962
rect 6884 23908 6890 23910
rect 6946 23908 6970 23910
rect 7026 23908 7050 23910
rect 7106 23908 7130 23910
rect 7186 23908 7192 23910
rect 6884 23899 7192 23908
rect 6736 23520 6788 23526
rect 6736 23462 6788 23468
rect 6736 23044 6788 23050
rect 6736 22986 6788 22992
rect 6472 22936 6684 22964
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6366 20632 6422 20641
rect 6366 20567 6422 20576
rect 6380 20233 6408 20567
rect 6366 20224 6422 20233
rect 6366 20159 6422 20168
rect 6472 19802 6500 22936
rect 6550 22808 6606 22817
rect 6606 22766 6684 22794
rect 6550 22743 6606 22752
rect 6656 22522 6684 22766
rect 6748 22642 6776 22986
rect 6884 22876 7192 22885
rect 6884 22874 6890 22876
rect 6946 22874 6970 22876
rect 7026 22874 7050 22876
rect 7106 22874 7130 22876
rect 7186 22874 7192 22876
rect 6946 22822 6948 22874
rect 7128 22822 7130 22874
rect 6884 22820 6890 22822
rect 6946 22820 6970 22822
rect 7026 22820 7050 22822
rect 7106 22820 7130 22822
rect 7186 22820 7192 22822
rect 6884 22811 7192 22820
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6656 22494 6868 22522
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6552 22160 6604 22166
rect 6604 22108 6684 22114
rect 6552 22102 6684 22108
rect 6564 22086 6684 22102
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 20856 6592 21966
rect 6656 21622 6684 22086
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6748 21486 6776 22374
rect 6840 22030 6868 22494
rect 7392 22094 7420 32728
rect 7852 32450 7880 33487
rect 7944 33454 7972 35158
rect 8024 33992 8076 33998
rect 8024 33934 8076 33940
rect 8036 33504 8064 33934
rect 8128 33640 8156 35974
rect 8128 33612 8248 33640
rect 8116 33516 8168 33522
rect 8036 33476 8116 33504
rect 8116 33458 8168 33464
rect 7932 33448 7984 33454
rect 7932 33390 7984 33396
rect 7576 32422 7880 32450
rect 7576 31754 7604 32422
rect 7576 31726 7788 31754
rect 7656 31680 7708 31686
rect 7656 31622 7708 31628
rect 7668 31482 7696 31622
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7484 29850 7512 30534
rect 7564 30252 7616 30258
rect 7564 30194 7616 30200
rect 7472 29844 7524 29850
rect 7472 29786 7524 29792
rect 7470 29744 7526 29753
rect 7470 29679 7526 29688
rect 7484 28994 7512 29679
rect 7576 29628 7604 30194
rect 7760 29730 7788 31726
rect 7944 31346 7972 33390
rect 8128 33114 8156 33458
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 8220 32994 8248 33612
rect 8036 32966 8248 32994
rect 7932 31340 7984 31346
rect 7932 31282 7984 31288
rect 7840 31136 7892 31142
rect 7840 31078 7892 31084
rect 7852 30569 7880 31078
rect 7838 30560 7894 30569
rect 7838 30495 7894 30504
rect 8036 30258 8064 32966
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8128 30666 8156 32846
rect 8208 32428 8260 32434
rect 8208 32370 8260 32376
rect 8220 31142 8248 32370
rect 8312 32314 8340 36110
rect 8404 35630 8432 36518
rect 8392 35624 8444 35630
rect 8392 35566 8444 35572
rect 8496 35476 8524 36654
rect 8588 36122 8616 36858
rect 8680 36718 8708 37198
rect 8668 36712 8720 36718
rect 8668 36654 8720 36660
rect 8588 36094 8708 36122
rect 8576 36032 8628 36038
rect 8576 35974 8628 35980
rect 8588 35766 8616 35974
rect 8576 35760 8628 35766
rect 8576 35702 8628 35708
rect 8404 35448 8524 35476
rect 8404 32434 8432 35448
rect 8484 34604 8536 34610
rect 8484 34546 8536 34552
rect 8496 34134 8524 34546
rect 8484 34128 8536 34134
rect 8484 34070 8536 34076
rect 8392 32428 8444 32434
rect 8392 32370 8444 32376
rect 8312 32286 8432 32314
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 8116 30660 8168 30666
rect 8116 30602 8168 30608
rect 8114 30424 8170 30433
rect 8114 30359 8170 30368
rect 8024 30252 8076 30258
rect 8024 30194 8076 30200
rect 7840 30048 7892 30054
rect 7840 29990 7892 29996
rect 7852 29850 7880 29990
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 8128 29730 8156 30359
rect 7760 29702 7880 29730
rect 7576 29600 7696 29628
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7576 28994 7604 29106
rect 7484 28966 7604 28994
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 7300 22066 7420 22094
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6884 21788 7192 21797
rect 6884 21786 6890 21788
rect 6946 21786 6970 21788
rect 7026 21786 7050 21788
rect 7106 21786 7130 21788
rect 7186 21786 7192 21788
rect 6946 21734 6948 21786
rect 7128 21734 7130 21786
rect 6884 21732 6890 21734
rect 6946 21732 6970 21734
rect 7026 21732 7050 21734
rect 7106 21732 7130 21734
rect 7186 21732 7192 21734
rect 6884 21723 7192 21732
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 7116 21146 7144 21626
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 6564 20828 6684 20856
rect 6550 20768 6606 20777
rect 6550 20703 6606 20712
rect 6380 19774 6500 19802
rect 6380 19514 6408 19774
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6472 19009 6500 19654
rect 6458 19000 6514 19009
rect 6458 18935 6514 18944
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6380 17610 6408 18702
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6380 16658 6408 17546
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6012 16510 6316 16538
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 5722 12336 5778 12345
rect 5722 12271 5778 12280
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5408 8044 5488 8072
rect 5356 8026 5408 8032
rect 5460 7410 5488 8044
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5460 6474 5488 7346
rect 5552 7002 5580 7346
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5460 6446 5580 6474
rect 5644 6458 5672 9862
rect 5736 7721 5764 12271
rect 5828 10810 5856 14350
rect 5920 13938 5948 14758
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5920 13462 5948 13874
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5722 7712 5778 7721
rect 5722 7647 5778 7656
rect 5828 6798 5856 10610
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5722 6488 5778 6497
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5914 5396 6054
rect 5460 5914 5488 6326
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5552 5794 5580 6446
rect 5632 6452 5684 6458
rect 5722 6423 5724 6432
rect 5632 6394 5684 6400
rect 5776 6423 5778 6432
rect 5724 6394 5776 6400
rect 5368 5766 5580 5794
rect 5920 5778 5948 13262
rect 6012 10266 6040 16510
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6288 16182 6316 16390
rect 6276 16176 6328 16182
rect 6196 16124 6276 16130
rect 6196 16118 6328 16124
rect 6196 16102 6316 16118
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6104 14074 6132 14350
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6104 12850 6132 13330
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6104 12238 6132 12582
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6104 10130 6132 12038
rect 6196 10674 6224 16102
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6288 15502 6316 15982
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6288 13190 6316 15438
rect 6472 15314 6500 18022
rect 6380 15286 6500 15314
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6380 12986 6408 15286
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6472 14890 6500 15098
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 14385 6500 14418
rect 6458 14376 6514 14385
rect 6458 14311 6514 14320
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6274 12336 6330 12345
rect 6274 12271 6330 12280
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 5998 10024 6054 10033
rect 5998 9959 6054 9968
rect 5908 5772 5960 5778
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5368 5234 5396 5766
rect 5908 5714 5960 5720
rect 5816 5704 5868 5710
rect 5446 5672 5502 5681
rect 5816 5646 5868 5652
rect 5446 5607 5502 5616
rect 5356 5228 5408 5234
rect 5276 5188 5356 5216
rect 5276 4826 5304 5188
rect 5356 5170 5408 5176
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5368 2922 5396 4694
rect 5460 3534 5488 5607
rect 5828 5370 5856 5646
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5552 4826 5580 5102
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 6012 2774 6040 9959
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6104 7313 6132 8366
rect 6196 7410 6224 10134
rect 6288 7954 6316 12271
rect 6366 12200 6422 12209
rect 6366 12135 6422 12144
rect 6380 11898 6408 12135
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6472 10962 6500 13874
rect 6380 10934 6500 10962
rect 6380 10266 6408 10934
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6472 10130 6500 10746
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6380 9722 6408 10066
rect 6458 10024 6514 10033
rect 6458 9959 6514 9968
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6090 7304 6146 7313
rect 6090 7239 6092 7248
rect 6144 7239 6146 7248
rect 6092 7210 6144 7216
rect 6104 5914 6132 7210
rect 6288 6322 6316 7890
rect 6380 7886 6408 9454
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6276 6316 6328 6322
rect 6380 6304 6408 7822
rect 6472 7460 6500 9959
rect 6564 7562 6592 20703
rect 6656 20534 6684 20828
rect 6884 20700 7192 20709
rect 6884 20698 6890 20700
rect 6946 20698 6970 20700
rect 7026 20698 7050 20700
rect 7106 20698 7130 20700
rect 7186 20698 7192 20700
rect 6946 20646 6948 20698
rect 7128 20646 7130 20698
rect 6884 20644 6890 20646
rect 6946 20644 6970 20646
rect 7026 20644 7050 20646
rect 7106 20644 7130 20646
rect 7186 20644 7192 20646
rect 6884 20635 7192 20644
rect 6644 20528 6696 20534
rect 6696 20488 6776 20516
rect 6644 20470 6696 20476
rect 6748 19786 6776 20488
rect 7300 20262 7328 22066
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21622 7420 21830
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 7288 19848 7340 19854
rect 6826 19816 6882 19825
rect 6736 19780 6788 19786
rect 7288 19790 7340 19796
rect 7380 19848 7432 19854
rect 7484 19825 7512 28358
rect 7576 28082 7604 28966
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7562 27704 7618 27713
rect 7668 27690 7696 29600
rect 7748 28620 7800 28626
rect 7748 28562 7800 28568
rect 7618 27662 7696 27690
rect 7562 27639 7618 27648
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 26897 7696 27270
rect 7760 26994 7788 28562
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7654 26888 7710 26897
rect 7654 26823 7710 26832
rect 7852 26382 7880 29702
rect 8036 29702 8156 29730
rect 7932 29640 7984 29646
rect 7932 29582 7984 29588
rect 7944 29238 7972 29582
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 7944 27538 7972 29174
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 7840 26376 7892 26382
rect 7892 26336 7972 26364
rect 7840 26318 7892 26324
rect 7564 26240 7616 26246
rect 7564 26182 7616 26188
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7576 25838 7604 26182
rect 7852 26042 7880 26182
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7668 25650 7696 25842
rect 7668 25622 7788 25650
rect 7760 25498 7788 25622
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7576 25106 7604 25230
rect 7576 25078 7788 25106
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7576 23118 7604 24006
rect 7668 23866 7696 24074
rect 7656 23860 7708 23866
rect 7656 23802 7708 23808
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7668 22094 7696 23462
rect 7576 22066 7696 22094
rect 7576 21434 7604 22066
rect 7656 21616 7708 21622
rect 7654 21584 7656 21593
rect 7708 21584 7710 21593
rect 7654 21519 7710 21528
rect 7576 21406 7696 21434
rect 7562 20768 7618 20777
rect 7562 20703 7618 20712
rect 7380 19790 7432 19796
rect 7470 19816 7526 19825
rect 6826 19751 6828 19760
rect 6736 19722 6788 19728
rect 6880 19751 6882 19760
rect 6828 19722 6880 19728
rect 6748 18834 6776 19722
rect 6884 19612 7192 19621
rect 6884 19610 6890 19612
rect 6946 19610 6970 19612
rect 7026 19610 7050 19612
rect 7106 19610 7130 19612
rect 7186 19610 7192 19612
rect 6946 19558 6948 19610
rect 7128 19558 7130 19610
rect 6884 19556 6890 19558
rect 6946 19556 6970 19558
rect 7026 19556 7050 19558
rect 7106 19556 7130 19558
rect 7186 19556 7192 19558
rect 6884 19547 7192 19556
rect 7194 19408 7250 19417
rect 7194 19343 7196 19352
rect 7248 19343 7250 19352
rect 7196 19314 7248 19320
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 7104 18692 7156 18698
rect 7300 18680 7328 19790
rect 7392 19378 7420 19790
rect 7470 19751 7526 19760
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7484 18970 7512 19314
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7156 18652 7328 18680
rect 7104 18634 7156 18640
rect 6884 18524 7192 18533
rect 6884 18522 6890 18524
rect 6946 18522 6970 18524
rect 7026 18522 7050 18524
rect 7106 18522 7130 18524
rect 7186 18522 7192 18524
rect 6946 18470 6948 18522
rect 7128 18470 7130 18522
rect 6884 18468 6890 18470
rect 6946 18468 6970 18470
rect 7026 18468 7050 18470
rect 7106 18468 7130 18470
rect 7186 18468 7192 18470
rect 6884 18459 7192 18468
rect 6918 18184 6974 18193
rect 6918 18119 6974 18128
rect 6932 17678 6960 18119
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 7286 17640 7342 17649
rect 7286 17575 7342 17584
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6748 17338 6776 17478
rect 6884 17436 7192 17445
rect 6884 17434 6890 17436
rect 6946 17434 6970 17436
rect 7026 17434 7050 17436
rect 7106 17434 7130 17436
rect 7186 17434 7192 17436
rect 6946 17382 6948 17434
rect 7128 17382 7130 17434
rect 6884 17380 6890 17382
rect 6946 17380 6970 17382
rect 7026 17380 7050 17382
rect 7106 17380 7130 17382
rect 7186 17380 7192 17382
rect 6884 17371 7192 17380
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6644 17264 6696 17270
rect 6642 17232 6644 17241
rect 6696 17232 6698 17241
rect 6932 17202 6960 17274
rect 6642 17167 6698 17176
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 6840 17105 6868 17138
rect 6826 17096 6882 17105
rect 6826 17031 6882 17040
rect 7208 16969 7236 17138
rect 7194 16960 7250 16969
rect 7194 16895 7250 16904
rect 7300 16810 7328 17575
rect 7576 16810 7604 20703
rect 7668 19922 7696 21406
rect 7760 20754 7788 25078
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7852 23186 7880 23462
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7944 22953 7972 26336
rect 8036 24818 8064 29702
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 8128 29306 8156 29582
rect 8206 29336 8262 29345
rect 8116 29300 8168 29306
rect 8206 29271 8262 29280
rect 8116 29242 8168 29248
rect 8116 29028 8168 29034
rect 8220 29016 8248 29271
rect 8168 28988 8248 29016
rect 8116 28970 8168 28976
rect 8116 28552 8168 28558
rect 8116 28494 8168 28500
rect 8128 28082 8156 28494
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 8312 27554 8340 31826
rect 8128 27526 8340 27554
rect 8128 26994 8156 27526
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8128 25158 8156 26930
rect 8220 25906 8248 27270
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 8220 24954 8248 25842
rect 8300 25832 8352 25838
rect 8300 25774 8352 25780
rect 8312 24954 8340 25774
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8300 24948 8352 24954
rect 8300 24890 8352 24896
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 8312 24682 8340 24890
rect 8300 24676 8352 24682
rect 8300 24618 8352 24624
rect 8298 24304 8354 24313
rect 8404 24290 8432 32286
rect 8496 31890 8524 34070
rect 8680 33946 8708 36094
rect 8588 33918 8708 33946
rect 8588 32609 8616 33918
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8680 33658 8708 33798
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8574 32600 8630 32609
rect 8574 32535 8630 32544
rect 8576 32496 8628 32502
rect 8576 32438 8628 32444
rect 8484 31884 8536 31890
rect 8484 31826 8536 31832
rect 8496 31793 8524 31826
rect 8482 31784 8538 31793
rect 8482 31719 8538 31728
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8496 25945 8524 31622
rect 8588 30802 8616 32438
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8576 30796 8628 30802
rect 8576 30738 8628 30744
rect 8482 25936 8538 25945
rect 8482 25871 8538 25880
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8354 24262 8432 24290
rect 8298 24239 8354 24248
rect 8116 24064 8168 24070
rect 8116 24006 8168 24012
rect 8128 23798 8156 24006
rect 8116 23792 8168 23798
rect 8116 23734 8168 23740
rect 8208 23724 8260 23730
rect 8208 23666 8260 23672
rect 8220 23526 8248 23666
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 23118 8432 23462
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 7930 22944 7986 22953
rect 7930 22879 7986 22888
rect 8116 22772 8168 22778
rect 8116 22714 8168 22720
rect 7840 22704 7892 22710
rect 7840 22646 7892 22652
rect 7852 20942 7880 22646
rect 7840 20936 7892 20942
rect 7892 20896 8064 20924
rect 7840 20878 7892 20884
rect 8036 20777 8064 20896
rect 8022 20768 8078 20777
rect 7760 20726 7972 20754
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 19310 7696 19654
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7760 17320 7788 19450
rect 7852 19446 7880 20538
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7852 18698 7880 19382
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7944 18465 7972 20726
rect 8022 20703 8078 20712
rect 8024 19916 8076 19922
rect 8024 19858 8076 19864
rect 8036 19378 8064 19858
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 7930 18456 7986 18465
rect 7930 18391 7986 18400
rect 7838 18048 7894 18057
rect 7944 18034 7972 18391
rect 8024 18352 8076 18358
rect 8024 18294 8076 18300
rect 7894 18006 7972 18034
rect 7838 17983 7894 17992
rect 7760 17292 7972 17320
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7656 17128 7708 17134
rect 7708 17088 7788 17116
rect 7656 17070 7708 17076
rect 7024 16782 7512 16810
rect 7576 16782 7696 16810
rect 6828 16720 6880 16726
rect 6826 16688 6828 16697
rect 6880 16688 6882 16697
rect 6736 16652 6788 16658
rect 7024 16658 7052 16782
rect 6826 16623 6882 16632
rect 7012 16652 7064 16658
rect 6736 16594 6788 16600
rect 7012 16594 7064 16600
rect 7196 16652 7248 16658
rect 7248 16612 7420 16640
rect 7196 16594 7248 16600
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 15065 6684 16526
rect 6642 15056 6698 15065
rect 6642 14991 6698 15000
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6656 12832 6684 14894
rect 6748 14414 6776 16594
rect 6884 16348 7192 16357
rect 6884 16346 6890 16348
rect 6946 16346 6970 16348
rect 7026 16346 7050 16348
rect 7106 16346 7130 16348
rect 7186 16346 7192 16348
rect 6946 16294 6948 16346
rect 7128 16294 7130 16346
rect 6884 16292 6890 16294
rect 6946 16292 6970 16294
rect 7026 16292 7050 16294
rect 7106 16292 7130 16294
rect 7186 16292 7192 16294
rect 6884 16283 7192 16292
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7300 15706 7328 15982
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 6884 15260 7192 15269
rect 6884 15258 6890 15260
rect 6946 15258 6970 15260
rect 7026 15258 7050 15260
rect 7106 15258 7130 15260
rect 7186 15258 7192 15260
rect 6946 15206 6948 15258
rect 7128 15206 7130 15258
rect 6884 15204 6890 15206
rect 6946 15204 6970 15206
rect 7026 15204 7050 15206
rect 7106 15204 7130 15206
rect 7186 15204 7192 15206
rect 6884 15195 7192 15204
rect 7300 14822 7328 15302
rect 7392 15162 7420 16612
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7484 15026 7512 16782
rect 7564 16720 7616 16726
rect 7564 16662 7616 16668
rect 7576 15706 7604 16662
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 6840 14482 6868 14758
rect 7576 14618 7604 14894
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7668 14498 7696 16782
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 7576 14470 7696 14498
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6918 14376 6974 14385
rect 6918 14311 6974 14320
rect 7380 14340 7432 14346
rect 6932 14278 6960 14311
rect 7380 14282 7432 14288
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6748 14074 6776 14214
rect 6884 14172 7192 14181
rect 6884 14170 6890 14172
rect 6946 14170 6970 14172
rect 7026 14170 7050 14172
rect 7106 14170 7130 14172
rect 7186 14170 7192 14172
rect 6946 14118 6948 14170
rect 7128 14118 7130 14170
rect 6884 14116 6890 14118
rect 6946 14116 6970 14118
rect 7026 14116 7050 14118
rect 7106 14116 7130 14118
rect 7186 14116 7192 14118
rect 6884 14107 7192 14116
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 7012 14000 7064 14006
rect 6840 13960 7012 13988
rect 6840 13870 6868 13960
rect 7392 13977 7420 14282
rect 7012 13942 7064 13948
rect 7378 13968 7434 13977
rect 7378 13903 7434 13912
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 6884 13084 7192 13093
rect 6884 13082 6890 13084
rect 6946 13082 6970 13084
rect 7026 13082 7050 13084
rect 7106 13082 7130 13084
rect 7186 13082 7192 13084
rect 6946 13030 6948 13082
rect 7128 13030 7130 13082
rect 6884 13028 6890 13030
rect 6946 13028 6970 13030
rect 7026 13028 7050 13030
rect 7106 13028 7130 13030
rect 7186 13028 7192 13030
rect 6884 13019 7192 13028
rect 7300 12986 7328 13126
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6736 12844 6788 12850
rect 6656 12804 6736 12832
rect 6736 12786 6788 12792
rect 6826 12472 6882 12481
rect 7102 12472 7158 12481
rect 6932 12442 7102 12458
rect 6826 12407 6882 12416
rect 6920 12436 7102 12442
rect 6840 12306 6868 12407
rect 6972 12430 7102 12436
rect 7102 12407 7158 12416
rect 6920 12378 6972 12384
rect 6932 12347 6960 12378
rect 6828 12300 6880 12306
rect 6656 12260 6828 12288
rect 6656 10112 6684 12260
rect 6828 12242 6880 12248
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11354 6776 12038
rect 6884 11996 7192 12005
rect 6884 11994 6890 11996
rect 6946 11994 6970 11996
rect 7026 11994 7050 11996
rect 7106 11994 7130 11996
rect 7186 11994 7192 11996
rect 6946 11942 6948 11994
rect 7128 11942 7130 11994
rect 6884 11940 6890 11942
rect 6946 11940 6970 11942
rect 7026 11940 7050 11942
rect 7106 11940 7130 11942
rect 7186 11940 7192 11942
rect 6884 11931 7192 11940
rect 7300 11762 7328 12922
rect 7392 12617 7420 12922
rect 7378 12608 7434 12617
rect 7378 12543 7434 12552
rect 7392 12442 7420 12543
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7576 12356 7604 14470
rect 7656 14408 7708 14414
rect 7656 14350 7708 14356
rect 7668 14074 7696 14350
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7576 12328 7696 12356
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7378 12200 7434 12209
rect 7378 12135 7434 12144
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 7024 11082 7052 11494
rect 7392 11150 7420 12135
rect 7484 11354 7512 12242
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6884 10908 7192 10917
rect 6884 10906 6890 10908
rect 6946 10906 6970 10908
rect 7026 10906 7050 10908
rect 7106 10906 7130 10908
rect 7186 10906 7192 10908
rect 6946 10854 6948 10906
rect 7128 10854 7130 10906
rect 6884 10852 6890 10854
rect 6946 10852 6970 10854
rect 7026 10852 7050 10854
rect 7106 10852 7130 10854
rect 7186 10852 7192 10854
rect 6884 10843 7192 10852
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 6736 10124 6788 10130
rect 6656 10084 6736 10112
rect 6736 10066 6788 10072
rect 6840 9926 6868 10406
rect 7392 10266 7420 10406
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6884 9820 7192 9829
rect 6884 9818 6890 9820
rect 6946 9818 6970 9820
rect 7026 9818 7050 9820
rect 7106 9818 7130 9820
rect 7186 9818 7192 9820
rect 6946 9766 6948 9818
rect 7128 9766 7130 9818
rect 6884 9764 6890 9766
rect 6946 9764 6970 9766
rect 7026 9764 7050 9766
rect 7106 9764 7130 9766
rect 7186 9764 7192 9766
rect 6884 9755 7192 9764
rect 6884 8732 7192 8741
rect 6884 8730 6890 8732
rect 6946 8730 6970 8732
rect 7026 8730 7050 8732
rect 7106 8730 7130 8732
rect 7186 8730 7192 8732
rect 6946 8678 6948 8730
rect 7128 8678 7130 8730
rect 6884 8676 6890 8678
rect 6946 8676 6970 8678
rect 7026 8676 7050 8678
rect 7106 8676 7130 8678
rect 7186 8676 7192 8678
rect 6884 8667 7192 8676
rect 7300 8616 7328 10202
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7208 8588 7328 8616
rect 7208 8294 7236 8588
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 8090 7236 8230
rect 7300 8090 7328 8434
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7194 7984 7250 7993
rect 7392 7970 7420 9658
rect 7484 9178 7512 10746
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7576 10266 7604 10678
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7484 8566 7512 8910
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7194 7919 7196 7928
rect 7248 7919 7250 7928
rect 7300 7942 7420 7970
rect 7196 7890 7248 7896
rect 6884 7644 7192 7653
rect 6884 7642 6890 7644
rect 6946 7642 6970 7644
rect 7026 7642 7050 7644
rect 7106 7642 7130 7644
rect 7186 7642 7192 7644
rect 6946 7590 6948 7642
rect 7128 7590 7130 7642
rect 6884 7588 6890 7590
rect 6946 7588 6970 7590
rect 7026 7588 7050 7590
rect 7106 7588 7130 7590
rect 7186 7588 7192 7590
rect 6884 7579 7192 7588
rect 6564 7534 6776 7562
rect 6472 7432 6592 7460
rect 6460 6316 6512 6322
rect 6380 6276 6460 6304
rect 6276 6258 6328 6264
rect 6460 6258 6512 6264
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6104 4146 6132 5850
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6380 5234 6408 5510
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6366 3768 6422 3777
rect 6366 3703 6368 3712
rect 6420 3703 6422 3712
rect 6368 3674 6420 3680
rect 6472 3618 6500 5238
rect 6380 3590 6500 3618
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6104 2990 6132 3334
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6196 2922 6224 3431
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 6288 2825 6316 3130
rect 5092 2746 5304 2774
rect 3700 2644 3752 2650
rect 3700 2586 3752 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3974 2272 4030 2281
rect 3974 2207 4030 2216
rect 3988 2106 4016 2207
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 4160 1964 4212 1970
rect 4212 1924 4292 1952
rect 4160 1906 4212 1912
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3804 1426 3832 1906
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 4264 1442 4292 1924
rect 3792 1420 3844 1426
rect 3792 1362 3844 1368
rect 4080 1414 4292 1442
rect 3884 1284 3936 1290
rect 3884 1226 3936 1232
rect 3792 1216 3844 1222
rect 3792 1158 3844 1164
rect 3804 160 3832 1158
rect 3896 1018 3924 1226
rect 3884 1012 3936 1018
rect 3884 954 3936 960
rect 4080 160 4108 1414
rect 4356 950 4384 2746
rect 4894 2680 4950 2689
rect 4894 2615 4950 2624
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4436 1284 4488 1290
rect 4436 1226 4488 1232
rect 4344 944 4396 950
rect 4344 886 4396 892
rect 4448 678 4476 1226
rect 4436 672 4488 678
rect 4436 614 4488 620
rect 3514 82 3570 160
rect 3436 54 3570 82
rect 3514 0 3570 54
rect 3790 0 3846 160
rect 4066 0 4122 160
rect 4342 82 4398 160
rect 4540 82 4568 2382
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 4632 160 4660 1974
rect 4908 1562 4936 2615
rect 5276 2514 5304 2746
rect 5644 2746 6040 2774
rect 6274 2816 6330 2825
rect 6274 2751 6330 2760
rect 5644 2650 5672 2746
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6182 2544 6238 2553
rect 5264 2508 5316 2514
rect 6182 2479 6238 2488
rect 5264 2450 5316 2456
rect 4988 2440 5040 2446
rect 5448 2440 5500 2446
rect 5040 2400 5212 2428
rect 4988 2382 5040 2388
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4986 2136 5042 2145
rect 4986 2071 4988 2080
rect 5040 2071 5042 2080
rect 4988 2042 5040 2048
rect 5092 1970 5120 2246
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 5080 1760 5132 1766
rect 5078 1728 5080 1737
rect 5132 1728 5134 1737
rect 5078 1663 5134 1672
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 4712 1420 4764 1426
rect 4712 1362 4764 1368
rect 4724 1034 4752 1362
rect 4988 1216 5040 1222
rect 5080 1216 5132 1222
rect 4988 1158 5040 1164
rect 5078 1184 5080 1193
rect 5132 1184 5134 1193
rect 4724 1006 4936 1034
rect 4908 160 4936 1006
rect 5000 542 5028 1158
rect 5078 1119 5134 1128
rect 5184 950 5212 2400
rect 5500 2400 5764 2428
rect 5448 2382 5500 2388
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5276 2106 5304 2246
rect 5368 2106 5396 2246
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5264 1352 5316 1358
rect 5264 1294 5316 1300
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 4988 536 5040 542
rect 4988 478 5040 484
rect 4342 54 4568 82
rect 4342 0 4398 54
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5170 82 5226 160
rect 5276 82 5304 1294
rect 5460 160 5488 2246
rect 5540 1352 5592 1358
rect 5538 1320 5540 1329
rect 5736 1340 5764 2400
rect 5814 2272 5870 2281
rect 5814 2207 5870 2216
rect 5828 2038 5856 2207
rect 5816 2032 5868 2038
rect 5816 1974 5868 1980
rect 6196 1970 6224 2479
rect 6380 1986 6408 3590
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3126 6500 3334
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 6564 2961 6592 7432
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6656 5642 6684 6938
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6550 2952 6606 2961
rect 6460 2916 6512 2922
rect 6550 2887 6606 2896
rect 6460 2858 6512 2864
rect 6472 2446 6500 2858
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 2106 6500 2246
rect 6656 2106 6684 3130
rect 6748 2106 6776 7534
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 7300 3670 7328 7942
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7392 6322 7420 7822
rect 7484 7546 7512 7822
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7576 7426 7604 8434
rect 7484 7398 7604 7426
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7392 5030 7420 6054
rect 7484 5234 7512 7398
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 5914 7604 6258
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7576 5234 7604 5578
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7392 3670 7420 4150
rect 7576 4146 7604 5034
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7380 3664 7432 3670
rect 7380 3606 7432 3612
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6840 2961 6868 2994
rect 6826 2952 6882 2961
rect 6826 2887 6882 2896
rect 6932 2650 6960 2994
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 6184 1964 6236 1970
rect 6380 1958 6500 1986
rect 6184 1906 6236 1912
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5592 1320 5594 1329
rect 5736 1312 5856 1340
rect 5538 1255 5594 1264
rect 5828 1018 5856 1312
rect 5920 1034 5948 1838
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6276 1216 6328 1222
rect 6276 1158 6328 1164
rect 5816 1012 5868 1018
rect 5920 1006 6040 1034
rect 5816 954 5868 960
rect 5540 672 5592 678
rect 5592 632 5764 660
rect 5540 614 5592 620
rect 5736 160 5764 632
rect 6012 160 6040 1006
rect 6288 160 6316 1158
rect 6380 678 6408 1294
rect 6472 1222 6500 1958
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6564 1562 6592 1906
rect 7300 1850 7328 2994
rect 7392 2650 7420 3606
rect 7668 2774 7696 12328
rect 7760 11218 7788 17088
rect 7852 16590 7880 17138
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7838 14920 7894 14929
rect 7838 14855 7894 14864
rect 7852 14074 7880 14855
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 12782 7880 13670
rect 7944 12986 7972 17292
rect 8036 14414 8064 18294
rect 8128 17270 8156 22714
rect 8496 22166 8524 25434
rect 8588 24410 8616 30738
rect 8680 25226 8708 31078
rect 8772 29850 8800 41386
rect 8864 39098 8892 41670
rect 9048 41670 9352 41698
rect 8944 40384 8996 40390
rect 8944 40326 8996 40332
rect 8852 39092 8904 39098
rect 8852 39034 8904 39040
rect 8852 38344 8904 38350
rect 8852 38286 8904 38292
rect 8864 36174 8892 38286
rect 8956 37942 8984 40326
rect 8944 37936 8996 37942
rect 8944 37878 8996 37884
rect 8852 36168 8904 36174
rect 8852 36110 8904 36116
rect 8956 35834 8984 37878
rect 8944 35828 8996 35834
rect 8944 35770 8996 35776
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 8864 35601 8892 35634
rect 8850 35592 8906 35601
rect 8850 35527 8906 35536
rect 8956 35193 8984 35770
rect 8942 35184 8998 35193
rect 8942 35119 8998 35128
rect 8944 35080 8996 35086
rect 8944 35022 8996 35028
rect 8850 34232 8906 34241
rect 8850 34167 8906 34176
rect 8864 34066 8892 34167
rect 8852 34060 8904 34066
rect 8852 34002 8904 34008
rect 8850 33960 8906 33969
rect 8850 33895 8906 33904
rect 8760 29844 8812 29850
rect 8760 29786 8812 29792
rect 8758 29336 8814 29345
rect 8758 29271 8814 29280
rect 8772 29238 8800 29271
rect 8760 29232 8812 29238
rect 8760 29174 8812 29180
rect 8758 29064 8814 29073
rect 8758 28999 8814 29008
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8576 24064 8628 24070
rect 8576 24006 8628 24012
rect 8588 23662 8616 24006
rect 8576 23656 8628 23662
rect 8576 23598 8628 23604
rect 8484 22160 8536 22166
rect 8484 22102 8536 22108
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8220 21457 8248 21966
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8206 21448 8262 21457
rect 8404 21434 8432 21830
rect 8496 21690 8524 22102
rect 8576 22024 8628 22030
rect 8576 21966 8628 21972
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8206 21383 8262 21392
rect 8312 21406 8432 21434
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8312 21298 8340 21406
rect 8220 21270 8340 21298
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8220 21010 8248 21270
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8208 20800 8260 20806
rect 8260 20760 8340 20788
rect 8208 20742 8260 20748
rect 8206 19952 8262 19961
rect 8206 19887 8262 19896
rect 8220 19514 8248 19887
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8312 19394 8340 20760
rect 8220 19366 8340 19394
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8128 16250 8156 16594
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8220 15978 8248 19366
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18426 8340 19110
rect 8404 18873 8432 21286
rect 8496 21146 8524 21422
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8390 18864 8446 18873
rect 8390 18799 8446 18808
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8312 16266 8340 18362
rect 8496 18290 8524 20946
rect 8588 20466 8616 21966
rect 8680 21894 8708 24754
rect 8772 24614 8800 28999
rect 8864 28558 8892 33895
rect 8852 28552 8904 28558
rect 8852 28494 8904 28500
rect 8850 28112 8906 28121
rect 8850 28047 8906 28056
rect 8864 25498 8892 28047
rect 8956 26874 8984 35022
rect 9048 34746 9076 41670
rect 9416 41562 9444 43318
rect 9496 43308 9548 43314
rect 9496 43250 9548 43256
rect 9956 43308 10008 43314
rect 10152 43296 10180 44463
rect 10008 43268 10180 43296
rect 10324 43308 10376 43314
rect 9956 43250 10008 43256
rect 10428 43296 10456 44463
rect 10508 43648 10560 43654
rect 10508 43590 10560 43596
rect 10520 43450 10548 43590
rect 10508 43444 10560 43450
rect 10508 43386 10560 43392
rect 10704 43314 10732 44463
rect 10376 43268 10456 43296
rect 10692 43308 10744 43314
rect 10324 43250 10376 43256
rect 10980 43296 11008 44463
rect 11152 43376 11204 43382
rect 11152 43318 11204 43324
rect 11060 43308 11112 43314
rect 10980 43268 11060 43296
rect 10692 43250 10744 43256
rect 11060 43250 11112 43256
rect 9508 42906 9536 43250
rect 9680 43240 9732 43246
rect 9680 43182 9732 43188
rect 9692 42906 9720 43182
rect 10600 43172 10652 43178
rect 10600 43114 10652 43120
rect 9772 43104 9824 43110
rect 9772 43046 9824 43052
rect 10140 43104 10192 43110
rect 10192 43064 10272 43092
rect 10140 43046 10192 43052
rect 9496 42900 9548 42906
rect 9496 42842 9548 42848
rect 9680 42900 9732 42906
rect 9680 42842 9732 42848
rect 9588 42696 9640 42702
rect 9588 42638 9640 42644
rect 9494 42256 9550 42265
rect 9494 42191 9496 42200
rect 9548 42191 9550 42200
rect 9496 42162 9548 42168
rect 9600 41585 9628 42638
rect 9784 42566 9812 43046
rect 9851 43004 10159 43013
rect 9851 43002 9857 43004
rect 9913 43002 9937 43004
rect 9993 43002 10017 43004
rect 10073 43002 10097 43004
rect 10153 43002 10159 43004
rect 9913 42950 9915 43002
rect 10095 42950 10097 43002
rect 9851 42948 9857 42950
rect 9913 42948 9937 42950
rect 9993 42948 10017 42950
rect 10073 42948 10097 42950
rect 10153 42948 10159 42950
rect 9851 42939 10159 42948
rect 9772 42560 9824 42566
rect 9772 42502 9824 42508
rect 9772 42288 9824 42294
rect 9824 42265 9904 42276
rect 9824 42256 9918 42265
rect 9824 42248 9862 42256
rect 9772 42230 9824 42236
rect 9862 42191 9918 42200
rect 9772 42016 9824 42022
rect 9772 41958 9824 41964
rect 9784 41800 9812 41958
rect 9851 41916 10159 41925
rect 9851 41914 9857 41916
rect 9913 41914 9937 41916
rect 9993 41914 10017 41916
rect 10073 41914 10097 41916
rect 10153 41914 10159 41916
rect 9913 41862 9915 41914
rect 10095 41862 10097 41914
rect 9851 41860 9857 41862
rect 9913 41860 9937 41862
rect 9993 41860 10017 41862
rect 10073 41860 10097 41862
rect 10153 41860 10159 41862
rect 9851 41851 10159 41860
rect 9784 41772 9996 41800
rect 9680 41608 9732 41614
rect 9324 41534 9444 41562
rect 9586 41576 9642 41585
rect 9128 40384 9180 40390
rect 9128 40326 9180 40332
rect 9140 40118 9168 40326
rect 9324 40118 9352 41534
rect 9864 41608 9916 41614
rect 9732 41585 9812 41596
rect 9732 41576 9826 41585
rect 9732 41568 9770 41576
rect 9680 41550 9732 41556
rect 9586 41511 9642 41520
rect 9692 41414 9720 41550
rect 9864 41550 9916 41556
rect 9770 41511 9826 41520
rect 9416 41386 9720 41414
rect 9128 40112 9180 40118
rect 9128 40054 9180 40060
rect 9312 40112 9364 40118
rect 9312 40054 9364 40060
rect 9324 38876 9352 40054
rect 9416 39438 9444 41386
rect 9692 41138 9720 41386
rect 9680 41132 9732 41138
rect 9680 41074 9732 41080
rect 9496 41064 9548 41070
rect 9496 41006 9548 41012
rect 9508 40633 9536 41006
rect 9876 41002 9904 41550
rect 9968 41478 9996 41772
rect 9956 41472 10008 41478
rect 9956 41414 10008 41420
rect 9864 40996 9916 41002
rect 9864 40938 9916 40944
rect 9588 40928 9640 40934
rect 9588 40870 9640 40876
rect 9494 40624 9550 40633
rect 9494 40559 9550 40568
rect 9600 39982 9628 40870
rect 9851 40828 10159 40837
rect 9851 40826 9857 40828
rect 9913 40826 9937 40828
rect 9993 40826 10017 40828
rect 10073 40826 10097 40828
rect 10153 40826 10159 40828
rect 9913 40774 9915 40826
rect 10095 40774 10097 40826
rect 9851 40772 9857 40774
rect 9913 40772 9937 40774
rect 9993 40772 10017 40774
rect 10073 40772 10097 40774
rect 10153 40772 10159 40774
rect 9851 40763 10159 40772
rect 9772 40112 9824 40118
rect 9772 40054 9824 40060
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9588 39976 9640 39982
rect 9588 39918 9640 39924
rect 9404 39432 9456 39438
rect 9404 39374 9456 39380
rect 9232 38848 9352 38876
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9140 37806 9168 38694
rect 9232 38554 9260 38848
rect 9416 38740 9444 39374
rect 9324 38712 9444 38740
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 9232 37942 9260 38490
rect 9220 37936 9272 37942
rect 9220 37878 9272 37884
rect 9128 37800 9180 37806
rect 9128 37742 9180 37748
rect 9126 36816 9182 36825
rect 9126 36751 9128 36760
rect 9180 36751 9182 36760
rect 9128 36722 9180 36728
rect 9140 36174 9168 36722
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 9232 35834 9260 37878
rect 9220 35828 9272 35834
rect 9220 35770 9272 35776
rect 9324 35680 9352 38712
rect 9692 38593 9720 39986
rect 9784 39642 9812 40054
rect 9851 39740 10159 39749
rect 9851 39738 9857 39740
rect 9913 39738 9937 39740
rect 9993 39738 10017 39740
rect 10073 39738 10097 39740
rect 10153 39738 10159 39740
rect 9913 39686 9915 39738
rect 10095 39686 10097 39738
rect 9851 39684 9857 39686
rect 9913 39684 9937 39686
rect 9993 39684 10017 39686
rect 10073 39684 10097 39686
rect 10153 39684 10159 39686
rect 9851 39675 10159 39684
rect 9772 39636 9824 39642
rect 9772 39578 9824 39584
rect 9772 39432 9824 39438
rect 9772 39374 9824 39380
rect 9678 38584 9734 38593
rect 9678 38519 9734 38528
rect 9404 38344 9456 38350
rect 9404 38286 9456 38292
rect 9416 36281 9444 38286
rect 9692 37874 9720 38519
rect 9680 37868 9732 37874
rect 9680 37810 9732 37816
rect 9402 36272 9458 36281
rect 9402 36207 9458 36216
rect 9588 35828 9640 35834
rect 9588 35770 9640 35776
rect 9404 35760 9456 35766
rect 9140 35652 9352 35680
rect 9402 35728 9404 35737
rect 9456 35728 9458 35737
rect 9402 35663 9458 35672
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 9034 34232 9090 34241
rect 9034 34167 9090 34176
rect 9048 33658 9076 34167
rect 9036 33652 9088 33658
rect 9036 33594 9088 33600
rect 9140 32434 9168 35652
rect 9600 35612 9628 35770
rect 9692 35766 9720 37810
rect 9784 36650 9812 39374
rect 9851 38652 10159 38661
rect 9851 38650 9857 38652
rect 9913 38650 9937 38652
rect 9993 38650 10017 38652
rect 10073 38650 10097 38652
rect 10153 38650 10159 38652
rect 9913 38598 9915 38650
rect 10095 38598 10097 38650
rect 9851 38596 9857 38598
rect 9913 38596 9937 38598
rect 9993 38596 10017 38598
rect 10073 38596 10097 38598
rect 10153 38596 10159 38598
rect 9851 38587 10159 38596
rect 10140 38208 10192 38214
rect 10140 38150 10192 38156
rect 10152 38010 10180 38150
rect 10140 38004 10192 38010
rect 10140 37946 10192 37952
rect 9851 37564 10159 37573
rect 9851 37562 9857 37564
rect 9913 37562 9937 37564
rect 9993 37562 10017 37564
rect 10073 37562 10097 37564
rect 10153 37562 10159 37564
rect 9913 37510 9915 37562
rect 10095 37510 10097 37562
rect 9851 37508 9857 37510
rect 9913 37508 9937 37510
rect 9993 37508 10017 37510
rect 10073 37508 10097 37510
rect 10153 37508 10159 37510
rect 9851 37499 10159 37508
rect 10048 37324 10100 37330
rect 10048 37266 10100 37272
rect 10060 36718 10088 37266
rect 10048 36712 10100 36718
rect 10048 36654 10100 36660
rect 9772 36644 9824 36650
rect 9772 36586 9824 36592
rect 9851 36476 10159 36485
rect 9851 36474 9857 36476
rect 9913 36474 9937 36476
rect 9993 36474 10017 36476
rect 10073 36474 10097 36476
rect 10153 36474 10159 36476
rect 9913 36422 9915 36474
rect 10095 36422 10097 36474
rect 9851 36420 9857 36422
rect 9913 36420 9937 36422
rect 9993 36420 10017 36422
rect 10073 36420 10097 36422
rect 10153 36420 10159 36422
rect 9851 36411 10159 36420
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 9680 35760 9732 35766
rect 9680 35702 9732 35708
rect 9324 35584 9628 35612
rect 9680 35624 9732 35630
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 9036 32224 9088 32230
rect 9036 32166 9088 32172
rect 9048 31906 9076 32166
rect 9048 31878 9168 31906
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 9048 30938 9076 31282
rect 9140 31278 9168 31878
rect 9232 31686 9260 32846
rect 9220 31680 9272 31686
rect 9220 31622 9272 31628
rect 9324 31414 9352 35584
rect 9680 35566 9732 35572
rect 9404 35488 9456 35494
rect 9404 35430 9456 35436
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9416 34202 9444 35430
rect 9600 35290 9628 35430
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 9692 34678 9720 35566
rect 9784 35086 9812 36110
rect 9851 35388 10159 35397
rect 9851 35386 9857 35388
rect 9913 35386 9937 35388
rect 9993 35386 10017 35388
rect 10073 35386 10097 35388
rect 10153 35386 10159 35388
rect 9913 35334 9915 35386
rect 10095 35334 10097 35386
rect 9851 35332 9857 35334
rect 9913 35332 9937 35334
rect 9993 35332 10017 35334
rect 10073 35332 10097 35334
rect 10153 35332 10159 35334
rect 9851 35323 10159 35332
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9680 34672 9732 34678
rect 9680 34614 9732 34620
rect 9496 34604 9548 34610
rect 9496 34546 9548 34552
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 9508 34241 9536 34546
rect 9494 34232 9550 34241
rect 9404 34196 9456 34202
rect 9494 34167 9550 34176
rect 9404 34138 9456 34144
rect 9402 33960 9458 33969
rect 9458 33930 9536 33946
rect 9458 33924 9548 33930
rect 9458 33918 9496 33924
rect 9402 33895 9458 33904
rect 9496 33866 9548 33872
rect 9404 33856 9456 33862
rect 9404 33798 9456 33804
rect 9416 33046 9444 33798
rect 9600 33658 9628 34546
rect 9772 34400 9824 34406
rect 9772 34342 9824 34348
rect 9784 34202 9812 34342
rect 9851 34300 10159 34309
rect 9851 34298 9857 34300
rect 9913 34298 9937 34300
rect 9993 34298 10017 34300
rect 10073 34298 10097 34300
rect 10153 34298 10159 34300
rect 9913 34246 9915 34298
rect 10095 34246 10097 34298
rect 9851 34244 9857 34246
rect 9913 34244 9937 34246
rect 9993 34244 10017 34246
rect 10073 34244 10097 34246
rect 10153 34244 10159 34246
rect 9851 34235 10159 34244
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9770 33552 9826 33561
rect 9770 33487 9772 33496
rect 9824 33487 9826 33496
rect 9864 33516 9916 33522
rect 9772 33458 9824 33464
rect 9864 33458 9916 33464
rect 9876 33300 9904 33458
rect 9784 33272 9904 33300
rect 9404 33040 9456 33046
rect 9404 32982 9456 32988
rect 9784 32910 9812 33272
rect 9851 33212 10159 33221
rect 9851 33210 9857 33212
rect 9913 33210 9937 33212
rect 9993 33210 10017 33212
rect 10073 33210 10097 33212
rect 10153 33210 10159 33212
rect 9913 33158 9915 33210
rect 10095 33158 10097 33210
rect 9851 33156 9857 33158
rect 9913 33156 9937 33158
rect 9993 33156 10017 33158
rect 10073 33156 10097 33158
rect 10153 33156 10159 33158
rect 9851 33147 10159 33156
rect 9772 32904 9824 32910
rect 9772 32846 9824 32852
rect 9494 32600 9550 32609
rect 9494 32535 9550 32544
rect 9312 31408 9364 31414
rect 9312 31350 9364 31356
rect 9404 31340 9456 31346
rect 9404 31282 9456 31288
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 9036 30932 9088 30938
rect 9036 30874 9088 30880
rect 9220 30728 9272 30734
rect 9218 30696 9220 30705
rect 9272 30696 9274 30705
rect 9218 30631 9274 30640
rect 9416 30433 9444 31282
rect 9402 30424 9458 30433
rect 9402 30359 9458 30368
rect 9036 30116 9088 30122
rect 9036 30058 9088 30064
rect 9048 29850 9076 30058
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 9048 29170 9076 29786
rect 9508 29753 9536 32535
rect 9680 31952 9732 31958
rect 9678 31920 9680 31929
rect 9732 31920 9734 31929
rect 9678 31855 9734 31864
rect 9784 31754 9812 32846
rect 10140 32836 10192 32842
rect 10140 32778 10192 32784
rect 10152 32570 10180 32778
rect 10140 32564 10192 32570
rect 10140 32506 10192 32512
rect 9851 32124 10159 32133
rect 9851 32122 9857 32124
rect 9913 32122 9937 32124
rect 9993 32122 10017 32124
rect 10073 32122 10097 32124
rect 10153 32122 10159 32124
rect 9913 32070 9915 32122
rect 10095 32070 10097 32122
rect 9851 32068 9857 32070
rect 9913 32068 9937 32070
rect 9993 32068 10017 32070
rect 10073 32068 10097 32070
rect 10153 32068 10159 32070
rect 9851 32059 10159 32068
rect 9692 31726 9812 31754
rect 9692 31090 9720 31726
rect 9772 31340 9824 31346
rect 9772 31282 9824 31288
rect 9784 31249 9812 31282
rect 9770 31240 9826 31249
rect 9770 31175 9826 31184
rect 9692 31062 9812 31090
rect 9784 30734 9812 31062
rect 9851 31036 10159 31045
rect 9851 31034 9857 31036
rect 9913 31034 9937 31036
rect 9993 31034 10017 31036
rect 10073 31034 10097 31036
rect 10153 31034 10159 31036
rect 9913 30982 9915 31034
rect 10095 30982 10097 31034
rect 9851 30980 9857 30982
rect 9913 30980 9937 30982
rect 9993 30980 10017 30982
rect 10073 30980 10097 30982
rect 10153 30980 10159 30982
rect 9851 30971 10159 30980
rect 10138 30832 10194 30841
rect 10138 30767 10194 30776
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9586 30424 9642 30433
rect 9586 30359 9642 30368
rect 9494 29744 9550 29753
rect 9494 29679 9550 29688
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9048 28994 9076 29106
rect 9048 28966 9444 28994
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9140 27674 9168 28154
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 9220 27532 9272 27538
rect 9220 27474 9272 27480
rect 8956 26846 9168 26874
rect 9140 26314 9168 26846
rect 9128 26308 9180 26314
rect 9128 26250 9180 26256
rect 9232 25838 9260 27474
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9324 26382 9352 26794
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 8852 25492 8904 25498
rect 8852 25434 8904 25440
rect 8852 25356 8904 25362
rect 8852 25298 8904 25304
rect 8864 24886 8892 25298
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 8760 24608 8812 24614
rect 8760 24550 8812 24556
rect 8772 23798 8800 24550
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8760 23792 8812 23798
rect 8760 23734 8812 23740
rect 8758 23624 8814 23633
rect 8758 23559 8814 23568
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8404 16998 8432 17614
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8392 16448 8444 16454
rect 8496 16436 8524 18226
rect 8444 16408 8524 16436
rect 8392 16390 8444 16396
rect 8312 16238 8432 16266
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8220 14906 8248 15574
rect 8220 14878 8340 14906
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14618 8248 14758
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8036 13802 8064 13942
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8036 12782 8064 13194
rect 7840 12776 7892 12782
rect 8024 12776 8076 12782
rect 7840 12718 7892 12724
rect 7930 12744 7986 12753
rect 8024 12718 8076 12724
rect 7930 12679 7986 12688
rect 7944 12442 7972 12679
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8036 12345 8064 12718
rect 8022 12336 8078 12345
rect 8022 12271 8078 12280
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8036 11898 8064 12174
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8022 11656 8078 11665
rect 7852 11614 8022 11642
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7760 4486 7788 11018
rect 7852 9722 7880 11614
rect 8022 11591 8078 11600
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7852 9489 7880 9522
rect 7838 9480 7894 9489
rect 7838 9415 7894 9424
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7852 8974 7880 9114
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 7852 7002 7880 8910
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4486 7880 4626
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7576 2746 7696 2774
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7484 2394 7512 2450
rect 7208 1834 7328 1850
rect 7196 1828 7328 1834
rect 7248 1822 7328 1828
rect 7392 2366 7512 2394
rect 7196 1770 7248 1776
rect 6552 1556 6604 1562
rect 6552 1498 6604 1504
rect 6736 1284 6788 1290
rect 6564 1244 6736 1272
rect 6460 1216 6512 1222
rect 6460 1158 6512 1164
rect 6368 672 6420 678
rect 6368 614 6420 620
rect 6564 160 6592 1244
rect 6736 1226 6788 1232
rect 7012 1284 7064 1290
rect 7064 1244 7328 1272
rect 7012 1226 7064 1232
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 6736 1012 6788 1018
rect 6736 954 6788 960
rect 6748 898 6776 954
rect 6920 944 6972 950
rect 6748 870 6868 898
rect 6972 892 7144 898
rect 6920 886 7144 892
rect 6932 870 7144 886
rect 6840 160 6868 870
rect 7116 160 7144 870
rect 7300 610 7328 1244
rect 7288 604 7340 610
rect 7288 546 7340 552
rect 7392 160 7420 2366
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 2106 7512 2246
rect 7576 2106 7604 2746
rect 7760 2514 7788 2994
rect 7944 2774 7972 11086
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 8498 8064 10406
rect 8128 9602 8156 14418
rect 8312 13818 8340 14878
rect 8220 13790 8340 13818
rect 8220 11558 8248 13790
rect 8404 13716 8432 16238
rect 8312 13688 8432 13716
rect 8482 13696 8538 13705
rect 8312 11694 8340 13688
rect 8482 13631 8538 13640
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8404 12889 8432 13398
rect 8390 12880 8446 12889
rect 8390 12815 8446 12824
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12220 8432 12718
rect 8496 12481 8524 13631
rect 8482 12472 8538 12481
rect 8482 12407 8538 12416
rect 8496 12374 8524 12407
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8404 12192 8524 12220
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8312 10606 8340 11630
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8496 9704 8524 12192
rect 8588 11762 8616 20402
rect 8680 18630 8708 21490
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8666 16688 8722 16697
rect 8666 16623 8668 16632
rect 8720 16623 8722 16632
rect 8668 16594 8720 16600
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8680 10810 8708 15914
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8404 9676 8524 9704
rect 8128 9574 8248 9602
rect 8404 9586 8432 9676
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8128 8634 8156 9386
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8128 7993 8156 8298
rect 8114 7984 8170 7993
rect 8114 7919 8170 7928
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8036 7342 8064 7754
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8036 5574 8064 7278
rect 8128 6254 8156 7919
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8022 4584 8078 4593
rect 8022 4519 8024 4528
rect 8076 4519 8078 4528
rect 8024 4490 8076 4496
rect 8128 2922 8156 6190
rect 8116 2916 8168 2922
rect 8116 2858 8168 2864
rect 7944 2746 8156 2774
rect 8128 2689 8156 2746
rect 8114 2680 8170 2689
rect 8114 2615 8170 2624
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7564 1216 7616 1222
rect 7564 1158 7616 1164
rect 7576 921 7604 1158
rect 7562 912 7618 921
rect 7562 847 7618 856
rect 7668 160 7696 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 1222 7788 2246
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 5170 54 5304 82
rect 5170 0 5226 54
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7852 82 7880 2382
rect 7930 2272 7986 2281
rect 7930 2207 7986 2216
rect 7944 1970 7972 2207
rect 8022 2000 8078 2009
rect 7932 1964 7984 1970
rect 8022 1935 8078 1944
rect 7932 1906 7984 1912
rect 8036 1834 8064 1935
rect 8024 1828 8076 1834
rect 8024 1770 8076 1776
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 7944 1018 7972 1158
rect 7932 1012 7984 1018
rect 7932 954 7984 960
rect 8036 950 8064 1294
rect 8024 944 8076 950
rect 8024 886 8076 892
rect 7930 82 7986 160
rect 7852 54 7986 82
rect 8128 82 8156 2382
rect 8220 2378 8248 9574
rect 8390 9580 8442 9586
rect 8390 9522 8442 9528
rect 8300 8492 8352 8498
rect 8300 8434 8352 8440
rect 8312 5098 8340 8434
rect 8404 8362 8432 9522
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 8838 8524 9454
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7546 8524 7686
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8588 6905 8616 10610
rect 8772 8401 8800 23559
rect 8956 23118 8984 24142
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8864 21146 8892 21490
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8956 21010 8984 23054
rect 9048 22030 9076 25162
rect 9232 24886 9260 25774
rect 9220 24880 9272 24886
rect 9220 24822 9272 24828
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9232 23322 9260 23666
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 9126 21720 9182 21729
rect 9126 21655 9182 21664
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8956 20874 8984 20946
rect 9140 20942 9168 21655
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 8944 20868 8996 20874
rect 8944 20810 8996 20816
rect 9128 20800 9180 20806
rect 9128 20742 9180 20748
rect 8850 20224 8906 20233
rect 8850 20159 8906 20168
rect 8864 16561 8892 20159
rect 9140 19786 9168 20742
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9140 19514 9168 19722
rect 9232 19514 9260 21490
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 8942 19000 8998 19009
rect 8942 18935 8998 18944
rect 8956 18358 8984 18935
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 9140 18426 9168 18770
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 9324 17678 9352 26318
rect 9416 25362 9444 28966
rect 9508 28529 9536 29106
rect 9600 29073 9628 30359
rect 9680 29640 9732 29646
rect 9680 29582 9732 29588
rect 9586 29064 9642 29073
rect 9586 28999 9642 29008
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9494 28520 9550 28529
rect 9600 28506 9628 28902
rect 9692 28626 9720 29582
rect 9784 28762 9812 30670
rect 10152 30258 10180 30767
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 9851 29948 10159 29957
rect 9851 29946 9857 29948
rect 9913 29946 9937 29948
rect 9993 29946 10017 29948
rect 10073 29946 10097 29948
rect 10153 29946 10159 29948
rect 9913 29894 9915 29946
rect 10095 29894 10097 29946
rect 9851 29892 9857 29894
rect 9913 29892 9937 29894
rect 9993 29892 10017 29894
rect 10073 29892 10097 29894
rect 10153 29892 10159 29894
rect 9851 29883 10159 29892
rect 10140 29708 10192 29714
rect 10140 29650 10192 29656
rect 10152 29345 10180 29650
rect 10138 29336 10194 29345
rect 10138 29271 10194 29280
rect 10244 28994 10272 43064
rect 10612 42906 10640 43114
rect 10968 43104 11020 43110
rect 10968 43046 11020 43052
rect 10600 42900 10652 42906
rect 10600 42842 10652 42848
rect 10784 42696 10836 42702
rect 10784 42638 10836 42644
rect 10324 42560 10376 42566
rect 10324 42502 10376 42508
rect 10336 42129 10364 42502
rect 10322 42120 10378 42129
rect 10322 42055 10378 42064
rect 10508 41676 10560 41682
rect 10508 41618 10560 41624
rect 10416 41132 10468 41138
rect 10416 41074 10468 41080
rect 10428 41041 10456 41074
rect 10414 41032 10470 41041
rect 10414 40967 10470 40976
rect 10324 40656 10376 40662
rect 10324 40598 10376 40604
rect 10336 40118 10364 40598
rect 10428 40508 10456 40967
rect 10520 40662 10548 41618
rect 10600 41540 10652 41546
rect 10600 41482 10652 41488
rect 10508 40656 10560 40662
rect 10508 40598 10560 40604
rect 10428 40480 10548 40508
rect 10324 40112 10376 40118
rect 10324 40054 10376 40060
rect 10336 37874 10364 40054
rect 10416 39840 10468 39846
rect 10416 39782 10468 39788
rect 10428 39370 10456 39782
rect 10416 39364 10468 39370
rect 10416 39306 10468 39312
rect 10520 39302 10548 40480
rect 10508 39296 10560 39302
rect 10508 39238 10560 39244
rect 10612 38842 10640 41482
rect 10796 41414 10824 42638
rect 10796 41386 10916 41414
rect 10784 40520 10836 40526
rect 10784 40462 10836 40468
rect 10796 40050 10824 40462
rect 10784 40044 10836 40050
rect 10784 39986 10836 39992
rect 10782 38856 10838 38865
rect 10612 38814 10782 38842
rect 10782 38791 10838 38800
rect 10324 37868 10376 37874
rect 10324 37810 10376 37816
rect 10336 35737 10364 37810
rect 10600 37664 10652 37670
rect 10600 37606 10652 37612
rect 10416 36712 10468 36718
rect 10416 36654 10468 36660
rect 10322 35728 10378 35737
rect 10322 35663 10378 35672
rect 10428 35578 10456 36654
rect 10612 36281 10640 37606
rect 10784 36644 10836 36650
rect 10784 36586 10836 36592
rect 10598 36272 10654 36281
rect 10598 36207 10654 36216
rect 10508 36168 10560 36174
rect 10508 36110 10560 36116
rect 10336 35550 10456 35578
rect 10336 33318 10364 35550
rect 10416 35488 10468 35494
rect 10416 35430 10468 35436
rect 10428 35290 10456 35430
rect 10416 35284 10468 35290
rect 10416 35226 10468 35232
rect 10416 35148 10468 35154
rect 10520 35136 10548 36110
rect 10796 35170 10824 36586
rect 10468 35108 10548 35136
rect 10704 35142 10824 35170
rect 10416 35090 10468 35096
rect 10704 34610 10732 35142
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10692 34604 10744 34610
rect 10692 34546 10744 34552
rect 10796 34241 10824 35022
rect 10782 34232 10838 34241
rect 10782 34167 10838 34176
rect 10692 34128 10744 34134
rect 10692 34070 10744 34076
rect 10784 34128 10836 34134
rect 10784 34070 10836 34076
rect 10324 33312 10376 33318
rect 10508 33312 10560 33318
rect 10376 33272 10456 33300
rect 10324 33254 10376 33260
rect 10428 32434 10456 33272
rect 10508 33254 10560 33260
rect 10520 32978 10548 33254
rect 10704 32978 10732 34070
rect 10508 32972 10560 32978
rect 10508 32914 10560 32920
rect 10692 32972 10744 32978
rect 10692 32914 10744 32920
rect 10600 32564 10652 32570
rect 10600 32506 10652 32512
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 10416 32428 10468 32434
rect 10416 32370 10468 32376
rect 10336 31958 10364 32370
rect 10508 32020 10560 32026
rect 10508 31962 10560 31968
rect 10324 31952 10376 31958
rect 10324 31894 10376 31900
rect 10416 31204 10468 31210
rect 10416 31146 10468 31152
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10336 29714 10364 31078
rect 10324 29708 10376 29714
rect 10324 29650 10376 29656
rect 10428 29646 10456 31146
rect 10520 31113 10548 31962
rect 10506 31104 10562 31113
rect 10506 31039 10562 31048
rect 10612 30954 10640 32506
rect 10704 31210 10732 32914
rect 10692 31204 10744 31210
rect 10692 31146 10744 31152
rect 10520 30926 10640 30954
rect 10520 29782 10548 30926
rect 10796 30841 10824 34070
rect 10782 30832 10838 30841
rect 10782 30767 10838 30776
rect 10692 30728 10744 30734
rect 10598 30696 10654 30705
rect 10692 30670 10744 30676
rect 10598 30631 10654 30640
rect 10508 29776 10560 29782
rect 10508 29718 10560 29724
rect 10612 29646 10640 30631
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10612 28994 10640 29582
rect 10244 28966 10456 28994
rect 9851 28860 10159 28869
rect 9851 28858 9857 28860
rect 9913 28858 9937 28860
rect 9993 28858 10017 28860
rect 10073 28858 10097 28860
rect 10153 28858 10159 28860
rect 9913 28806 9915 28858
rect 10095 28806 10097 28858
rect 9851 28804 9857 28806
rect 9913 28804 9937 28806
rect 9993 28804 10017 28806
rect 10073 28804 10097 28806
rect 10153 28804 10159 28806
rect 9851 28795 10159 28804
rect 9772 28756 9824 28762
rect 9772 28698 9824 28704
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9600 28478 9812 28506
rect 9494 28455 9550 28464
rect 9496 28416 9548 28422
rect 9496 28358 9548 28364
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9416 22982 9444 25298
rect 9508 24070 9536 28358
rect 9588 27532 9640 27538
rect 9588 27474 9640 27480
rect 9600 27130 9628 27474
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9586 26616 9642 26625
rect 9692 26602 9720 28358
rect 9784 27554 9812 28478
rect 10324 28416 10376 28422
rect 10324 28358 10376 28364
rect 10046 28248 10102 28257
rect 9968 28206 10046 28234
rect 9968 28082 9996 28206
rect 10046 28183 10102 28192
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9851 27772 10159 27781
rect 9851 27770 9857 27772
rect 9913 27770 9937 27772
rect 9993 27770 10017 27772
rect 10073 27770 10097 27772
rect 10153 27770 10159 27772
rect 9913 27718 9915 27770
rect 10095 27718 10097 27770
rect 9851 27716 9857 27718
rect 9913 27716 9937 27718
rect 9993 27716 10017 27718
rect 10073 27716 10097 27718
rect 10153 27716 10159 27718
rect 9851 27707 10159 27716
rect 9784 27526 9996 27554
rect 10336 27538 10364 28358
rect 9864 27464 9916 27470
rect 9864 27406 9916 27412
rect 9876 26908 9904 27406
rect 9968 27033 9996 27526
rect 10048 27532 10100 27538
rect 10324 27532 10376 27538
rect 10100 27492 10272 27520
rect 10048 27474 10100 27480
rect 10244 27418 10272 27492
rect 10324 27474 10376 27480
rect 10244 27390 10364 27418
rect 9954 27024 10010 27033
rect 9954 26959 10010 26968
rect 9876 26880 10272 26908
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9642 26574 9720 26602
rect 9586 26551 9642 26560
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9692 25770 9720 26454
rect 9784 25888 9812 26726
rect 9851 26684 10159 26693
rect 9851 26682 9857 26684
rect 9913 26682 9937 26684
rect 9993 26682 10017 26684
rect 10073 26682 10097 26684
rect 10153 26682 10159 26684
rect 9913 26630 9915 26682
rect 10095 26630 10097 26682
rect 9851 26628 9857 26630
rect 9913 26628 9937 26630
rect 9993 26628 10017 26630
rect 10073 26628 10097 26630
rect 10153 26628 10159 26630
rect 9851 26619 10159 26628
rect 10138 26480 10194 26489
rect 9968 26450 10138 26466
rect 9956 26444 10138 26450
rect 10008 26438 10138 26444
rect 10138 26415 10194 26424
rect 9956 26386 10008 26392
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10048 25900 10100 25906
rect 9784 25860 10048 25888
rect 10048 25842 10100 25848
rect 9588 25764 9640 25770
rect 9588 25706 9640 25712
rect 9680 25764 9732 25770
rect 9680 25706 9732 25712
rect 9600 25226 9628 25706
rect 9588 25220 9640 25226
rect 9588 25162 9640 25168
rect 9692 24682 9720 25706
rect 10152 25684 10180 26318
rect 9784 25656 10180 25684
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9496 24064 9548 24070
rect 9600 24041 9628 24142
rect 9496 24006 9548 24012
rect 9586 24032 9642 24041
rect 9586 23967 9642 23976
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 22098 9444 22918
rect 9586 22672 9642 22681
rect 9692 22642 9720 24346
rect 9784 23730 9812 25656
rect 9851 25596 10159 25605
rect 9851 25594 9857 25596
rect 9913 25594 9937 25596
rect 9993 25594 10017 25596
rect 10073 25594 10097 25596
rect 10153 25594 10159 25596
rect 9913 25542 9915 25594
rect 10095 25542 10097 25594
rect 9851 25540 9857 25542
rect 9913 25540 9937 25542
rect 9993 25540 10017 25542
rect 10073 25540 10097 25542
rect 10153 25540 10159 25542
rect 9851 25531 10159 25540
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 10152 24682 10180 25162
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 9851 24508 10159 24517
rect 9851 24506 9857 24508
rect 9913 24506 9937 24508
rect 9993 24506 10017 24508
rect 10073 24506 10097 24508
rect 10153 24506 10159 24508
rect 9913 24454 9915 24506
rect 10095 24454 10097 24506
rect 9851 24452 9857 24454
rect 9913 24452 9937 24454
rect 9993 24452 10017 24454
rect 10073 24452 10097 24454
rect 10153 24452 10159 24454
rect 9851 24443 10159 24452
rect 10048 24336 10100 24342
rect 10048 24278 10100 24284
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9968 23576 9996 23734
rect 10060 23662 10088 24278
rect 10138 24168 10194 24177
rect 10138 24103 10194 24112
rect 10152 23866 10180 24103
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9784 23548 9996 23576
rect 9586 22607 9642 22616
rect 9680 22636 9732 22642
rect 9496 22160 9548 22166
rect 9496 22102 9548 22108
rect 9404 22092 9456 22098
rect 9404 22034 9456 22040
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9416 21321 9444 21490
rect 9508 21468 9536 22102
rect 9600 21729 9628 22607
rect 9680 22578 9732 22584
rect 9784 22001 9812 23548
rect 9851 23420 10159 23429
rect 9851 23418 9857 23420
rect 9913 23418 9937 23420
rect 9993 23418 10017 23420
rect 10073 23418 10097 23420
rect 10153 23418 10159 23420
rect 9913 23366 9915 23418
rect 10095 23366 10097 23418
rect 9851 23364 9857 23366
rect 9913 23364 9937 23366
rect 9993 23364 10017 23366
rect 10073 23364 10097 23366
rect 10153 23364 10159 23366
rect 9851 23355 10159 23364
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 10060 22817 10088 22986
rect 10046 22808 10102 22817
rect 10046 22743 10102 22752
rect 9851 22332 10159 22341
rect 9851 22330 9857 22332
rect 9913 22330 9937 22332
rect 9993 22330 10017 22332
rect 10073 22330 10097 22332
rect 10153 22330 10159 22332
rect 9913 22278 9915 22330
rect 10095 22278 10097 22330
rect 9851 22276 9857 22278
rect 9913 22276 9937 22278
rect 9993 22276 10017 22278
rect 10073 22276 10097 22278
rect 10153 22276 10159 22278
rect 9851 22267 10159 22276
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9770 21992 9826 22001
rect 9770 21927 9826 21936
rect 9784 21894 9812 21927
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9586 21720 9642 21729
rect 9876 21706 9904 22034
rect 9586 21655 9642 21664
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9784 21678 9904 21706
rect 9588 21480 9640 21486
rect 9508 21440 9588 21468
rect 9588 21422 9640 21428
rect 9402 21312 9458 21321
rect 9402 21247 9458 21256
rect 9692 20806 9720 21626
rect 9784 21010 9812 21678
rect 9851 21244 10159 21253
rect 9851 21242 9857 21244
rect 9913 21242 9937 21244
rect 9993 21242 10017 21244
rect 10073 21242 10097 21244
rect 10153 21242 10159 21244
rect 9913 21190 9915 21242
rect 10095 21190 10097 21242
rect 9851 21188 9857 21190
rect 9913 21188 9937 21190
rect 9993 21188 10017 21190
rect 10073 21188 10097 21190
rect 10153 21188 10159 21190
rect 9851 21179 10159 21188
rect 9862 21040 9918 21049
rect 9772 21004 9824 21010
rect 9862 20975 9918 20984
rect 10138 21040 10194 21049
rect 10138 20975 10140 20984
rect 9772 20946 9824 20952
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9416 18766 9444 20266
rect 9784 20058 9812 20946
rect 9876 20942 9904 20975
rect 10192 20975 10194 20984
rect 10140 20946 10192 20952
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 9956 20528 10008 20534
rect 9954 20496 9956 20505
rect 10008 20496 10010 20505
rect 9954 20431 10010 20440
rect 10152 20380 10180 20742
rect 10244 20534 10272 26880
rect 10336 26450 10364 27390
rect 10428 26994 10456 28966
rect 10520 28966 10640 28994
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10336 25945 10364 26386
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10322 25936 10378 25945
rect 10322 25871 10378 25880
rect 10428 25838 10456 26318
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 10428 25498 10456 25774
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10152 20352 10272 20380
rect 9851 20156 10159 20165
rect 9851 20154 9857 20156
rect 9913 20154 9937 20156
rect 9993 20154 10017 20156
rect 10073 20154 10097 20156
rect 10153 20154 10159 20156
rect 9913 20102 9915 20154
rect 10095 20102 10097 20154
rect 9851 20100 9857 20102
rect 9913 20100 9937 20102
rect 9993 20100 10017 20102
rect 10073 20100 10097 20102
rect 10153 20100 10159 20102
rect 9851 20091 10159 20100
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9862 19952 9918 19961
rect 9784 19910 9862 19938
rect 9494 19408 9550 19417
rect 9494 19343 9550 19352
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9140 17105 9168 17274
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9126 17096 9182 17105
rect 9126 17031 9182 17040
rect 8850 16552 8906 16561
rect 8850 16487 8906 16496
rect 8864 14770 8892 16487
rect 9036 16108 9088 16114
rect 9232 16096 9260 17138
rect 9088 16068 9260 16096
rect 9036 16050 9088 16056
rect 9232 15638 9260 16068
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8864 14742 8984 14770
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8758 8392 8814 8401
rect 8758 8327 8814 8336
rect 8864 7410 8892 14554
rect 8956 12850 8984 14742
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 9048 12782 9076 15302
rect 9140 13394 9168 15438
rect 9232 15026 9260 15574
rect 9324 15366 9352 17614
rect 9402 15600 9458 15609
rect 9402 15535 9458 15544
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9416 15162 9444 15535
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9416 14414 9444 15098
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9508 14260 9536 19343
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18766 9720 19110
rect 9784 18766 9812 19910
rect 10244 19938 10272 20352
rect 9862 19887 9918 19896
rect 10152 19910 10272 19938
rect 10152 19174 10180 19910
rect 10230 19408 10286 19417
rect 10230 19343 10286 19352
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 9851 19068 10159 19077
rect 9851 19066 9857 19068
rect 9913 19066 9937 19068
rect 9993 19066 10017 19068
rect 10073 19066 10097 19068
rect 10153 19066 10159 19068
rect 9913 19014 9915 19066
rect 10095 19014 10097 19066
rect 9851 19012 9857 19014
rect 9913 19012 9937 19014
rect 9993 19012 10017 19014
rect 10073 19012 10097 19014
rect 10153 19012 10159 19014
rect 9851 19003 10159 19012
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9968 18578 9996 18634
rect 9692 18550 9996 18578
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 17377 9628 18158
rect 9586 17368 9642 17377
rect 9586 17303 9642 17312
rect 9600 17202 9628 17303
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16794 9628 17002
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9324 14232 9536 14260
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9140 12986 9168 13330
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9232 12850 9260 13670
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 9048 12170 9076 12718
rect 9324 12434 9352 14232
rect 9404 13932 9456 13938
rect 9600 13920 9628 16730
rect 9692 16046 9720 18550
rect 9851 17980 10159 17989
rect 9851 17978 9857 17980
rect 9913 17978 9937 17980
rect 9993 17978 10017 17980
rect 10073 17978 10097 17980
rect 10153 17978 10159 17980
rect 9913 17926 9915 17978
rect 10095 17926 10097 17978
rect 9851 17924 9857 17926
rect 9913 17924 9937 17926
rect 9993 17924 10017 17926
rect 10073 17924 10097 17926
rect 10153 17924 10159 17926
rect 9851 17915 10159 17924
rect 9772 17740 9824 17746
rect 10244 17728 10272 19343
rect 10336 18290 10364 22578
rect 10520 22094 10548 28966
rect 10704 28642 10732 30670
rect 10784 29776 10836 29782
rect 10784 29718 10836 29724
rect 10796 28994 10824 29718
rect 10888 29306 10916 41386
rect 10980 40730 11008 43046
rect 11164 42838 11192 43318
rect 11256 43314 11284 44463
rect 11532 43602 11560 44463
rect 11808 44146 11836 44463
rect 11808 44118 11928 44146
rect 11532 43574 11652 43602
rect 11244 43308 11296 43314
rect 11244 43250 11296 43256
rect 11244 43104 11296 43110
rect 11244 43046 11296 43052
rect 11152 42832 11204 42838
rect 11152 42774 11204 42780
rect 11256 41414 11284 43046
rect 11624 42702 11652 43574
rect 11900 42702 11928 44118
rect 12084 43314 12112 44463
rect 12360 43364 12388 44463
rect 12440 43376 12492 43382
rect 12360 43336 12440 43364
rect 12636 43364 12664 44463
rect 12912 43738 12940 44463
rect 13188 43874 13216 44463
rect 13188 43846 13308 43874
rect 12912 43710 13216 43738
rect 12818 43548 13126 43557
rect 12818 43546 12824 43548
rect 12880 43546 12904 43548
rect 12960 43546 12984 43548
rect 13040 43546 13064 43548
rect 13120 43546 13126 43548
rect 12880 43494 12882 43546
rect 13062 43494 13064 43546
rect 12818 43492 12824 43494
rect 12880 43492 12904 43494
rect 12960 43492 12984 43494
rect 13040 43492 13064 43494
rect 13120 43492 13126 43494
rect 12818 43483 13126 43492
rect 12808 43376 12860 43382
rect 12636 43336 12808 43364
rect 12440 43318 12492 43324
rect 13188 43364 13216 43710
rect 12808 43318 12860 43324
rect 12898 43344 12954 43353
rect 12072 43308 12124 43314
rect 12898 43279 12954 43288
rect 13004 43336 13216 43364
rect 13280 43364 13308 43846
rect 13360 43376 13412 43382
rect 13280 43336 13360 43364
rect 12072 43250 12124 43256
rect 12912 43110 12940 43279
rect 11980 43104 12032 43110
rect 11980 43046 12032 43052
rect 12532 43104 12584 43110
rect 12532 43046 12584 43052
rect 12900 43104 12952 43110
rect 12900 43046 12952 43052
rect 11612 42696 11664 42702
rect 11612 42638 11664 42644
rect 11888 42696 11940 42702
rect 11888 42638 11940 42644
rect 11796 42560 11848 42566
rect 11796 42502 11848 42508
rect 11704 42152 11756 42158
rect 11704 42094 11756 42100
rect 11256 41386 11468 41414
rect 11060 40928 11112 40934
rect 11060 40870 11112 40876
rect 10968 40724 11020 40730
rect 10968 40666 11020 40672
rect 11072 40594 11100 40870
rect 11060 40588 11112 40594
rect 11060 40530 11112 40536
rect 11152 40384 11204 40390
rect 11204 40332 11284 40338
rect 11152 40326 11284 40332
rect 11164 40310 11284 40326
rect 11256 39982 11284 40310
rect 11244 39976 11296 39982
rect 11244 39918 11296 39924
rect 11152 38344 11204 38350
rect 11152 38286 11204 38292
rect 11164 37942 11192 38286
rect 11152 37936 11204 37942
rect 11152 37878 11204 37884
rect 11256 37788 11284 39918
rect 11164 37760 11284 37788
rect 10968 37664 11020 37670
rect 10968 37606 11020 37612
rect 10980 33674 11008 37606
rect 11060 37120 11112 37126
rect 11060 37062 11112 37068
rect 11072 36378 11100 37062
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 11164 36122 11192 37760
rect 11242 36272 11298 36281
rect 11242 36207 11244 36216
rect 11296 36207 11298 36216
rect 11244 36178 11296 36184
rect 11336 36168 11388 36174
rect 11164 36116 11336 36122
rect 11164 36110 11388 36116
rect 11164 36094 11376 36110
rect 11060 35488 11112 35494
rect 11060 35430 11112 35436
rect 11072 35290 11100 35430
rect 11060 35284 11112 35290
rect 11060 35226 11112 35232
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 11072 34406 11100 35022
rect 11060 34400 11112 34406
rect 11060 34342 11112 34348
rect 10980 33646 11192 33674
rect 10968 33584 11020 33590
rect 10968 33526 11020 33532
rect 10980 30870 11008 33526
rect 11060 33448 11112 33454
rect 11060 33390 11112 33396
rect 11072 33114 11100 33390
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 11164 32994 11192 33646
rect 11072 32966 11192 32994
rect 10968 30864 11020 30870
rect 10968 30806 11020 30812
rect 10966 30696 11022 30705
rect 10966 30631 11022 30640
rect 10876 29300 10928 29306
rect 10876 29242 10928 29248
rect 10980 28994 11008 30631
rect 11072 30297 11100 32966
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 11256 32858 11284 36094
rect 11336 36032 11388 36038
rect 11336 35974 11388 35980
rect 11348 32978 11376 35974
rect 11336 32972 11388 32978
rect 11336 32914 11388 32920
rect 11164 32570 11192 32846
rect 11256 32830 11376 32858
rect 11242 32736 11298 32745
rect 11242 32671 11298 32680
rect 11152 32564 11204 32570
rect 11152 32506 11204 32512
rect 11152 31408 11204 31414
rect 11150 31376 11152 31385
rect 11204 31376 11206 31385
rect 11150 31311 11206 31320
rect 11256 30802 11284 32671
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11244 30796 11296 30802
rect 11244 30738 11296 30744
rect 11164 30394 11192 30738
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 11058 30288 11114 30297
rect 11058 30223 11114 30232
rect 11164 29782 11192 30330
rect 11244 30252 11296 30258
rect 11244 30194 11296 30200
rect 11256 30161 11284 30194
rect 11242 30152 11298 30161
rect 11242 30087 11298 30096
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 11348 29306 11376 32830
rect 11440 29594 11468 41386
rect 11716 41070 11744 42094
rect 11808 41993 11836 42502
rect 11794 41984 11850 41993
rect 11794 41919 11850 41928
rect 11704 41064 11756 41070
rect 11704 41006 11756 41012
rect 11612 40588 11664 40594
rect 11612 40530 11664 40536
rect 11624 39506 11652 40530
rect 11796 39840 11848 39846
rect 11796 39782 11848 39788
rect 11612 39500 11664 39506
rect 11612 39442 11664 39448
rect 11624 39030 11652 39442
rect 11704 39364 11756 39370
rect 11704 39306 11756 39312
rect 11612 39024 11664 39030
rect 11612 38966 11664 38972
rect 11520 38888 11572 38894
rect 11520 38830 11572 38836
rect 11532 37738 11560 38830
rect 11612 38480 11664 38486
rect 11612 38422 11664 38428
rect 11520 37732 11572 37738
rect 11520 37674 11572 37680
rect 11624 36038 11652 38422
rect 11612 36032 11664 36038
rect 11612 35974 11664 35980
rect 11518 35864 11574 35873
rect 11518 35799 11574 35808
rect 11532 35766 11560 35799
rect 11716 35766 11744 39306
rect 11808 38214 11836 39782
rect 11992 39001 12020 43046
rect 12544 42945 12572 43046
rect 12530 42936 12586 42945
rect 12530 42871 12586 42880
rect 12256 42764 12308 42770
rect 12256 42706 12308 42712
rect 12072 42560 12124 42566
rect 12072 42502 12124 42508
rect 12084 42129 12112 42502
rect 12070 42120 12126 42129
rect 12070 42055 12126 42064
rect 12268 41414 12296 42706
rect 13004 42702 13032 43336
rect 13360 43318 13412 43324
rect 13464 43296 13492 44463
rect 13636 43308 13688 43314
rect 13464 43268 13636 43296
rect 13636 43250 13688 43256
rect 13636 43172 13688 43178
rect 13636 43114 13688 43120
rect 12992 42696 13044 42702
rect 12992 42638 13044 42644
rect 13096 42634 13308 42650
rect 13084 42628 13308 42634
rect 13136 42622 13308 42628
rect 13084 42570 13136 42576
rect 12818 42460 13126 42469
rect 12818 42458 12824 42460
rect 12880 42458 12904 42460
rect 12960 42458 12984 42460
rect 13040 42458 13064 42460
rect 13120 42458 13126 42460
rect 12880 42406 12882 42458
rect 13062 42406 13064 42458
rect 12818 42404 12824 42406
rect 12880 42404 12904 42406
rect 12960 42404 12984 42406
rect 13040 42404 13064 42406
rect 13120 42404 13126 42406
rect 12818 42395 13126 42404
rect 12532 41812 12584 41818
rect 12532 41754 12584 41760
rect 12084 41386 12296 41414
rect 11978 38992 12034 39001
rect 11978 38927 12034 38936
rect 12084 38536 12112 41386
rect 12440 41200 12492 41206
rect 12440 41142 12492 41148
rect 12452 40458 12480 41142
rect 12440 40452 12492 40458
rect 12440 40394 12492 40400
rect 12164 40384 12216 40390
rect 12164 40326 12216 40332
rect 12348 40384 12400 40390
rect 12348 40326 12400 40332
rect 12176 39846 12204 40326
rect 12360 39982 12388 40326
rect 12348 39976 12400 39982
rect 12348 39918 12400 39924
rect 12164 39840 12216 39846
rect 12164 39782 12216 39788
rect 11900 38508 12112 38536
rect 11796 38208 11848 38214
rect 11796 38150 11848 38156
rect 11796 37664 11848 37670
rect 11796 37606 11848 37612
rect 11808 37398 11836 37606
rect 11796 37392 11848 37398
rect 11796 37334 11848 37340
rect 11900 35834 11928 38508
rect 12176 38418 12204 39782
rect 12256 39364 12308 39370
rect 12256 39306 12308 39312
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 12164 38412 12216 38418
rect 12164 38354 12216 38360
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 11992 35766 12020 38354
rect 12268 38332 12296 39306
rect 12452 38434 12480 40394
rect 12544 39030 12572 41754
rect 12818 41372 13126 41381
rect 12818 41370 12824 41372
rect 12880 41370 12904 41372
rect 12960 41370 12984 41372
rect 13040 41370 13064 41372
rect 13120 41370 13126 41372
rect 12880 41318 12882 41370
rect 13062 41318 13064 41370
rect 12818 41316 12824 41318
rect 12880 41316 12904 41318
rect 12960 41316 12984 41318
rect 13040 41316 13064 41318
rect 13120 41316 13126 41318
rect 12818 41307 13126 41316
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12728 40050 12756 40462
rect 12818 40284 13126 40293
rect 12818 40282 12824 40284
rect 12880 40282 12904 40284
rect 12960 40282 12984 40284
rect 13040 40282 13064 40284
rect 13120 40282 13126 40284
rect 12880 40230 12882 40282
rect 13062 40230 13064 40282
rect 12818 40228 12824 40230
rect 12880 40228 12904 40230
rect 12960 40228 12984 40230
rect 13040 40228 13064 40230
rect 13120 40228 13126 40230
rect 12818 40219 13126 40228
rect 12716 40044 12768 40050
rect 12716 39986 12768 39992
rect 12818 39196 13126 39205
rect 12818 39194 12824 39196
rect 12880 39194 12904 39196
rect 12960 39194 12984 39196
rect 13040 39194 13064 39196
rect 13120 39194 13126 39196
rect 12880 39142 12882 39194
rect 13062 39142 13064 39194
rect 12818 39140 12824 39142
rect 12880 39140 12904 39142
rect 12960 39140 12984 39142
rect 13040 39140 13064 39142
rect 13120 39140 13126 39142
rect 12818 39131 13126 39140
rect 12532 39024 12584 39030
rect 12532 38966 12584 38972
rect 12532 38752 12584 38758
rect 12532 38694 12584 38700
rect 12544 38554 12572 38694
rect 13280 38554 13308 42622
rect 13360 39976 13412 39982
rect 13360 39918 13412 39924
rect 13372 39642 13400 39918
rect 13360 39636 13412 39642
rect 13360 39578 13412 39584
rect 13452 39092 13504 39098
rect 13452 39034 13504 39040
rect 12532 38548 12584 38554
rect 12532 38490 12584 38496
rect 13268 38548 13320 38554
rect 13268 38490 13320 38496
rect 12452 38406 12572 38434
rect 12440 38344 12492 38350
rect 12268 38304 12440 38332
rect 12440 38286 12492 38292
rect 12164 38208 12216 38214
rect 12544 38196 12572 38406
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 12164 38150 12216 38156
rect 12452 38168 12572 38196
rect 12070 36952 12126 36961
rect 12070 36887 12126 36896
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11704 35760 11756 35766
rect 11704 35702 11756 35708
rect 11980 35760 12032 35766
rect 11980 35702 12032 35708
rect 11532 33386 11560 35702
rect 11612 35692 11664 35698
rect 11612 35634 11664 35640
rect 11624 35154 11652 35634
rect 11612 35148 11664 35154
rect 11612 35090 11664 35096
rect 11716 34626 11744 35702
rect 12084 35086 12112 36887
rect 12176 35766 12204 38150
rect 12254 37224 12310 37233
rect 12254 37159 12310 37168
rect 12268 36038 12296 37159
rect 12256 36032 12308 36038
rect 12256 35974 12308 35980
rect 12164 35760 12216 35766
rect 12164 35702 12216 35708
rect 12072 35080 12124 35086
rect 12070 35048 12072 35057
rect 12124 35048 12126 35057
rect 12070 34983 12126 34992
rect 11624 34598 11744 34626
rect 11624 34066 11652 34598
rect 11888 34536 11940 34542
rect 11888 34478 11940 34484
rect 11704 34468 11756 34474
rect 11704 34410 11756 34416
rect 11612 34060 11664 34066
rect 11612 34002 11664 34008
rect 11624 33658 11652 34002
rect 11612 33652 11664 33658
rect 11612 33594 11664 33600
rect 11520 33380 11572 33386
rect 11520 33322 11572 33328
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11532 30802 11560 32914
rect 11716 31498 11744 34410
rect 11900 34066 11928 34478
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 11796 33652 11848 33658
rect 11796 33594 11848 33600
rect 11624 31470 11744 31498
rect 11624 31414 11652 31470
rect 11612 31408 11664 31414
rect 11612 31350 11664 31356
rect 11808 31226 11836 33594
rect 11900 32978 11928 34002
rect 12176 33522 12204 35702
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 12164 33380 12216 33386
rect 12164 33322 12216 33328
rect 11888 32972 11940 32978
rect 11888 32914 11940 32920
rect 11980 32428 12032 32434
rect 11980 32370 12032 32376
rect 11624 31198 11836 31226
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 11532 30598 11560 30738
rect 11624 30705 11652 31198
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 11610 30696 11666 30705
rect 11610 30631 11666 30640
rect 11520 30592 11572 30598
rect 11520 30534 11572 30540
rect 11624 29714 11652 30631
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11440 29566 11652 29594
rect 11336 29300 11388 29306
rect 11336 29242 11388 29248
rect 11060 29232 11112 29238
rect 11058 29200 11060 29209
rect 11112 29200 11114 29209
rect 11058 29135 11114 29144
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11152 29028 11204 29034
rect 10796 28966 10916 28994
rect 10980 28966 11100 28994
rect 11152 28970 11204 28976
rect 10612 28614 10732 28642
rect 10612 25922 10640 28614
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10704 26042 10732 28494
rect 10888 28422 10916 28966
rect 11072 28642 11100 28966
rect 11164 28762 11192 28970
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 11072 28614 11192 28642
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10782 27432 10838 27441
rect 10782 27367 10784 27376
rect 10836 27367 10838 27376
rect 10784 27338 10836 27344
rect 10782 26480 10838 26489
rect 10782 26415 10784 26424
rect 10836 26415 10838 26424
rect 10784 26386 10836 26392
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10612 25894 10732 25922
rect 10598 24304 10654 24313
rect 10598 24239 10654 24248
rect 10428 22066 10548 22094
rect 10428 19281 10456 22066
rect 10612 20618 10640 24239
rect 10704 20806 10732 25894
rect 10888 25294 10916 28358
rect 10980 26586 11008 28494
rect 11164 28404 11192 28614
rect 11348 28558 11376 29106
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11440 28762 11468 28902
rect 11624 28762 11652 29566
rect 11428 28756 11480 28762
rect 11428 28698 11480 28704
rect 11612 28756 11664 28762
rect 11612 28698 11664 28704
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11164 28376 11376 28404
rect 11348 28082 11376 28376
rect 11624 28082 11652 28494
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11072 26450 11100 27814
rect 11244 26784 11296 26790
rect 11244 26726 11296 26732
rect 11152 26512 11204 26518
rect 11152 26454 11204 26460
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 11164 26042 11192 26454
rect 11256 26314 11284 26726
rect 11348 26489 11376 28018
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11334 26480 11390 26489
rect 11334 26415 11390 26424
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10796 22778 10824 24142
rect 10888 23905 10916 25230
rect 10968 24676 11020 24682
rect 10968 24618 11020 24624
rect 10874 23896 10930 23905
rect 10874 23831 10930 23840
rect 10874 23488 10930 23497
rect 10874 23423 10930 23432
rect 10888 23118 10916 23423
rect 10876 23112 10928 23118
rect 10876 23054 10928 23060
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 10980 22658 11008 24618
rect 11152 23656 11204 23662
rect 11152 23598 11204 23604
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 11072 22778 11100 23122
rect 11164 23050 11192 23598
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 11150 22944 11206 22953
rect 11150 22879 11206 22888
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10796 22630 11008 22658
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10612 20590 10732 20618
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10414 19272 10470 19281
rect 10414 19207 10470 19216
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10428 18766 10456 19110
rect 10520 18970 10548 20470
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10612 20058 10640 20402
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10598 19816 10654 19825
rect 10598 19751 10654 19760
rect 10612 19378 10640 19751
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10428 18057 10456 18566
rect 10508 18080 10560 18086
rect 10414 18048 10470 18057
rect 10508 18022 10560 18028
rect 10414 17983 10470 17992
rect 10520 17814 10548 18022
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10244 17700 10456 17728
rect 9772 17682 9824 17688
rect 9784 17338 9812 17682
rect 10140 17672 10192 17678
rect 10192 17632 10272 17660
rect 10140 17614 10192 17620
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9851 16892 10159 16901
rect 9851 16890 9857 16892
rect 9913 16890 9937 16892
rect 9993 16890 10017 16892
rect 10073 16890 10097 16892
rect 10153 16890 10159 16892
rect 9913 16838 9915 16890
rect 10095 16838 10097 16890
rect 9851 16836 9857 16838
rect 9913 16836 9937 16838
rect 9993 16836 10017 16838
rect 10073 16836 10097 16838
rect 10153 16836 10159 16838
rect 9851 16827 10159 16836
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15706 9720 15846
rect 9851 15804 10159 15813
rect 9851 15802 9857 15804
rect 9913 15802 9937 15804
rect 9993 15802 10017 15804
rect 10073 15802 10097 15804
rect 10153 15802 10159 15804
rect 9913 15750 9915 15802
rect 10095 15750 10097 15802
rect 9851 15748 9857 15750
rect 9913 15748 9937 15750
rect 9993 15748 10017 15750
rect 10073 15748 10097 15750
rect 10153 15748 10159 15750
rect 9851 15739 10159 15748
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9956 15564 10008 15570
rect 10008 15524 10088 15552
rect 9956 15506 10008 15512
rect 9692 15366 9720 15506
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9876 15178 9904 15438
rect 9954 15192 10010 15201
rect 9876 15150 9954 15178
rect 9954 15127 10010 15136
rect 10060 15042 10088 15524
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10244 15450 10272 17632
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10336 16794 10364 17138
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15570 10364 15846
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10152 15162 10180 15438
rect 10244 15422 10364 15450
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10060 15014 10272 15042
rect 9851 14716 10159 14725
rect 9851 14714 9857 14716
rect 9913 14714 9937 14716
rect 9993 14714 10017 14716
rect 10073 14714 10097 14716
rect 10153 14714 10159 14716
rect 9913 14662 9915 14714
rect 10095 14662 10097 14714
rect 9851 14660 9857 14662
rect 9913 14660 9937 14662
rect 9993 14660 10017 14662
rect 10073 14660 10097 14662
rect 10153 14660 10159 14662
rect 9851 14651 10159 14660
rect 10140 14544 10192 14550
rect 10140 14486 10192 14492
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 9784 14232 9996 14260
rect 10060 14249 10088 14350
rect 9784 14074 9812 14232
rect 9772 14068 9824 14074
rect 9968 14056 9996 14232
rect 10046 14240 10102 14249
rect 10046 14175 10102 14184
rect 10048 14068 10100 14074
rect 9968 14028 10048 14056
rect 9772 14010 9824 14016
rect 10048 14010 10100 14016
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9864 14000 9916 14006
rect 10152 13954 10180 14486
rect 9916 13948 10180 13954
rect 9864 13942 10180 13948
rect 9456 13892 9628 13920
rect 9404 13874 9456 13880
rect 9416 12866 9444 13874
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 13462 9536 13738
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12986 9536 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9416 12838 9536 12866
rect 9324 12406 9444 12434
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 10962 9076 11698
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9140 11150 9168 11494
rect 9324 11354 9352 11494
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9048 10934 9168 10962
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9042 9076 9862
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8942 8936 8998 8945
rect 8942 8871 8998 8880
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8956 7206 8984 8871
rect 9048 8430 9076 8978
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9034 7848 9090 7857
rect 9140 7834 9168 10934
rect 9416 10674 9444 12406
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9090 7806 9168 7834
rect 9232 7818 9260 10542
rect 9310 9616 9366 9625
rect 9310 9551 9312 9560
rect 9364 9551 9366 9560
rect 9404 9580 9456 9586
rect 9312 9522 9364 9528
rect 9404 9522 9456 9528
rect 9416 9382 9444 9522
rect 9404 9376 9456 9382
rect 9324 9336 9404 9364
rect 9220 7812 9272 7818
rect 9034 7783 9090 7792
rect 9220 7754 9272 7760
rect 9232 7410 9260 7754
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9324 7290 9352 9336
rect 9404 9318 9456 9324
rect 9402 8936 9458 8945
rect 9508 8922 9536 12838
rect 9692 12186 9720 13942
rect 9874 13926 10180 13942
rect 9851 13628 10159 13637
rect 9851 13626 9857 13628
rect 9913 13626 9937 13628
rect 9993 13626 10017 13628
rect 10073 13626 10097 13628
rect 10153 13626 10159 13628
rect 9913 13574 9915 13626
rect 10095 13574 10097 13626
rect 9851 13572 9857 13574
rect 9913 13572 9937 13574
rect 9993 13572 10017 13574
rect 10073 13572 10097 13574
rect 10153 13572 10159 13574
rect 9851 13563 10159 13572
rect 10244 13462 10272 15014
rect 10336 14362 10364 15422
rect 10428 14482 10456 17700
rect 10612 17270 10640 19314
rect 10704 18086 10732 20590
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10796 17882 10824 22630
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10874 21584 10930 21593
rect 10874 21519 10930 21528
rect 10888 19854 10916 21519
rect 10980 20890 11008 22374
rect 11058 21992 11114 22001
rect 11058 21927 11114 21936
rect 11072 21690 11100 21927
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11164 20942 11192 22879
rect 11256 22094 11284 26250
rect 11348 24818 11376 26415
rect 11336 24812 11388 24818
rect 11336 24754 11388 24760
rect 11334 24168 11390 24177
rect 11334 24103 11336 24112
rect 11388 24103 11390 24112
rect 11336 24074 11388 24080
rect 11440 23050 11468 27338
rect 11532 27130 11560 27406
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11532 25906 11560 27066
rect 11612 26988 11664 26994
rect 11612 26930 11664 26936
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 11532 24818 11560 25094
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11518 23216 11574 23225
rect 11518 23151 11574 23160
rect 11336 23044 11388 23050
rect 11336 22986 11388 22992
rect 11428 23044 11480 23050
rect 11428 22986 11480 22992
rect 11348 22545 11376 22986
rect 11440 22778 11468 22986
rect 11532 22982 11560 23151
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11334 22536 11390 22545
rect 11334 22471 11390 22480
rect 11256 22066 11468 22094
rect 11440 21978 11468 22066
rect 11256 21950 11468 21978
rect 11256 21894 11284 21950
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11152 20936 11204 20942
rect 10980 20874 11100 20890
rect 11152 20878 11204 20884
rect 10980 20868 11112 20874
rect 10980 20862 11060 20868
rect 11060 20810 11112 20816
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20398 11008 20742
rect 11256 20602 11284 21830
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10692 17672 10744 17678
rect 10888 17660 10916 18634
rect 11072 17882 11100 19178
rect 11164 18154 11192 20470
rect 11348 20398 11376 21422
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11336 20392 11388 20398
rect 11242 20360 11298 20369
rect 11336 20334 11388 20340
rect 11242 20295 11244 20304
rect 11296 20295 11298 20304
rect 11244 20266 11296 20272
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11348 19718 11376 20198
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11440 19417 11468 21286
rect 11520 20868 11572 20874
rect 11520 20810 11572 20816
rect 11426 19408 11482 19417
rect 11426 19343 11482 19352
rect 11532 19310 11560 20810
rect 11244 19304 11296 19310
rect 11520 19304 11572 19310
rect 11426 19272 11482 19281
rect 11244 19246 11296 19252
rect 11256 18766 11284 19246
rect 11348 19230 11426 19258
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11164 17746 11192 18090
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 10744 17632 10916 17660
rect 10692 17614 10744 17620
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 14550 10548 15846
rect 10612 15706 10640 16050
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10690 14920 10746 14929
rect 10690 14855 10746 14864
rect 10508 14544 10560 14550
rect 10508 14486 10560 14492
rect 10416 14476 10468 14482
rect 10416 14418 10468 14424
rect 10336 14334 10640 14362
rect 10414 14240 10470 14249
rect 10414 14175 10470 14184
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10336 13462 10364 14010
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10324 13456 10376 13462
rect 10324 13398 10376 13404
rect 9876 12850 9904 13398
rect 10140 13388 10192 13394
rect 10428 13376 10456 14175
rect 10428 13348 10548 13376
rect 10140 13330 10192 13336
rect 10152 13274 10180 13330
rect 10414 13288 10470 13297
rect 9956 13252 10008 13258
rect 10152 13246 10272 13274
rect 10008 13212 10088 13240
rect 9956 13194 10008 13200
rect 10060 13138 10088 13212
rect 10138 13152 10194 13161
rect 10060 13110 10138 13138
rect 10138 13087 10194 13096
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9851 12540 10159 12549
rect 9851 12538 9857 12540
rect 9913 12538 9937 12540
rect 9993 12538 10017 12540
rect 10073 12538 10097 12540
rect 10153 12538 10159 12540
rect 9913 12486 9915 12538
rect 10095 12486 10097 12538
rect 9851 12484 9857 12486
rect 9913 12484 9937 12486
rect 9993 12484 10017 12486
rect 10073 12484 10097 12486
rect 10153 12484 10159 12486
rect 9851 12475 10159 12484
rect 9692 12158 9812 12186
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11354 9720 12038
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9784 10810 9812 12158
rect 9851 11452 10159 11461
rect 9851 11450 9857 11452
rect 9913 11450 9937 11452
rect 9993 11450 10017 11452
rect 10073 11450 10097 11452
rect 10153 11450 10159 11452
rect 9913 11398 9915 11450
rect 10095 11398 10097 11450
rect 9851 11396 9857 11398
rect 9913 11396 9937 11398
rect 9993 11396 10017 11398
rect 10073 11396 10097 11398
rect 10153 11396 10159 11398
rect 9851 11387 10159 11396
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9876 11150 9904 11290
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9968 10656 9996 11086
rect 10152 10810 10180 11086
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 9692 10628 9996 10656
rect 9692 9625 9720 10628
rect 9851 10364 10159 10373
rect 9851 10362 9857 10364
rect 9913 10362 9937 10364
rect 9993 10362 10017 10364
rect 10073 10362 10097 10364
rect 10153 10362 10159 10364
rect 9913 10310 9915 10362
rect 10095 10310 10097 10362
rect 9851 10308 9857 10310
rect 9913 10308 9937 10310
rect 9993 10308 10017 10310
rect 10073 10308 10097 10310
rect 10153 10308 10159 10310
rect 9851 10299 10159 10308
rect 9770 10160 9826 10169
rect 9770 10095 9826 10104
rect 9678 9616 9734 9625
rect 9678 9551 9734 9560
rect 9588 9512 9640 9518
rect 9586 9480 9588 9489
rect 9640 9480 9642 9489
rect 9586 9415 9642 9424
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9178 9628 9318
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9458 8894 9536 8922
rect 9402 8871 9458 8880
rect 9692 7528 9720 9551
rect 9784 7993 9812 10095
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10152 9518 10180 9658
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 9851 9276 10159 9285
rect 9851 9274 9857 9276
rect 9913 9274 9937 9276
rect 9993 9274 10017 9276
rect 10073 9274 10097 9276
rect 10153 9274 10159 9276
rect 9913 9222 9915 9274
rect 10095 9222 10097 9274
rect 9851 9220 9857 9222
rect 9913 9220 9937 9222
rect 9993 9220 10017 9222
rect 10073 9220 10097 9222
rect 10153 9220 10159 9222
rect 9851 9211 10159 9220
rect 9851 8188 10159 8197
rect 9851 8186 9857 8188
rect 9913 8186 9937 8188
rect 9993 8186 10017 8188
rect 10073 8186 10097 8188
rect 10153 8186 10159 8188
rect 9913 8134 9915 8186
rect 10095 8134 10097 8186
rect 9851 8132 9857 8134
rect 9913 8132 9937 8134
rect 9993 8132 10017 8134
rect 10073 8132 10097 8134
rect 10153 8132 10159 8134
rect 9851 8123 10159 8132
rect 9770 7984 9826 7993
rect 9770 7919 9772 7928
rect 9824 7919 9826 7928
rect 9772 7890 9824 7896
rect 9140 7262 9352 7290
rect 9508 7500 9720 7528
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6934 9076 7142
rect 9036 6928 9088 6934
rect 8574 6896 8630 6905
rect 9036 6870 9088 6876
rect 8574 6831 8630 6840
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8680 5030 8708 6802
rect 8956 6458 8984 6802
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9048 6458 9076 6666
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8680 3466 8708 4014
rect 8864 3534 8892 4762
rect 9140 4282 9168 7262
rect 9220 7200 9272 7206
rect 9508 7154 9536 7500
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9220 7142 9272 7148
rect 9232 5302 9260 7142
rect 9416 7126 9536 7154
rect 9312 6792 9364 6798
rect 9416 6780 9444 7126
rect 9364 6752 9444 6780
rect 9312 6734 9364 6740
rect 9416 6254 9444 6752
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9310 6080 9366 6089
rect 9310 6015 9366 6024
rect 9324 5545 9352 6015
rect 9508 5914 9536 6122
rect 9496 5908 9548 5914
rect 9600 5896 9628 7346
rect 10244 7342 10272 13246
rect 10414 13223 10470 13232
rect 10324 9580 10376 9586
rect 10428 9568 10456 13223
rect 10520 12918 10548 13348
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10520 12345 10548 12854
rect 10506 12336 10562 12345
rect 10506 12271 10562 12280
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10520 9586 10548 9862
rect 10612 9722 10640 14334
rect 10704 13326 10732 14855
rect 10692 13320 10744 13326
rect 10690 13288 10692 13297
rect 10744 13288 10746 13297
rect 10690 13223 10746 13232
rect 10796 13138 10824 17274
rect 10704 13110 10824 13138
rect 10704 10062 10732 13110
rect 10888 12434 10916 17632
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10980 17338 11008 17614
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11058 17232 11114 17241
rect 11058 17167 11060 17176
rect 11112 17167 11114 17176
rect 11060 17138 11112 17144
rect 11256 16998 11284 18702
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 16794 11284 16934
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11348 16538 11376 19230
rect 11520 19246 11572 19252
rect 11426 19207 11482 19216
rect 11428 18692 11480 18698
rect 11428 18634 11480 18640
rect 11072 16510 11376 16538
rect 11072 14278 11100 16510
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 15094 11192 15438
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11152 15088 11204 15094
rect 11152 15030 11204 15036
rect 11164 14618 11192 15030
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11256 14482 11284 15370
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 13977 11192 14214
rect 11150 13968 11206 13977
rect 11150 13903 11206 13912
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10980 12986 11008 13262
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10888 12406 11008 12434
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10782 10296 10838 10305
rect 10782 10231 10838 10240
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10704 9926 10732 9998
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10376 9540 10456 9568
rect 10324 9522 10376 9528
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 8634 10364 9318
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 9851 7100 10159 7109
rect 9851 7098 9857 7100
rect 9913 7098 9937 7100
rect 9993 7098 10017 7100
rect 10073 7098 10097 7100
rect 10153 7098 10159 7100
rect 9913 7046 9915 7098
rect 10095 7046 10097 7098
rect 9851 7044 9857 7046
rect 9913 7044 9937 7046
rect 9993 7044 10017 7046
rect 10073 7044 10097 7046
rect 10153 7044 10159 7046
rect 9851 7035 10159 7044
rect 10336 6866 10364 7142
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9772 6248 9824 6254
rect 9876 6236 9904 6734
rect 9968 6322 9996 6734
rect 10428 6338 10456 9540
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 9178 10640 9522
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10704 8786 10732 9658
rect 9956 6316 10008 6322
rect 10060 6310 10456 6338
rect 10060 6304 10088 6310
rect 10008 6276 10088 6304
rect 9956 6258 10008 6264
rect 9824 6208 9904 6236
rect 10232 6248 10284 6254
rect 9772 6190 9824 6196
rect 10232 6190 10284 6196
rect 9600 5868 9720 5896
rect 9496 5850 9548 5856
rect 9692 5778 9720 5868
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9678 5672 9734 5681
rect 9678 5607 9734 5616
rect 9692 5574 9720 5607
rect 9680 5568 9732 5574
rect 9310 5536 9366 5545
rect 9680 5510 9732 5516
rect 9310 5471 9366 5480
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9232 4729 9260 5102
rect 9218 4720 9274 4729
rect 9218 4655 9274 4664
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9140 3890 9168 4218
rect 9312 4140 9364 4146
rect 9784 4128 9812 6190
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9968 5098 9996 5578
rect 10152 5574 10180 5646
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10244 5370 10272 6190
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 10244 4758 10272 5102
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9312 4082 9364 4088
rect 9416 4100 9812 4128
rect 9048 3862 9168 3890
rect 9048 3641 9076 3862
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9034 3632 9090 3641
rect 9034 3567 9036 3576
rect 9088 3567 9090 3576
rect 9036 3538 9088 3544
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8312 3194 8340 3402
rect 8300 3188 8352 3194
rect 9140 3176 9168 3674
rect 9140 3148 9260 3176
rect 8300 3130 8352 3136
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 8300 2848 8352 2854
rect 8576 2848 8628 2854
rect 8352 2796 8524 2802
rect 8300 2790 8524 2796
rect 8576 2790 8628 2796
rect 8312 2774 8524 2790
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8312 1970 8340 2586
rect 8404 2514 8432 2586
rect 8496 2514 8524 2774
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8588 2446 8616 2790
rect 8576 2440 8628 2446
rect 8944 2440 8996 2446
rect 8576 2382 8628 2388
rect 8772 2400 8944 2428
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8312 950 8340 1158
rect 8300 944 8352 950
rect 8300 886 8352 892
rect 8496 160 8524 2314
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8588 2106 8616 2246
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8668 1216 8720 1222
rect 8668 1158 8720 1164
rect 8680 882 8708 1158
rect 8668 876 8720 882
rect 8668 818 8720 824
rect 8772 160 8800 2400
rect 8944 2382 8996 2388
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 2106 8984 2246
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 8852 1488 8904 1494
rect 9036 1488 9088 1494
rect 8904 1436 9036 1442
rect 8852 1430 9088 1436
rect 8864 1414 9076 1430
rect 9036 1352 9088 1358
rect 9034 1320 9036 1329
rect 9088 1320 9090 1329
rect 9034 1255 9090 1264
rect 8206 82 8262 160
rect 8128 54 8262 82
rect 7930 0 7986 54
rect 8206 0 8262 54
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 82 9090 160
rect 9140 82 9168 2994
rect 9232 1290 9260 3148
rect 9324 2106 9352 4082
rect 9416 3942 9444 4100
rect 9876 4026 9904 4626
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 10060 4078 10088 4218
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 9508 3998 9904 4026
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9416 3738 9444 3878
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9508 3602 9536 3998
rect 9680 3936 9732 3942
rect 10060 3924 10088 4014
rect 9680 3878 9732 3884
rect 9784 3896 10088 3924
rect 9692 3777 9720 3878
rect 9678 3768 9734 3777
rect 9678 3703 9734 3712
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9678 3360 9734 3369
rect 9678 3295 9734 3304
rect 9692 3194 9720 3295
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9220 1284 9272 1290
rect 9220 1226 9272 1232
rect 9324 160 9352 1498
rect 9600 160 9628 2926
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9692 2446 9720 2586
rect 9784 2582 9812 3896
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 10048 3596 10100 3602
rect 10244 3584 10272 4150
rect 10336 4146 10364 4558
rect 10428 4146 10456 6310
rect 10612 8758 10732 8786
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10520 5817 10548 6122
rect 10612 5914 10640 8758
rect 10796 7886 10824 10231
rect 10888 10130 10916 10678
rect 10980 10169 11008 12406
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11354 11100 11562
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10966 10160 11022 10169
rect 10876 10124 10928 10130
rect 10966 10095 11022 10104
rect 10876 10066 10928 10072
rect 10888 9722 10916 10066
rect 10876 9716 10928 9722
rect 11164 9674 11192 13903
rect 11256 12714 11284 14418
rect 11440 14414 11468 18634
rect 11624 18426 11652 26930
rect 11716 26217 11744 31078
rect 11886 30560 11942 30569
rect 11886 30495 11942 30504
rect 11794 30288 11850 30297
rect 11794 30223 11850 30232
rect 11808 29238 11836 30223
rect 11796 29232 11848 29238
rect 11796 29174 11848 29180
rect 11794 29064 11850 29073
rect 11900 29034 11928 30495
rect 11992 29510 12020 32370
rect 12072 31680 12124 31686
rect 12072 31622 12124 31628
rect 12084 30802 12112 31622
rect 12072 30796 12124 30802
rect 12072 30738 12124 30744
rect 12084 29714 12112 30738
rect 12072 29708 12124 29714
rect 12072 29650 12124 29656
rect 11980 29504 12032 29510
rect 11980 29446 12032 29452
rect 11992 29102 12020 29446
rect 12176 29238 12204 33322
rect 12164 29232 12216 29238
rect 12164 29174 12216 29180
rect 11980 29096 12032 29102
rect 11980 29038 12032 29044
rect 11794 28999 11796 29008
rect 11848 28999 11850 29008
rect 11888 29028 11940 29034
rect 11796 28970 11848 28976
rect 11888 28970 11940 28976
rect 12072 28484 12124 28490
rect 12072 28426 12124 28432
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 11702 26208 11758 26217
rect 11702 26143 11758 26152
rect 11808 25401 11836 28018
rect 11900 26314 11928 28358
rect 12084 28257 12112 28426
rect 12070 28248 12126 28257
rect 12070 28183 12126 28192
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 11886 26072 11942 26081
rect 11886 26007 11942 26016
rect 11900 25974 11928 26007
rect 11888 25968 11940 25974
rect 11888 25910 11940 25916
rect 11794 25392 11850 25401
rect 11794 25327 11850 25336
rect 11704 25220 11756 25226
rect 11704 25162 11756 25168
rect 11716 24682 11744 25162
rect 11808 24750 11836 25327
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11704 24676 11756 24682
rect 11704 24618 11756 24624
rect 11900 24313 11928 25910
rect 12084 25158 12112 27950
rect 12164 27940 12216 27946
rect 12164 27882 12216 27888
rect 12072 25152 12124 25158
rect 11978 25120 12034 25129
rect 12072 25094 12124 25100
rect 11978 25055 12034 25064
rect 11886 24304 11942 24313
rect 11886 24239 11942 24248
rect 11992 23866 12020 25055
rect 12176 24886 12204 27882
rect 12268 27470 12296 35974
rect 12452 35873 12480 38168
rect 12636 38010 12664 38286
rect 12818 38108 13126 38117
rect 12818 38106 12824 38108
rect 12880 38106 12904 38108
rect 12960 38106 12984 38108
rect 13040 38106 13064 38108
rect 13120 38106 13126 38108
rect 12880 38054 12882 38106
rect 13062 38054 13064 38106
rect 12818 38052 12824 38054
rect 12880 38052 12904 38054
rect 12960 38052 12984 38054
rect 13040 38052 13064 38054
rect 13120 38052 13126 38054
rect 12818 38043 13126 38052
rect 12624 38004 12676 38010
rect 12624 37946 12676 37952
rect 12818 37020 13126 37029
rect 12818 37018 12824 37020
rect 12880 37018 12904 37020
rect 12960 37018 12984 37020
rect 13040 37018 13064 37020
rect 13120 37018 13126 37020
rect 12880 36966 12882 37018
rect 13062 36966 13064 37018
rect 12818 36964 12824 36966
rect 12880 36964 12904 36966
rect 12960 36964 12984 36966
rect 13040 36964 13064 36966
rect 13120 36964 13126 36966
rect 12818 36955 13126 36964
rect 12532 36576 12584 36582
rect 12532 36518 12584 36524
rect 12544 36242 12572 36518
rect 12532 36236 12584 36242
rect 12532 36178 12584 36184
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12438 35864 12494 35873
rect 12438 35799 12494 35808
rect 12636 35698 12664 35974
rect 12818 35932 13126 35941
rect 12818 35930 12824 35932
rect 12880 35930 12904 35932
rect 12960 35930 12984 35932
rect 13040 35930 13064 35932
rect 13120 35930 13126 35932
rect 12880 35878 12882 35930
rect 13062 35878 13064 35930
rect 12818 35876 12824 35878
rect 12880 35876 12904 35878
rect 12960 35876 12984 35878
rect 13040 35876 13064 35878
rect 13120 35876 13126 35878
rect 12818 35867 13126 35876
rect 12624 35692 12676 35698
rect 12624 35634 12676 35640
rect 12808 35624 12860 35630
rect 12808 35566 12860 35572
rect 12990 35592 13046 35601
rect 12820 35290 12848 35566
rect 12990 35527 12992 35536
rect 13044 35527 13046 35536
rect 12992 35498 13044 35504
rect 13464 35465 13492 39034
rect 13544 37868 13596 37874
rect 13544 37810 13596 37816
rect 13450 35456 13506 35465
rect 13450 35391 13506 35400
rect 13556 35290 13584 37810
rect 12808 35284 12860 35290
rect 12808 35226 12860 35232
rect 13544 35284 13596 35290
rect 13544 35226 13596 35232
rect 13358 35184 13414 35193
rect 13358 35119 13414 35128
rect 12818 34844 13126 34853
rect 12818 34842 12824 34844
rect 12880 34842 12904 34844
rect 12960 34842 12984 34844
rect 13040 34842 13064 34844
rect 13120 34842 13126 34844
rect 12880 34790 12882 34842
rect 13062 34790 13064 34842
rect 12818 34788 12824 34790
rect 12880 34788 12904 34790
rect 12960 34788 12984 34790
rect 13040 34788 13064 34790
rect 13120 34788 13126 34790
rect 12818 34779 13126 34788
rect 13266 34776 13322 34785
rect 13266 34711 13322 34720
rect 13082 34504 13138 34513
rect 13138 34462 13216 34490
rect 13082 34439 13138 34448
rect 12530 34096 12586 34105
rect 12530 34031 12532 34040
rect 12584 34031 12586 34040
rect 12532 34002 12584 34008
rect 12346 33960 12402 33969
rect 12346 33895 12348 33904
rect 12400 33895 12402 33904
rect 12530 33960 12586 33969
rect 12586 33930 12664 33946
rect 12586 33924 12676 33930
rect 12586 33918 12624 33924
rect 12530 33895 12586 33904
rect 12348 33866 12400 33872
rect 12624 33866 12676 33872
rect 12818 33756 13126 33765
rect 12818 33754 12824 33756
rect 12880 33754 12904 33756
rect 12960 33754 12984 33756
rect 13040 33754 13064 33756
rect 13120 33754 13126 33756
rect 12880 33702 12882 33754
rect 13062 33702 13064 33754
rect 12818 33700 12824 33702
rect 12880 33700 12904 33702
rect 12960 33700 12984 33702
rect 13040 33700 13064 33702
rect 13120 33700 13126 33702
rect 12818 33691 13126 33700
rect 12716 33652 12768 33658
rect 12716 33594 12768 33600
rect 12728 33522 12756 33594
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 12900 33312 12952 33318
rect 12900 33254 12952 33260
rect 12912 33114 12940 33254
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12440 31340 12492 31346
rect 12440 31282 12492 31288
rect 12348 30592 12400 30598
rect 12348 30534 12400 30540
rect 12360 29714 12388 30534
rect 12452 30054 12480 31282
rect 12544 30938 12572 31758
rect 12636 31521 12664 32846
rect 12716 32836 12768 32842
rect 12716 32778 12768 32784
rect 12622 31512 12678 31521
rect 12622 31447 12678 31456
rect 12728 31464 12756 32778
rect 12818 32668 13126 32677
rect 12818 32666 12824 32668
rect 12880 32666 12904 32668
rect 12960 32666 12984 32668
rect 13040 32666 13064 32668
rect 13120 32666 13126 32668
rect 12880 32614 12882 32666
rect 13062 32614 13064 32666
rect 12818 32612 12824 32614
rect 12880 32612 12904 32614
rect 12960 32612 12984 32614
rect 13040 32612 13064 32614
rect 13120 32612 13126 32614
rect 12818 32603 13126 32612
rect 12818 31580 13126 31589
rect 12818 31578 12824 31580
rect 12880 31578 12904 31580
rect 12960 31578 12984 31580
rect 13040 31578 13064 31580
rect 13120 31578 13126 31580
rect 12880 31526 12882 31578
rect 13062 31526 13064 31578
rect 12818 31524 12824 31526
rect 12880 31524 12904 31526
rect 12960 31524 12984 31526
rect 13040 31524 13064 31526
rect 13120 31524 13126 31526
rect 12818 31515 13126 31524
rect 13188 31464 13216 34462
rect 13280 31958 13308 34711
rect 13268 31952 13320 31958
rect 13268 31894 13320 31900
rect 12728 31436 12848 31464
rect 12820 31346 12848 31436
rect 13096 31436 13216 31464
rect 12808 31340 12860 31346
rect 12808 31282 12860 31288
rect 12622 31240 12678 31249
rect 12622 31175 12678 31184
rect 12532 30932 12584 30938
rect 12532 30874 12584 30880
rect 12636 30433 12664 31175
rect 13096 30580 13124 31436
rect 13280 31346 13308 31894
rect 13268 31340 13320 31346
rect 13268 31282 13320 31288
rect 13188 31210 13308 31226
rect 13188 31204 13320 31210
rect 13188 31198 13268 31204
rect 13188 30870 13216 31198
rect 13268 31146 13320 31152
rect 13266 31104 13322 31113
rect 13266 31039 13322 31048
rect 13176 30864 13228 30870
rect 13176 30806 13228 30812
rect 13096 30552 13216 30580
rect 12818 30492 13126 30501
rect 12818 30490 12824 30492
rect 12880 30490 12904 30492
rect 12960 30490 12984 30492
rect 13040 30490 13064 30492
rect 13120 30490 13126 30492
rect 12880 30438 12882 30490
rect 13062 30438 13064 30490
rect 12818 30436 12824 30438
rect 12880 30436 12904 30438
rect 12960 30436 12984 30438
rect 13040 30436 13064 30438
rect 13120 30436 13126 30438
rect 12622 30424 12678 30433
rect 12818 30427 13126 30436
rect 12622 30359 12678 30368
rect 12440 30048 12492 30054
rect 12440 29990 12492 29996
rect 12348 29708 12400 29714
rect 12348 29650 12400 29656
rect 12452 29170 12480 29990
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12728 29084 12756 29582
rect 12818 29404 13126 29413
rect 12818 29402 12824 29404
rect 12880 29402 12904 29404
rect 12960 29402 12984 29404
rect 13040 29402 13064 29404
rect 13120 29402 13126 29404
rect 12880 29350 12882 29402
rect 13062 29350 13064 29402
rect 12818 29348 12824 29350
rect 12880 29348 12904 29350
rect 12960 29348 12984 29350
rect 13040 29348 13064 29350
rect 13120 29348 13126 29350
rect 12818 29339 13126 29348
rect 12544 29056 12756 29084
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12452 28121 12480 28970
rect 12544 28937 12572 29056
rect 12624 29006 12676 29012
rect 13188 28994 13216 30552
rect 12676 28966 12756 28994
rect 12624 28948 12676 28954
rect 12530 28928 12586 28937
rect 12530 28863 12586 28872
rect 12438 28112 12494 28121
rect 12438 28047 12494 28056
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12348 26308 12400 26314
rect 12348 26250 12400 26256
rect 12268 26042 12296 26250
rect 12256 26036 12308 26042
rect 12256 25978 12308 25984
rect 12268 25158 12296 25978
rect 12360 25838 12388 26250
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 12360 25294 12388 25638
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12452 25226 12480 27270
rect 12544 26042 12572 28863
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12636 26926 12664 27950
rect 12728 27520 12756 28966
rect 13096 28966 13216 28994
rect 13096 28422 13124 28966
rect 13280 28642 13308 31039
rect 13188 28614 13308 28642
rect 13084 28416 13136 28422
rect 13084 28358 13136 28364
rect 12818 28316 13126 28325
rect 12818 28314 12824 28316
rect 12880 28314 12904 28316
rect 12960 28314 12984 28316
rect 13040 28314 13064 28316
rect 13120 28314 13126 28316
rect 12880 28262 12882 28314
rect 13062 28262 13064 28314
rect 12818 28260 12824 28262
rect 12880 28260 12904 28262
rect 12960 28260 12984 28262
rect 13040 28260 13064 28262
rect 13120 28260 13126 28262
rect 12818 28251 13126 28260
rect 12808 27532 12860 27538
rect 12728 27492 12808 27520
rect 12728 27130 12756 27492
rect 12808 27474 12860 27480
rect 13188 27441 13216 28614
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 13174 27432 13230 27441
rect 13174 27367 13230 27376
rect 13280 27316 13308 28358
rect 13188 27288 13308 27316
rect 12818 27228 13126 27237
rect 12818 27226 12824 27228
rect 12880 27226 12904 27228
rect 12960 27226 12984 27228
rect 13040 27226 13064 27228
rect 13120 27226 13126 27228
rect 12880 27174 12882 27226
rect 13062 27174 13064 27226
rect 12818 27172 12824 27174
rect 12880 27172 12904 27174
rect 12960 27172 12984 27174
rect 13040 27172 13064 27174
rect 13120 27172 13126 27174
rect 12818 27163 13126 27172
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12544 25362 12572 25638
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12636 25226 12664 26182
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12360 24970 12388 25094
rect 12728 24970 12756 26930
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12912 26586 12940 26862
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12818 26140 13126 26149
rect 12818 26138 12824 26140
rect 12880 26138 12904 26140
rect 12960 26138 12984 26140
rect 13040 26138 13064 26140
rect 13120 26138 13126 26140
rect 12880 26086 12882 26138
rect 13062 26086 13064 26138
rect 12818 26084 12824 26086
rect 12880 26084 12904 26086
rect 12960 26084 12984 26086
rect 13040 26084 13064 26086
rect 13120 26084 13126 26086
rect 12818 26075 13126 26084
rect 12818 25052 13126 25061
rect 12818 25050 12824 25052
rect 12880 25050 12904 25052
rect 12960 25050 12984 25052
rect 13040 25050 13064 25052
rect 13120 25050 13126 25052
rect 12880 24998 12882 25050
rect 13062 24998 13064 25050
rect 12818 24996 12824 24998
rect 12880 24996 12904 24998
rect 12960 24996 12984 24998
rect 13040 24996 13064 24998
rect 13120 24996 13126 24998
rect 12818 24987 13126 24996
rect 12268 24954 12388 24970
rect 12256 24948 12388 24954
rect 12308 24942 12388 24948
rect 12636 24942 12756 24970
rect 12256 24890 12308 24896
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 12072 24744 12124 24750
rect 12072 24686 12124 24692
rect 12084 24274 12112 24686
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 12176 24154 12204 24822
rect 12348 24200 12400 24206
rect 12176 24126 12296 24154
rect 12636 24177 12664 24942
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12348 24142 12400 24148
rect 12622 24168 12678 24177
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11716 21978 11744 23666
rect 11808 23338 11836 23734
rect 12070 23624 12126 23633
rect 12070 23559 12126 23568
rect 12084 23526 12112 23559
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11808 23310 12112 23338
rect 11796 23044 11848 23050
rect 11796 22986 11848 22992
rect 11808 22817 11836 22986
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11794 22808 11850 22817
rect 11794 22743 11850 22752
rect 11716 21962 11836 21978
rect 11716 21956 11848 21962
rect 11716 21950 11796 21956
rect 11716 21457 11744 21950
rect 11796 21898 11848 21904
rect 11796 21480 11848 21486
rect 11702 21448 11758 21457
rect 11796 21422 11848 21428
rect 11702 21383 11758 21392
rect 11808 21049 11836 21422
rect 11794 21040 11850 21049
rect 11794 20975 11796 20984
rect 11848 20975 11850 20984
rect 11796 20946 11848 20952
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11808 19378 11836 20470
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11518 17776 11574 17785
rect 11518 17711 11574 17720
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11242 12336 11298 12345
rect 11242 12271 11298 12280
rect 11256 12102 11284 12271
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 9722 11284 10610
rect 10876 9658 10928 9664
rect 10980 9646 11192 9674
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10506 5808 10562 5817
rect 10506 5743 10562 5752
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10100 3556 10272 3584
rect 10048 3538 10100 3544
rect 9954 3496 10010 3505
rect 9954 3431 10010 3440
rect 9864 3120 9916 3126
rect 9968 3108 9996 3431
rect 10336 3126 10364 3878
rect 10428 3194 10456 4082
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 9916 3080 9996 3108
rect 10324 3120 10376 3126
rect 9864 3062 9916 3068
rect 10324 3062 10376 3068
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10322 2272 10378 2281
rect 9692 1358 9720 2246
rect 10322 2207 10378 2216
rect 10336 1970 10364 2207
rect 10520 2106 10548 3538
rect 10612 2446 10640 5850
rect 10888 5302 10916 8570
rect 10980 8537 11008 9646
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 10966 8528 11022 8537
rect 10966 8463 11022 8472
rect 10980 7410 11008 8463
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 11072 7274 11100 9415
rect 11152 8424 11204 8430
rect 11152 8366 11204 8372
rect 11164 8090 11192 8366
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11256 8090 11284 8230
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11242 7032 11298 7041
rect 11242 6967 11298 6976
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10966 5944 11022 5953
rect 10966 5879 11022 5888
rect 10980 5574 11008 5879
rect 11072 5574 11100 6054
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10888 4622 10916 5238
rect 11164 5098 11192 5646
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11164 4758 11192 5034
rect 11152 4752 11204 4758
rect 11152 4694 11204 4700
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 11058 3768 11114 3777
rect 11058 3703 11060 3712
rect 11112 3703 11114 3712
rect 11152 3732 11204 3738
rect 11060 3674 11112 3680
rect 11152 3674 11204 3680
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10704 3369 10732 3402
rect 10690 3360 10746 3369
rect 10690 3295 10746 3304
rect 11060 3120 11112 3126
rect 11058 3088 11060 3097
rect 11112 3088 11114 3097
rect 10692 3052 10744 3058
rect 11058 3023 11114 3032
rect 10692 2994 10744 3000
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10508 2100 10560 2106
rect 10508 2042 10560 2048
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 10704 1562 10732 2994
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10796 2650 10824 2926
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11060 1760 11112 1766
rect 10980 1720 11060 1748
rect 10692 1556 10744 1562
rect 10692 1498 10744 1504
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9864 672 9916 678
rect 9864 614 9916 620
rect 9968 626 9996 1362
rect 10508 1216 10560 1222
rect 10508 1158 10560 1164
rect 9876 160 9904 614
rect 9968 598 10180 626
rect 10152 160 10180 598
rect 9034 54 9168 82
rect 9034 0 9090 54
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 82 10470 160
rect 10520 82 10548 1158
rect 10692 1012 10744 1018
rect 10692 954 10744 960
rect 10704 160 10732 954
rect 10980 160 11008 1720
rect 11060 1702 11112 1708
rect 11164 746 11192 3674
rect 11256 2650 11284 6967
rect 11348 5624 11376 12786
rect 11532 12434 11560 17711
rect 11624 15162 11652 18362
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 17134 11744 18022
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11808 15162 11836 19314
rect 11900 15450 11928 22918
rect 12084 21962 12112 23310
rect 12176 23118 12204 24006
rect 12268 23730 12296 24126
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12360 23322 12388 24142
rect 12622 24103 12678 24112
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12256 22772 12308 22778
rect 12256 22714 12308 22720
rect 12268 22250 12296 22714
rect 12360 22438 12388 23258
rect 12348 22432 12400 22438
rect 12348 22374 12400 22380
rect 12268 22222 12388 22250
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 12072 21956 12124 21962
rect 12072 21898 12124 21904
rect 11992 21690 12020 21898
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11992 20058 12020 20946
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12176 19334 12204 20878
rect 12256 20392 12308 20398
rect 12256 20334 12308 20340
rect 12084 19306 12204 19334
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 16658 12020 18566
rect 12084 17542 12112 19306
rect 12268 18714 12296 20334
rect 12360 19417 12388 22222
rect 12452 20534 12480 23802
rect 12636 23730 12664 24103
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12544 20602 12572 23598
rect 12622 23080 12678 23089
rect 12622 23015 12678 23024
rect 12636 22642 12664 23015
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12636 21554 12664 22374
rect 12728 21672 12756 24822
rect 13188 24698 13216 27288
rect 13268 26852 13320 26858
rect 13268 26794 13320 26800
rect 13280 25906 13308 26794
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13096 24670 13216 24698
rect 13096 24410 13124 24670
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 12818 23964 13126 23973
rect 12818 23962 12824 23964
rect 12880 23962 12904 23964
rect 12960 23962 12984 23964
rect 13040 23962 13064 23964
rect 13120 23962 13126 23964
rect 12880 23910 12882 23962
rect 13062 23910 13064 23962
rect 12818 23908 12824 23910
rect 12880 23908 12904 23910
rect 12960 23908 12984 23910
rect 13040 23908 13064 23910
rect 13120 23908 13126 23910
rect 12818 23899 13126 23908
rect 13188 23662 13216 24550
rect 13176 23656 13228 23662
rect 13280 23633 13308 25638
rect 13176 23598 13228 23604
rect 13266 23624 13322 23633
rect 13266 23559 13322 23568
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 12818 22876 13126 22885
rect 12818 22874 12824 22876
rect 12880 22874 12904 22876
rect 12960 22874 12984 22876
rect 13040 22874 13064 22876
rect 13120 22874 13126 22876
rect 12880 22822 12882 22874
rect 13062 22822 13064 22874
rect 12818 22820 12824 22822
rect 12880 22820 12904 22822
rect 12960 22820 12984 22822
rect 13040 22820 13064 22822
rect 13120 22820 13126 22822
rect 12818 22811 13126 22820
rect 13176 22704 13228 22710
rect 13176 22646 13228 22652
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12912 22234 12940 22578
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 12818 21788 13126 21797
rect 12818 21786 12824 21788
rect 12880 21786 12904 21788
rect 12960 21786 12984 21788
rect 13040 21786 13064 21788
rect 13120 21786 13126 21788
rect 12880 21734 12882 21786
rect 13062 21734 13064 21786
rect 12818 21732 12824 21734
rect 12880 21732 12904 21734
rect 12960 21732 12984 21734
rect 13040 21732 13064 21734
rect 13120 21732 13126 21734
rect 12818 21723 13126 21732
rect 12728 21644 12848 21672
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12636 20777 12664 20810
rect 12716 20800 12768 20806
rect 12622 20768 12678 20777
rect 12820 20788 12848 21644
rect 13188 20913 13216 22646
rect 13174 20904 13230 20913
rect 13174 20839 13230 20848
rect 12820 20760 13216 20788
rect 12716 20742 12768 20748
rect 12622 20703 12678 20712
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12728 20398 12756 20742
rect 12818 20700 13126 20709
rect 12818 20698 12824 20700
rect 12880 20698 12904 20700
rect 12960 20698 12984 20700
rect 13040 20698 13064 20700
rect 13120 20698 13126 20700
rect 12880 20646 12882 20698
rect 13062 20646 13064 20698
rect 12818 20644 12824 20646
rect 12880 20644 12904 20646
rect 12960 20644 12984 20646
rect 13040 20644 13064 20646
rect 13120 20644 13126 20646
rect 12818 20635 13126 20644
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12530 19952 12586 19961
rect 12452 19910 12530 19938
rect 12346 19408 12402 19417
rect 12346 19343 12402 19352
rect 12176 18686 12296 18714
rect 12176 18290 12204 18686
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 18358 12296 18566
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12176 17898 12204 18226
rect 12176 17870 12296 17898
rect 12268 17814 12296 17870
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12084 16114 12112 17070
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 12084 15570 12112 16050
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11900 15422 12112 15450
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11612 15156 11664 15162
rect 11796 15156 11848 15162
rect 11664 15116 11744 15144
rect 11612 15098 11664 15104
rect 11610 13152 11666 13161
rect 11610 13087 11666 13096
rect 11624 12986 11652 13087
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11612 12708 11664 12714
rect 11612 12650 11664 12656
rect 11440 12406 11560 12434
rect 11440 11626 11468 12406
rect 11624 12322 11652 12650
rect 11532 12294 11652 12322
rect 11532 11762 11560 12294
rect 11612 12096 11664 12102
rect 11716 12084 11744 15116
rect 11796 15098 11848 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11808 12434 11836 14962
rect 11900 14958 11928 15302
rect 11992 15026 12020 15302
rect 12084 15201 12112 15422
rect 12070 15192 12126 15201
rect 12070 15127 12126 15136
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 12084 14618 12112 14962
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11888 13728 11940 13734
rect 12084 13716 12112 14350
rect 11940 13688 12112 13716
rect 11888 13670 11940 13676
rect 11900 13326 11928 13670
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12850 12020 13262
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12084 12730 12112 12786
rect 11992 12702 12112 12730
rect 11992 12646 12020 12702
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 12072 12640 12124 12646
rect 12072 12582 12124 12588
rect 11808 12406 12020 12434
rect 11992 12170 12020 12406
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11664 12056 11744 12084
rect 11612 12038 11664 12044
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11440 9994 11468 10542
rect 11428 9988 11480 9994
rect 11428 9930 11480 9936
rect 11440 9586 11468 9930
rect 11624 9926 11652 12038
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11624 8566 11652 9862
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11624 6322 11652 8502
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 6798 11744 7686
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11716 6118 11744 6734
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11428 5636 11480 5642
rect 11348 5596 11428 5624
rect 11428 5578 11480 5584
rect 11440 4593 11468 5578
rect 11426 4584 11482 4593
rect 11426 4519 11482 4528
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 11244 1420 11296 1426
rect 11244 1362 11296 1368
rect 11152 740 11204 746
rect 11152 682 11204 688
rect 11256 160 11284 1362
rect 11348 1290 11376 3334
rect 11440 3233 11468 4519
rect 11716 4146 11744 6054
rect 11704 4140 11756 4146
rect 11808 4128 11836 10746
rect 11900 10606 11928 11494
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11992 9994 12020 12106
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11992 8498 12020 9930
rect 12084 9586 12112 12582
rect 12176 12434 12204 17682
rect 12254 17640 12310 17649
rect 12254 17575 12310 17584
rect 12268 17202 12296 17575
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 16114 12296 16390
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12360 15586 12388 19343
rect 12452 17678 12480 19910
rect 12530 19887 12586 19896
rect 12808 19848 12860 19854
rect 12636 19808 12808 19836
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18222 12572 19110
rect 12636 18465 12664 19808
rect 12808 19790 12860 19796
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12728 19446 12756 19654
rect 12818 19612 13126 19621
rect 12818 19610 12824 19612
rect 12880 19610 12904 19612
rect 12960 19610 12984 19612
rect 13040 19610 13064 19612
rect 13120 19610 13126 19612
rect 12880 19558 12882 19610
rect 13062 19558 13064 19610
rect 12818 19556 12824 19558
rect 12880 19556 12904 19558
rect 12960 19556 12984 19558
rect 13040 19556 13064 19558
rect 13120 19556 13126 19558
rect 12818 19547 13126 19556
rect 12716 19440 12768 19446
rect 12716 19382 12768 19388
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12622 18456 12678 18465
rect 12622 18391 12678 18400
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12728 18306 12756 18906
rect 12818 18524 13126 18533
rect 12818 18522 12824 18524
rect 12880 18522 12904 18524
rect 12960 18522 12984 18524
rect 13040 18522 13064 18524
rect 13120 18522 13126 18524
rect 12880 18470 12882 18522
rect 13062 18470 13064 18522
rect 12818 18468 12824 18470
rect 12880 18468 12904 18470
rect 12960 18468 12984 18470
rect 13040 18468 13064 18470
rect 13120 18468 13126 18470
rect 12818 18459 13126 18468
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12530 18048 12586 18057
rect 12530 17983 12586 17992
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12544 17082 12572 17983
rect 12452 17054 12572 17082
rect 12452 15706 12480 17054
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16697 12572 16934
rect 12530 16688 12586 16697
rect 12530 16623 12586 16632
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12268 15558 12388 15586
rect 12268 13326 12296 15558
rect 12346 15464 12402 15473
rect 12346 15399 12402 15408
rect 12256 13320 12308 13326
rect 12256 13262 12308 13268
rect 12176 12406 12296 12434
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11898 12204 12106
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 9994 12204 11834
rect 12268 10810 12296 12406
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12084 8634 12112 9522
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12176 8498 12204 9930
rect 12360 9761 12388 15399
rect 12636 15162 12664 18294
rect 12728 18278 12940 18306
rect 12912 18222 12940 18278
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12728 16250 12756 17682
rect 13096 17678 13124 18090
rect 13188 18057 13216 20760
rect 13280 20505 13308 23462
rect 13372 22094 13400 35119
rect 13556 33998 13584 35226
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13542 32872 13598 32881
rect 13542 32807 13544 32816
rect 13596 32807 13598 32816
rect 13544 32778 13596 32784
rect 13648 31754 13676 43114
rect 13740 42752 13768 44463
rect 14016 43602 14044 44463
rect 14292 43602 14320 44463
rect 14016 43574 14136 43602
rect 14292 43574 14412 43602
rect 14004 43444 14056 43450
rect 14004 43386 14056 43392
rect 13820 42764 13872 42770
rect 13740 42724 13820 42752
rect 13820 42706 13872 42712
rect 14016 38654 14044 43386
rect 14108 42702 14136 43574
rect 14188 43104 14240 43110
rect 14188 43046 14240 43052
rect 14280 43104 14332 43110
rect 14280 43046 14332 43052
rect 14096 42696 14148 42702
rect 14096 42638 14148 42644
rect 14200 41414 14228 43046
rect 14292 42945 14320 43046
rect 14278 42936 14334 42945
rect 14278 42871 14334 42880
rect 14384 42702 14412 43574
rect 14568 43364 14596 44463
rect 14844 43382 14872 44463
rect 14740 43376 14792 43382
rect 14568 43336 14740 43364
rect 14740 43318 14792 43324
rect 14832 43376 14884 43382
rect 14832 43318 14884 43324
rect 14924 43172 14976 43178
rect 14924 43114 14976 43120
rect 14936 42945 14964 43114
rect 14922 42936 14978 42945
rect 14922 42871 14978 42880
rect 15120 42752 15148 44463
rect 15396 43296 15424 44463
rect 15476 43308 15528 43314
rect 15396 43268 15476 43296
rect 15672 43296 15700 44463
rect 15948 43382 15976 44463
rect 16028 43716 16080 43722
rect 16028 43658 16080 43664
rect 15936 43376 15988 43382
rect 15936 43318 15988 43324
rect 16040 43314 16068 43658
rect 16224 43364 16252 44463
rect 16396 43376 16448 43382
rect 16224 43336 16396 43364
rect 16396 43318 16448 43324
rect 15844 43308 15896 43314
rect 15672 43268 15844 43296
rect 15476 43250 15528 43256
rect 15844 43250 15896 43256
rect 16028 43308 16080 43314
rect 16028 43250 16080 43256
rect 15292 43104 15344 43110
rect 15290 43072 15292 43081
rect 15844 43104 15896 43110
rect 15344 43072 15346 43081
rect 15290 43007 15346 43016
rect 15672 43064 15844 43092
rect 15200 42764 15252 42770
rect 15120 42724 15200 42752
rect 15200 42706 15252 42712
rect 14372 42696 14424 42702
rect 14372 42638 14424 42644
rect 15474 42664 15530 42673
rect 14924 42628 14976 42634
rect 15474 42599 15530 42608
rect 14924 42570 14976 42576
rect 14556 42560 14608 42566
rect 14556 42502 14608 42508
rect 14832 42560 14884 42566
rect 14832 42502 14884 42508
rect 14200 41386 14504 41414
rect 14476 38758 14504 41386
rect 14464 38752 14516 38758
rect 14464 38694 14516 38700
rect 14016 38626 14136 38654
rect 13912 37664 13964 37670
rect 13912 37606 13964 37612
rect 13728 37324 13780 37330
rect 13728 37266 13780 37272
rect 13740 35068 13768 37266
rect 13820 35760 13872 35766
rect 13820 35702 13872 35708
rect 13832 35222 13860 35702
rect 13820 35216 13872 35222
rect 13820 35158 13872 35164
rect 13740 35040 13860 35068
rect 13728 34128 13780 34134
rect 13728 34070 13780 34076
rect 13740 33658 13768 34070
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13832 31906 13860 35040
rect 13924 34542 13952 37606
rect 13912 34536 13964 34542
rect 13912 34478 13964 34484
rect 13924 33998 13952 34478
rect 13912 33992 13964 33998
rect 13910 33960 13912 33969
rect 13964 33960 13966 33969
rect 13910 33895 13966 33904
rect 14004 33924 14056 33930
rect 14004 33866 14056 33872
rect 14016 33658 14044 33866
rect 14004 33652 14056 33658
rect 14004 33594 14056 33600
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13924 32026 13952 33458
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 14016 32026 14044 32710
rect 13912 32020 13964 32026
rect 13912 31962 13964 31968
rect 14004 32020 14056 32026
rect 14004 31962 14056 31968
rect 13832 31878 13952 31906
rect 13820 31816 13872 31822
rect 13820 31758 13872 31764
rect 13556 31726 13676 31754
rect 13452 29504 13504 29510
rect 13452 29446 13504 29452
rect 13464 26926 13492 29446
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13452 26036 13504 26042
rect 13452 25978 13504 25984
rect 13464 23866 13492 25978
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13556 23474 13584 31726
rect 13728 31272 13780 31278
rect 13648 31220 13728 31226
rect 13648 31214 13780 31220
rect 13648 31198 13768 31214
rect 13648 30938 13676 31198
rect 13728 31136 13780 31142
rect 13728 31078 13780 31084
rect 13636 30932 13688 30938
rect 13636 30874 13688 30880
rect 13740 29696 13768 31078
rect 13832 30666 13860 31758
rect 13924 31657 13952 31878
rect 13910 31648 13966 31657
rect 13910 31583 13966 31592
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 13924 30802 13952 31282
rect 14004 31136 14056 31142
rect 14004 31078 14056 31084
rect 14016 30938 14044 31078
rect 14004 30932 14056 30938
rect 14004 30874 14056 30880
rect 13912 30796 13964 30802
rect 13912 30738 13964 30744
rect 13820 30660 13872 30666
rect 13820 30602 13872 30608
rect 13912 30388 13964 30394
rect 13912 30330 13964 30336
rect 13924 30190 13952 30330
rect 14004 30320 14056 30326
rect 14004 30262 14056 30268
rect 13912 30184 13964 30190
rect 13912 30126 13964 30132
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13648 29668 13768 29696
rect 13648 27033 13676 29668
rect 13832 29594 13860 29990
rect 13924 29714 13952 30126
rect 13912 29708 13964 29714
rect 13912 29650 13964 29656
rect 13832 29566 13952 29594
rect 13820 29232 13872 29238
rect 13820 29174 13872 29180
rect 13832 29073 13860 29174
rect 13818 29064 13874 29073
rect 13818 28999 13874 29008
rect 13728 28960 13780 28966
rect 13728 28902 13780 28908
rect 13820 28960 13872 28966
rect 13820 28902 13872 28908
rect 13740 27878 13768 28902
rect 13832 28762 13860 28902
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13924 28558 13952 29566
rect 14016 29306 14044 30262
rect 14004 29300 14056 29306
rect 14004 29242 14056 29248
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 13728 27872 13780 27878
rect 13728 27814 13780 27820
rect 13634 27024 13690 27033
rect 13634 26959 13690 26968
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13648 23730 13676 26522
rect 13740 25838 13768 27814
rect 13832 27402 13860 27950
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13832 26994 13860 27338
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13924 26382 13952 28494
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 14016 28082 14044 28358
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 14108 27849 14136 38626
rect 14464 38004 14516 38010
rect 14464 37946 14516 37952
rect 14476 37777 14504 37946
rect 14462 37768 14518 37777
rect 14462 37703 14518 37712
rect 14278 36136 14334 36145
rect 14278 36071 14334 36080
rect 14188 35488 14240 35494
rect 14188 35430 14240 35436
rect 14200 35018 14228 35430
rect 14188 35012 14240 35018
rect 14188 34954 14240 34960
rect 14188 34740 14240 34746
rect 14188 34682 14240 34688
rect 14094 27840 14150 27849
rect 14094 27775 14150 27784
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 14094 25936 14150 25945
rect 14094 25871 14150 25880
rect 14108 25838 14136 25871
rect 13728 25832 13780 25838
rect 14004 25832 14056 25838
rect 13728 25774 13780 25780
rect 13924 25792 14004 25820
rect 13726 24712 13782 24721
rect 13726 24647 13782 24656
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13464 23446 13584 23474
rect 13464 22710 13492 23446
rect 13740 23338 13768 24647
rect 13924 24342 13952 25792
rect 14004 25774 14056 25780
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23730 13860 24006
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13818 23624 13874 23633
rect 13818 23559 13874 23568
rect 13556 23310 13768 23338
rect 13452 22704 13504 22710
rect 13452 22646 13504 22652
rect 13372 22066 13492 22094
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13372 21010 13400 21966
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13266 20496 13322 20505
rect 13372 20466 13400 20946
rect 13464 20806 13492 22066
rect 13556 21350 13584 23310
rect 13832 22778 13860 23559
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13648 21554 13676 22170
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13648 20874 13676 21490
rect 13636 20868 13688 20874
rect 13636 20810 13688 20816
rect 13452 20800 13504 20806
rect 13452 20742 13504 20748
rect 13266 20431 13322 20440
rect 13360 20460 13412 20466
rect 13280 20346 13308 20431
rect 13360 20402 13412 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13280 20318 13492 20346
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13280 19258 13308 19994
rect 13464 19334 13492 20318
rect 13556 20058 13584 20402
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13542 19816 13598 19825
rect 13542 19751 13598 19760
rect 13556 19446 13584 19751
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13464 19306 13584 19334
rect 13280 19230 13400 19258
rect 13174 18048 13230 18057
rect 13174 17983 13230 17992
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 12818 17436 13126 17445
rect 12818 17434 12824 17436
rect 12880 17434 12904 17436
rect 12960 17434 12984 17436
rect 13040 17434 13064 17436
rect 13120 17434 13126 17436
rect 12880 17382 12882 17434
rect 13062 17382 13064 17434
rect 12818 17380 12824 17382
rect 12880 17380 12904 17382
rect 12960 17380 12984 17382
rect 13040 17380 13064 17382
rect 13120 17380 13126 17382
rect 12818 17371 13126 17380
rect 13280 17338 13308 17614
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 12820 17202 12848 17274
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 13372 16946 13400 19230
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13280 16918 13400 16946
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 12818 16348 13126 16357
rect 12818 16346 12824 16348
rect 12880 16346 12904 16348
rect 12960 16346 12984 16348
rect 13040 16346 13064 16348
rect 13120 16346 13126 16348
rect 12880 16294 12882 16346
rect 13062 16294 13064 16346
rect 12818 16292 12824 16294
rect 12880 16292 12904 16294
rect 12960 16292 12984 16294
rect 13040 16292 13064 16294
rect 13120 16292 13126 16294
rect 12818 16283 13126 16292
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12818 15260 13126 15269
rect 12818 15258 12824 15260
rect 12880 15258 12904 15260
rect 12960 15258 12984 15260
rect 13040 15258 13064 15260
rect 13120 15258 13126 15260
rect 12880 15206 12882 15258
rect 13062 15206 13064 15258
rect 12818 15204 12824 15206
rect 12880 15204 12904 15206
rect 12960 15204 12984 15206
rect 13040 15204 13064 15206
rect 13120 15204 13126 15206
rect 12818 15195 13126 15204
rect 12624 15156 12676 15162
rect 12544 15116 12624 15144
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 11898 12480 14962
rect 12544 12764 12572 15116
rect 12624 15098 12676 15104
rect 12808 14952 12860 14958
rect 12636 14912 12808 14940
rect 12636 14414 12664 14912
rect 12808 14894 12860 14900
rect 13188 14464 13216 16458
rect 13280 15434 13308 16918
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13372 16046 13400 16730
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 13004 14436 13308 14464
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12900 14408 12952 14414
rect 13004 14396 13032 14436
rect 12952 14368 13032 14396
rect 12900 14350 12952 14356
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12818 14172 13126 14181
rect 12818 14170 12824 14172
rect 12880 14170 12904 14172
rect 12960 14170 12984 14172
rect 13040 14170 13064 14172
rect 13120 14170 13126 14172
rect 12880 14118 12882 14170
rect 13062 14118 13064 14170
rect 12818 14116 12824 14118
rect 12880 14116 12904 14118
rect 12960 14116 12984 14118
rect 13040 14116 13064 14118
rect 13120 14116 13126 14118
rect 12818 14107 13126 14116
rect 13188 13954 13216 14214
rect 13096 13926 13216 13954
rect 13096 13870 13124 13926
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13084 13864 13136 13870
rect 13176 13864 13228 13870
rect 13084 13806 13136 13812
rect 13174 13832 13176 13841
rect 13228 13832 13230 13841
rect 12636 12866 12664 13806
rect 13004 13172 13032 13806
rect 13174 13767 13230 13776
rect 13176 13184 13228 13190
rect 13004 13144 13176 13172
rect 13176 13126 13228 13132
rect 12818 13084 13126 13093
rect 12818 13082 12824 13084
rect 12880 13082 12904 13084
rect 12960 13082 12984 13084
rect 13040 13082 13064 13084
rect 13120 13082 13126 13084
rect 12880 13030 12882 13082
rect 13062 13030 13064 13082
rect 12818 13028 12824 13030
rect 12880 13028 12904 13030
rect 12960 13028 12984 13030
rect 13040 13028 13064 13030
rect 13120 13028 13126 13030
rect 12818 13019 13126 13028
rect 12636 12838 12848 12866
rect 12544 12736 12664 12764
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12544 11898 12572 12242
rect 12636 12102 12664 12736
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 12238 12756 12582
rect 12820 12238 12848 12838
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12636 10146 12664 12038
rect 12818 11996 13126 12005
rect 12818 11994 12824 11996
rect 12880 11994 12904 11996
rect 12960 11994 12984 11996
rect 13040 11994 13064 11996
rect 13120 11994 13126 11996
rect 12880 11942 12882 11994
rect 13062 11942 13064 11994
rect 12818 11940 12824 11942
rect 12880 11940 12904 11942
rect 12960 11940 12984 11942
rect 13040 11940 13064 11942
rect 13120 11940 13126 11942
rect 12818 11931 13126 11940
rect 13188 11762 13216 12038
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12820 11642 12848 11698
rect 12820 11614 13032 11642
rect 13004 11558 13032 11614
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13188 11150 13216 11698
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 12544 10118 12664 10146
rect 12544 9926 12572 10118
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12346 9752 12402 9761
rect 12346 9687 12402 9696
rect 12348 9648 12400 9654
rect 12268 9608 12348 9636
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 11978 8392 12034 8401
rect 11978 8327 12034 8336
rect 11808 4100 11928 4128
rect 11704 4082 11756 4088
rect 11518 4040 11574 4049
rect 11518 3975 11574 3984
rect 11532 3534 11560 3975
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11426 3224 11482 3233
rect 11426 3159 11482 3168
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11532 1465 11560 2382
rect 11624 2038 11652 3334
rect 11716 2972 11744 4082
rect 11794 4040 11850 4049
rect 11794 3975 11850 3984
rect 11808 3534 11836 3975
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11900 3074 11928 4100
rect 11992 3194 12020 8327
rect 12084 8090 12112 8434
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12268 7886 12296 9608
rect 12348 9590 12400 9596
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12452 8838 12480 8910
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8634 12480 8774
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12544 8498 12572 9862
rect 12636 9722 12664 9998
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12072 7744 12124 7750
rect 12360 7732 12388 8434
rect 12072 7686 12124 7692
rect 12268 7704 12388 7732
rect 12084 3738 12112 7686
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12176 5914 12204 6122
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 4690 12204 5714
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11900 3058 12112 3074
rect 11900 3052 12124 3058
rect 11900 3046 12072 3052
rect 11796 2984 11848 2990
rect 11716 2944 11796 2972
rect 11900 2961 11928 3046
rect 12072 2994 12124 3000
rect 11980 2984 12032 2990
rect 11796 2926 11848 2932
rect 11886 2952 11942 2961
rect 11980 2926 12032 2932
rect 11886 2887 11942 2896
rect 11888 2848 11940 2854
rect 11808 2796 11888 2802
rect 11808 2790 11940 2796
rect 11808 2774 11928 2790
rect 11808 2446 11836 2774
rect 11992 2514 12020 2926
rect 12070 2680 12126 2689
rect 12070 2615 12126 2624
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 12084 2446 12112 2615
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 2106 11928 2246
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11888 1760 11940 1766
rect 11808 1720 11888 1748
rect 11518 1456 11574 1465
rect 11518 1391 11574 1400
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 11336 1284 11388 1290
rect 11336 1226 11388 1232
rect 11716 1018 11744 1294
rect 11704 1012 11756 1018
rect 11704 954 11756 960
rect 11520 944 11572 950
rect 11520 886 11572 892
rect 11532 160 11560 886
rect 11808 160 11836 1720
rect 11888 1702 11940 1708
rect 12176 1290 12204 2518
rect 12164 1284 12216 1290
rect 12164 1226 12216 1232
rect 11888 1216 11940 1222
rect 12072 1216 12124 1222
rect 11940 1164 12072 1170
rect 11888 1158 12124 1164
rect 11900 1142 12112 1158
rect 12072 876 12124 882
rect 12072 818 12124 824
rect 12084 160 12112 818
rect 12268 542 12296 7704
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12452 6265 12480 7278
rect 12544 6458 12572 8434
rect 12636 7954 12664 9318
rect 12728 8566 12756 11086
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 12818 10908 13126 10917
rect 12818 10906 12824 10908
rect 12880 10906 12904 10908
rect 12960 10906 12984 10908
rect 13040 10906 13064 10908
rect 13120 10906 13126 10908
rect 12880 10854 12882 10906
rect 13062 10854 13064 10906
rect 12818 10852 12824 10854
rect 12880 10852 12904 10854
rect 12960 10852 12984 10854
rect 13040 10852 13064 10854
rect 13120 10852 13126 10854
rect 12818 10843 13126 10852
rect 13188 10742 13216 10950
rect 13280 10810 13308 14436
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 12818 9820 13126 9829
rect 12818 9818 12824 9820
rect 12880 9818 12904 9820
rect 12960 9818 12984 9820
rect 13040 9818 13064 9820
rect 13120 9818 13126 9820
rect 12880 9766 12882 9818
rect 13062 9766 13064 9818
rect 12818 9764 12824 9766
rect 12880 9764 12904 9766
rect 12960 9764 12984 9766
rect 13040 9764 13064 9766
rect 13120 9764 13126 9766
rect 12818 9755 13126 9764
rect 12818 8732 13126 8741
rect 12818 8730 12824 8732
rect 12880 8730 12904 8732
rect 12960 8730 12984 8732
rect 13040 8730 13064 8732
rect 13120 8730 13126 8732
rect 12880 8678 12882 8730
rect 13062 8678 13064 8730
rect 12818 8676 12824 8678
rect 12880 8676 12904 8678
rect 12960 8676 12984 8678
rect 13040 8676 13064 8678
rect 13120 8676 13126 8678
rect 12818 8667 13126 8676
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12440 6259 12492 6265
rect 12440 6201 12492 6207
rect 12452 5914 12480 6201
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12452 5778 12480 5850
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12636 5234 12664 7414
rect 12728 6440 12756 8502
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 7886 13032 8230
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12818 7644 13126 7653
rect 12818 7642 12824 7644
rect 12880 7642 12904 7644
rect 12960 7642 12984 7644
rect 13040 7642 13064 7644
rect 13120 7642 13126 7644
rect 12880 7590 12882 7642
rect 13062 7590 13064 7642
rect 12818 7588 12824 7590
rect 12880 7588 12904 7590
rect 12960 7588 12984 7590
rect 13040 7588 13064 7590
rect 13120 7588 13126 7590
rect 12818 7579 13126 7588
rect 13188 6662 13216 10406
rect 13266 10024 13322 10033
rect 13266 9959 13322 9968
rect 13280 9722 13308 9959
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13280 8294 13308 8842
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13372 7818 13400 15982
rect 13464 15162 13492 17138
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14550 13492 14962
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13556 14090 13584 19306
rect 13648 16590 13676 20810
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 14618 13676 16050
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13464 14062 13584 14090
rect 13464 13841 13492 14062
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13544 13864 13596 13870
rect 13450 13832 13506 13841
rect 13544 13806 13596 13812
rect 13450 13767 13506 13776
rect 13556 13682 13584 13806
rect 13464 13654 13584 13682
rect 13464 13530 13492 13654
rect 13542 13560 13598 13569
rect 13452 13524 13504 13530
rect 13648 13530 13676 13874
rect 13542 13495 13598 13504
rect 13636 13524 13688 13530
rect 13452 13466 13504 13472
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13464 8566 13492 10678
rect 13556 8974 13584 13495
rect 13636 13466 13688 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 10470 13676 13330
rect 13740 12102 13768 18022
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13726 11928 13782 11937
rect 13726 11863 13782 11872
rect 13740 11694 13768 11863
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13832 11354 13860 20742
rect 13924 20398 13952 24278
rect 14004 23656 14056 23662
rect 14108 23644 14136 25774
rect 14056 23616 14136 23644
rect 14004 23598 14056 23604
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13912 19440 13964 19446
rect 13910 19408 13912 19417
rect 13964 19408 13966 19417
rect 13910 19343 13966 19352
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13924 15978 13952 17614
rect 14016 16522 14044 23462
rect 14200 22094 14228 34682
rect 14292 33862 14320 36071
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14292 31822 14320 33798
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14384 30394 14412 33458
rect 14476 32502 14504 34886
rect 14568 34649 14596 42502
rect 14740 42288 14792 42294
rect 14740 42230 14792 42236
rect 14648 41268 14700 41274
rect 14648 41210 14700 41216
rect 14554 34640 14610 34649
rect 14554 34575 14610 34584
rect 14464 32496 14516 32502
rect 14464 32438 14516 32444
rect 14660 31754 14688 41210
rect 14568 31726 14688 31754
rect 14372 30388 14424 30394
rect 14372 30330 14424 30336
rect 14568 29646 14596 31726
rect 14648 29844 14700 29850
rect 14648 29786 14700 29792
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14464 29504 14516 29510
rect 14464 29446 14516 29452
rect 14476 29306 14504 29446
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 14556 29232 14608 29238
rect 14660 29220 14688 29786
rect 14608 29192 14688 29220
rect 14556 29174 14608 29180
rect 14280 28960 14332 28966
rect 14332 28908 14412 28914
rect 14280 28902 14412 28908
rect 14292 28886 14412 28902
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 14292 25906 14320 28358
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14384 25786 14412 28886
rect 14462 27840 14518 27849
rect 14462 27775 14518 27784
rect 14292 25758 14412 25786
rect 14292 23526 14320 25758
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14292 22681 14320 23054
rect 14278 22672 14334 22681
rect 14278 22607 14334 22616
rect 14108 22066 14228 22094
rect 14108 20806 14136 22066
rect 14280 21548 14332 21554
rect 14280 21490 14332 21496
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14292 20466 14320 21490
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14108 18290 14136 19654
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14094 17232 14150 17241
rect 14094 17167 14150 17176
rect 14108 17134 14136 17167
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14094 16688 14150 16697
rect 14200 16674 14228 20334
rect 14292 20058 14320 20402
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14292 19514 14320 19790
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14292 18698 14320 19450
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14384 17338 14412 24006
rect 14476 23497 14504 27775
rect 14462 23488 14518 23497
rect 14462 23423 14518 23432
rect 14568 22982 14596 29174
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14660 27470 14688 27814
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14648 27328 14700 27334
rect 14648 27270 14700 27276
rect 14660 26926 14688 27270
rect 14648 26920 14700 26926
rect 14648 26862 14700 26868
rect 14752 26466 14780 42230
rect 14844 34610 14872 42502
rect 14832 34604 14884 34610
rect 14832 34546 14884 34552
rect 14832 32428 14884 32434
rect 14832 32370 14884 32376
rect 14844 31754 14872 32370
rect 14832 31748 14884 31754
rect 14832 31690 14884 31696
rect 14844 30870 14872 31690
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14844 30326 14872 30806
rect 14832 30320 14884 30326
rect 14936 30297 14964 42570
rect 15488 42566 15516 42599
rect 15476 42560 15528 42566
rect 15476 42502 15528 42508
rect 15568 42560 15620 42566
rect 15568 42502 15620 42508
rect 15384 42084 15436 42090
rect 15384 42026 15436 42032
rect 15108 41268 15160 41274
rect 15108 41210 15160 41216
rect 15120 40633 15148 41210
rect 15106 40624 15162 40633
rect 15106 40559 15162 40568
rect 15396 34746 15424 42026
rect 15476 37868 15528 37874
rect 15476 37810 15528 37816
rect 15488 35494 15516 37810
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15488 35154 15516 35430
rect 15476 35148 15528 35154
rect 15476 35090 15528 35096
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15384 34740 15436 34746
rect 15384 34682 15436 34688
rect 15016 34604 15068 34610
rect 15016 34546 15068 34552
rect 15028 34513 15056 34546
rect 15014 34504 15070 34513
rect 15014 34439 15070 34448
rect 15016 34400 15068 34406
rect 15016 34342 15068 34348
rect 15028 33862 15056 34342
rect 15200 34060 15252 34066
rect 15200 34002 15252 34008
rect 15016 33856 15068 33862
rect 15016 33798 15068 33804
rect 15108 33856 15160 33862
rect 15108 33798 15160 33804
rect 15120 33114 15148 33798
rect 15212 33522 15240 34002
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15304 32910 15332 34682
rect 15488 34066 15516 35090
rect 15476 34060 15528 34066
rect 15476 34002 15528 34008
rect 15384 33992 15436 33998
rect 15384 33934 15436 33940
rect 15396 33114 15424 33934
rect 15384 33108 15436 33114
rect 15384 33050 15436 33056
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 15108 32904 15160 32910
rect 15108 32846 15160 32852
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15382 32872 15438 32881
rect 15028 32570 15056 32846
rect 15016 32564 15068 32570
rect 15016 32506 15068 32512
rect 15028 30326 15056 32506
rect 15120 32502 15148 32846
rect 15382 32807 15438 32816
rect 15396 32774 15424 32807
rect 15292 32768 15344 32774
rect 15292 32710 15344 32716
rect 15384 32768 15436 32774
rect 15384 32710 15436 32716
rect 15304 32570 15332 32710
rect 15292 32564 15344 32570
rect 15292 32506 15344 32512
rect 15108 32496 15160 32502
rect 15108 32438 15160 32444
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15200 32360 15252 32366
rect 15200 32302 15252 32308
rect 15120 32026 15148 32302
rect 15108 32020 15160 32026
rect 15108 31962 15160 31968
rect 15212 31822 15240 32302
rect 15304 32026 15332 32506
rect 15292 32020 15344 32026
rect 15292 31962 15344 31968
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15290 31648 15346 31657
rect 15290 31583 15346 31592
rect 15016 30320 15068 30326
rect 14832 30262 14884 30268
rect 14922 30288 14978 30297
rect 15016 30262 15068 30268
rect 14922 30223 14978 30232
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14844 29306 14872 29990
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 14660 26438 14780 26466
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14476 19990 14504 22714
rect 14568 22409 14596 22918
rect 14554 22400 14610 22409
rect 14554 22335 14610 22344
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14464 19984 14516 19990
rect 14464 19926 14516 19932
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18834 14504 19110
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14568 18086 14596 20402
rect 14660 19334 14688 26438
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 14752 22778 14780 26318
rect 14844 24274 14872 29242
rect 14936 29102 14964 29990
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 15106 28656 15162 28665
rect 15106 28591 15162 28600
rect 15120 28558 15148 28591
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 14924 28076 14976 28082
rect 14924 28018 14976 28024
rect 14936 27713 14964 28018
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 14922 27704 14978 27713
rect 14922 27639 14978 27648
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 14832 23792 14884 23798
rect 14832 23734 14884 23740
rect 14844 23322 14872 23734
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22098 14872 22374
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14752 21690 14780 22034
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14936 21026 14964 27639
rect 15120 27538 15148 27950
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 15028 26042 15056 27270
rect 15212 27130 15240 28494
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 15108 26988 15160 26994
rect 15108 26930 15160 26936
rect 15120 26897 15148 26930
rect 15106 26888 15162 26897
rect 15162 26846 15240 26874
rect 15106 26823 15162 26832
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15016 24948 15068 24954
rect 15016 24890 15068 24896
rect 15028 24410 15056 24890
rect 15106 24576 15162 24585
rect 15106 24511 15162 24520
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15028 21554 15056 23258
rect 15120 23118 15148 24511
rect 15212 24177 15240 26846
rect 15304 25106 15332 31583
rect 15382 31240 15438 31249
rect 15382 31175 15438 31184
rect 15396 25362 15424 31175
rect 15488 30802 15516 31758
rect 15580 31482 15608 42502
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 15476 30796 15528 30802
rect 15476 30738 15528 30744
rect 15568 30728 15620 30734
rect 15568 30670 15620 30676
rect 15474 29200 15530 29209
rect 15474 29135 15476 29144
rect 15528 29135 15530 29144
rect 15476 29106 15528 29112
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15304 25078 15424 25106
rect 15290 24984 15346 24993
rect 15290 24919 15346 24928
rect 15198 24168 15254 24177
rect 15198 24103 15254 24112
rect 15304 23882 15332 24919
rect 15396 24721 15424 25078
rect 15382 24712 15438 24721
rect 15382 24647 15438 24656
rect 15488 24070 15516 29106
rect 15580 28558 15608 30670
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15672 26466 15700 43064
rect 15844 43046 15896 43052
rect 15785 43004 16093 43013
rect 15785 43002 15791 43004
rect 15847 43002 15871 43004
rect 15927 43002 15951 43004
rect 16007 43002 16031 43004
rect 16087 43002 16093 43004
rect 15847 42950 15849 43002
rect 16029 42950 16031 43002
rect 15785 42948 15791 42950
rect 15847 42948 15871 42950
rect 15927 42948 15951 42950
rect 16007 42948 16031 42950
rect 16087 42948 16093 42950
rect 15785 42939 16093 42948
rect 16500 42786 16528 44463
rect 16776 43364 16804 44463
rect 17052 43450 17080 44463
rect 17040 43444 17092 43450
rect 17040 43386 17092 43392
rect 16856 43376 16908 43382
rect 16776 43336 16856 43364
rect 16856 43318 16908 43324
rect 17328 43246 17356 44463
rect 17500 43648 17552 43654
rect 17500 43590 17552 43596
rect 17408 43308 17460 43314
rect 17408 43250 17460 43256
rect 17316 43240 17368 43246
rect 17316 43182 17368 43188
rect 16856 43104 16908 43110
rect 16856 43046 16908 43052
rect 16868 42906 16896 43046
rect 16856 42900 16908 42906
rect 16856 42842 16908 42848
rect 16500 42758 16620 42786
rect 16592 42702 16620 42758
rect 16488 42696 16540 42702
rect 16488 42638 16540 42644
rect 16580 42696 16632 42702
rect 16580 42638 16632 42644
rect 16120 42628 16172 42634
rect 16120 42570 16172 42576
rect 15785 41916 16093 41925
rect 15785 41914 15791 41916
rect 15847 41914 15871 41916
rect 15927 41914 15951 41916
rect 16007 41914 16031 41916
rect 16087 41914 16093 41916
rect 15847 41862 15849 41914
rect 16029 41862 16031 41914
rect 15785 41860 15791 41862
rect 15847 41860 15871 41862
rect 15927 41860 15951 41862
rect 16007 41860 16031 41862
rect 16087 41860 16093 41862
rect 15785 41851 16093 41860
rect 15785 40828 16093 40837
rect 15785 40826 15791 40828
rect 15847 40826 15871 40828
rect 15927 40826 15951 40828
rect 16007 40826 16031 40828
rect 16087 40826 16093 40828
rect 15847 40774 15849 40826
rect 16029 40774 16031 40826
rect 15785 40772 15791 40774
rect 15847 40772 15871 40774
rect 15927 40772 15951 40774
rect 16007 40772 16031 40774
rect 16087 40772 16093 40774
rect 15785 40763 16093 40772
rect 15785 39740 16093 39749
rect 15785 39738 15791 39740
rect 15847 39738 15871 39740
rect 15927 39738 15951 39740
rect 16007 39738 16031 39740
rect 16087 39738 16093 39740
rect 15847 39686 15849 39738
rect 16029 39686 16031 39738
rect 15785 39684 15791 39686
rect 15847 39684 15871 39686
rect 15927 39684 15951 39686
rect 16007 39684 16031 39686
rect 16087 39684 16093 39686
rect 15785 39675 16093 39684
rect 15785 38652 16093 38661
rect 15785 38650 15791 38652
rect 15847 38650 15871 38652
rect 15927 38650 15951 38652
rect 16007 38650 16031 38652
rect 16087 38650 16093 38652
rect 15847 38598 15849 38650
rect 16029 38598 16031 38650
rect 15785 38596 15791 38598
rect 15847 38596 15871 38598
rect 15927 38596 15951 38598
rect 16007 38596 16031 38598
rect 16087 38596 16093 38598
rect 15785 38587 16093 38596
rect 15785 37564 16093 37573
rect 15785 37562 15791 37564
rect 15847 37562 15871 37564
rect 15927 37562 15951 37564
rect 16007 37562 16031 37564
rect 16087 37562 16093 37564
rect 15847 37510 15849 37562
rect 16029 37510 16031 37562
rect 15785 37508 15791 37510
rect 15847 37508 15871 37510
rect 15927 37508 15951 37510
rect 16007 37508 16031 37510
rect 16087 37508 16093 37510
rect 15785 37499 16093 37508
rect 15785 36476 16093 36485
rect 15785 36474 15791 36476
rect 15847 36474 15871 36476
rect 15927 36474 15951 36476
rect 16007 36474 16031 36476
rect 16087 36474 16093 36476
rect 15847 36422 15849 36474
rect 16029 36422 16031 36474
rect 15785 36420 15791 36422
rect 15847 36420 15871 36422
rect 15927 36420 15951 36422
rect 16007 36420 16031 36422
rect 16087 36420 16093 36422
rect 15785 36411 16093 36420
rect 15785 35388 16093 35397
rect 15785 35386 15791 35388
rect 15847 35386 15871 35388
rect 15927 35386 15951 35388
rect 16007 35386 16031 35388
rect 16087 35386 16093 35388
rect 15847 35334 15849 35386
rect 16029 35334 16031 35386
rect 15785 35332 15791 35334
rect 15847 35332 15871 35334
rect 15927 35332 15951 35334
rect 16007 35332 16031 35334
rect 16087 35332 16093 35334
rect 15785 35323 16093 35332
rect 15785 34300 16093 34309
rect 15785 34298 15791 34300
rect 15847 34298 15871 34300
rect 15927 34298 15951 34300
rect 16007 34298 16031 34300
rect 16087 34298 16093 34300
rect 15847 34246 15849 34298
rect 16029 34246 16031 34298
rect 15785 34244 15791 34246
rect 15847 34244 15871 34246
rect 15927 34244 15951 34246
rect 16007 34244 16031 34246
rect 16087 34244 16093 34246
rect 15785 34235 16093 34244
rect 15785 33212 16093 33221
rect 15785 33210 15791 33212
rect 15847 33210 15871 33212
rect 15927 33210 15951 33212
rect 16007 33210 16031 33212
rect 16087 33210 16093 33212
rect 15847 33158 15849 33210
rect 16029 33158 16031 33210
rect 15785 33156 15791 33158
rect 15847 33156 15871 33158
rect 15927 33156 15951 33158
rect 16007 33156 16031 33158
rect 16087 33156 16093 33158
rect 15785 33147 16093 33156
rect 16132 33114 16160 42570
rect 16396 42560 16448 42566
rect 16396 42502 16448 42508
rect 16408 42294 16436 42502
rect 16396 42288 16448 42294
rect 16396 42230 16448 42236
rect 16500 42090 16528 42638
rect 16948 42560 17000 42566
rect 16948 42502 17000 42508
rect 17224 42560 17276 42566
rect 17224 42502 17276 42508
rect 17316 42560 17368 42566
rect 17316 42502 17368 42508
rect 16960 42294 16988 42502
rect 17236 42362 17264 42502
rect 17328 42362 17356 42502
rect 17224 42356 17276 42362
rect 17224 42298 17276 42304
rect 17316 42356 17368 42362
rect 17316 42298 17368 42304
rect 16948 42288 17000 42294
rect 16948 42230 17000 42236
rect 17040 42220 17092 42226
rect 17040 42162 17092 42168
rect 16488 42084 16540 42090
rect 16488 42026 16540 42032
rect 16948 42084 17000 42090
rect 16948 42026 17000 42032
rect 16304 42016 16356 42022
rect 16304 41958 16356 41964
rect 16212 34196 16264 34202
rect 16212 34138 16264 34144
rect 16224 33998 16252 34138
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16120 33108 16172 33114
rect 16120 33050 16172 33056
rect 15785 32124 16093 32133
rect 15785 32122 15791 32124
rect 15847 32122 15871 32124
rect 15927 32122 15951 32124
rect 16007 32122 16031 32124
rect 16087 32122 16093 32124
rect 15847 32070 15849 32122
rect 16029 32070 16031 32122
rect 15785 32068 15791 32070
rect 15847 32068 15871 32070
rect 15927 32068 15951 32070
rect 16007 32068 16031 32070
rect 16087 32068 16093 32070
rect 15785 32059 16093 32068
rect 15752 32020 15804 32026
rect 15752 31962 15804 31968
rect 15764 31822 15792 31962
rect 16224 31958 16252 33254
rect 16212 31952 16264 31958
rect 16212 31894 16264 31900
rect 15752 31816 15804 31822
rect 15804 31776 15884 31804
rect 15752 31758 15804 31764
rect 15752 31680 15804 31686
rect 15752 31622 15804 31628
rect 15764 31346 15792 31622
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15750 31240 15806 31249
rect 15856 31226 15884 31776
rect 16026 31784 16082 31793
rect 16026 31719 16082 31728
rect 16040 31686 16068 31719
rect 16028 31680 16080 31686
rect 16028 31622 16080 31628
rect 15806 31198 15884 31226
rect 15750 31175 15806 31184
rect 16120 31136 16172 31142
rect 16120 31078 16172 31084
rect 15785 31036 16093 31045
rect 15785 31034 15791 31036
rect 15847 31034 15871 31036
rect 15927 31034 15951 31036
rect 16007 31034 16031 31036
rect 16087 31034 16093 31036
rect 15847 30982 15849 31034
rect 16029 30982 16031 31034
rect 15785 30980 15791 30982
rect 15847 30980 15871 30982
rect 15927 30980 15951 30982
rect 16007 30980 16031 30982
rect 16087 30980 16093 30982
rect 15785 30971 16093 30980
rect 16132 30938 16160 31078
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 15785 29948 16093 29957
rect 15785 29946 15791 29948
rect 15847 29946 15871 29948
rect 15927 29946 15951 29948
rect 16007 29946 16031 29948
rect 16087 29946 16093 29948
rect 15847 29894 15849 29946
rect 16029 29894 16031 29946
rect 15785 29892 15791 29894
rect 15847 29892 15871 29894
rect 15927 29892 15951 29894
rect 16007 29892 16031 29894
rect 16087 29892 16093 29894
rect 15785 29883 16093 29892
rect 15752 29708 15804 29714
rect 15804 29668 15884 29696
rect 15752 29650 15804 29656
rect 15856 29345 15884 29668
rect 15936 29640 15988 29646
rect 15936 29582 15988 29588
rect 15948 29510 15976 29582
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15842 29336 15898 29345
rect 15842 29271 15898 29280
rect 15785 28860 16093 28869
rect 15785 28858 15791 28860
rect 15847 28858 15871 28860
rect 15927 28858 15951 28860
rect 16007 28858 16031 28860
rect 16087 28858 16093 28860
rect 15847 28806 15849 28858
rect 16029 28806 16031 28858
rect 15785 28804 15791 28806
rect 15847 28804 15871 28806
rect 15927 28804 15951 28806
rect 16007 28804 16031 28806
rect 16087 28804 16093 28806
rect 15785 28795 16093 28804
rect 16132 28558 16160 30670
rect 16224 29782 16252 31894
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 16212 28960 16264 28966
rect 16212 28902 16264 28908
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 15785 27772 16093 27781
rect 15785 27770 15791 27772
rect 15847 27770 15871 27772
rect 15927 27770 15951 27772
rect 16007 27770 16031 27772
rect 16087 27770 16093 27772
rect 15847 27718 15849 27770
rect 16029 27718 16031 27770
rect 15785 27716 15791 27718
rect 15847 27716 15871 27718
rect 15927 27716 15951 27718
rect 16007 27716 16031 27718
rect 16087 27716 16093 27718
rect 15785 27707 16093 27716
rect 15785 26684 16093 26693
rect 15785 26682 15791 26684
rect 15847 26682 15871 26684
rect 15927 26682 15951 26684
rect 16007 26682 16031 26684
rect 16087 26682 16093 26684
rect 15847 26630 15849 26682
rect 16029 26630 16031 26682
rect 15785 26628 15791 26630
rect 15847 26628 15871 26630
rect 15927 26628 15951 26630
rect 16007 26628 16031 26630
rect 16087 26628 16093 26630
rect 15785 26619 16093 26628
rect 15844 26580 15896 26586
rect 16028 26580 16080 26586
rect 15896 26540 16028 26568
rect 15844 26522 15896 26528
rect 16028 26522 16080 26528
rect 15580 26438 15700 26466
rect 15936 26444 15988 26450
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15304 23854 15516 23882
rect 15108 23112 15160 23118
rect 15108 23054 15160 23060
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15120 22094 15148 22918
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15292 22094 15344 22098
rect 15120 22092 15344 22094
rect 15120 22066 15292 22092
rect 15292 22034 15344 22040
rect 15108 22024 15160 22030
rect 15304 22003 15332 22034
rect 15108 21966 15160 21972
rect 15120 21604 15148 21966
rect 15396 21894 15424 22714
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15488 21672 15516 23854
rect 15396 21644 15516 21672
rect 15200 21616 15252 21622
rect 15120 21576 15200 21604
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15028 21078 15056 21286
rect 14752 20998 14964 21026
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 14752 20466 14780 20998
rect 14832 20936 14884 20942
rect 15120 20924 15148 21576
rect 15200 21558 15252 21564
rect 15396 21554 15424 21644
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15396 21162 15424 21490
rect 14832 20878 14884 20884
rect 14936 20896 15148 20924
rect 15304 21134 15424 21162
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14844 20262 14872 20878
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14660 19306 14780 19334
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14660 18426 14688 18634
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14554 17232 14610 17241
rect 14610 17190 14688 17218
rect 14554 17167 14610 17176
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14150 16646 14228 16674
rect 14094 16623 14150 16632
rect 14476 16590 14504 16934
rect 14464 16584 14516 16590
rect 14660 16574 14688 17190
rect 14464 16526 14516 16532
rect 14568 16546 14688 16574
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 14016 16402 14044 16458
rect 14016 16374 14228 16402
rect 14094 16144 14150 16153
rect 14094 16079 14150 16088
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13924 13394 13952 15914
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 14016 13870 14044 14758
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13924 11898 13952 12242
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13924 11234 13952 11494
rect 13740 11206 13952 11234
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13634 9888 13690 9897
rect 13634 9823 13690 9832
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 13464 7478 13492 8502
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 12728 6412 12848 6440
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12728 5846 12756 6258
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12820 5556 12848 6412
rect 12728 5528 12848 5556
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12728 4842 12756 5528
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 5001 13124 5102
rect 13082 4992 13138 5001
rect 13082 4927 13138 4936
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12728 4814 12848 4842
rect 12360 4282 12388 4762
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12728 4214 12756 4814
rect 12820 4622 12848 4814
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 13188 4282 13216 6598
rect 13280 6458 13308 7142
rect 13464 7002 13492 7278
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13358 6216 13414 6225
rect 13358 6151 13360 6160
rect 13412 6151 13414 6160
rect 13360 6122 13412 6128
rect 13450 6080 13506 6089
rect 13280 6038 13450 6066
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 12716 4208 12768 4214
rect 13188 4185 13216 4218
rect 12716 4150 12768 4156
rect 13174 4176 13230 4185
rect 13174 4111 13230 4120
rect 12532 3936 12584 3942
rect 12346 3904 12402 3913
rect 12532 3878 12584 3884
rect 12346 3839 12402 3848
rect 12360 3466 12388 3839
rect 12544 3602 12572 3878
rect 12898 3768 12954 3777
rect 12898 3703 12954 3712
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12912 3466 12940 3703
rect 13280 3618 13308 6038
rect 13450 6015 13506 6024
rect 13556 5930 13584 8570
rect 13464 5902 13584 5930
rect 13464 5273 13492 5902
rect 13648 5386 13676 9823
rect 13740 8634 13768 11206
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13818 9752 13874 9761
rect 13818 9687 13874 9696
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8514 13860 9687
rect 13740 8486 13860 8514
rect 13924 8498 13952 10678
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14016 10266 14044 10610
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9722 14044 9998
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 14016 9382 14044 9658
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9042 14044 9318
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13912 8492 13964 8498
rect 13740 7750 13768 8486
rect 13912 8434 13964 8440
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13832 8090 13860 8366
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13924 7970 13952 8434
rect 13832 7942 13952 7970
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13832 7478 13860 7942
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13924 6458 13952 7346
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13726 6352 13782 6361
rect 13726 6287 13728 6296
rect 13780 6287 13782 6296
rect 13728 6258 13780 6264
rect 13726 5536 13782 5545
rect 13726 5471 13782 5480
rect 13556 5358 13676 5386
rect 13450 5264 13506 5273
rect 13450 5199 13506 5208
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13372 4826 13400 5034
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13556 3720 13584 5358
rect 13556 3692 13676 3720
rect 13176 3596 13228 3602
rect 13280 3590 13584 3618
rect 13176 3538 13228 3544
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 12452 3194 12480 3402
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 2378 12572 3402
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12348 1420 12400 1426
rect 12348 1362 12400 1368
rect 12256 536 12308 542
rect 12256 478 12308 484
rect 12360 160 12388 1362
rect 12452 814 12480 2246
rect 12636 1970 12664 3062
rect 13188 2774 13216 3538
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13188 2746 13400 2774
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13280 2446 13308 2586
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12440 808 12492 814
rect 12440 750 12492 756
rect 12636 160 12664 1702
rect 13188 1562 13216 2246
rect 13176 1556 13228 1562
rect 13176 1498 13228 1504
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 12728 660 12756 1294
rect 13084 1216 13136 1222
rect 13136 1176 13216 1204
rect 13084 1158 13136 1164
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12728 632 12940 660
rect 12912 160 12940 632
rect 13188 160 13216 1176
rect 13372 1018 13400 2746
rect 13464 1408 13492 2790
rect 13556 2650 13584 3590
rect 13648 3534 13676 3692
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13740 3346 13768 5471
rect 13818 5264 13874 5273
rect 13818 5199 13874 5208
rect 13912 5228 13964 5234
rect 13832 5166 13860 5199
rect 13912 5170 13964 5176
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13924 3738 13952 5170
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13648 3318 13768 3346
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13544 2440 13596 2446
rect 13542 2408 13544 2417
rect 13596 2408 13598 2417
rect 13542 2343 13598 2352
rect 13648 2106 13676 3318
rect 13818 2680 13874 2689
rect 13818 2615 13874 2624
rect 13832 2446 13860 2615
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 13832 1873 13860 1906
rect 13818 1864 13874 1873
rect 13818 1799 13874 1808
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 13544 1420 13596 1426
rect 13464 1380 13544 1408
rect 13544 1362 13596 1368
rect 13648 1358 13676 1702
rect 13820 1556 13872 1562
rect 13820 1498 13872 1504
rect 13832 1408 13860 1498
rect 13740 1380 13860 1408
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13360 1012 13412 1018
rect 13360 954 13412 960
rect 13464 160 13492 1158
rect 13740 160 13768 1380
rect 13924 1358 13952 2518
rect 14016 2446 14044 7346
rect 14108 4826 14136 16079
rect 14200 12434 14228 16374
rect 14280 16108 14332 16114
rect 14332 16068 14412 16096
rect 14280 16050 14332 16056
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14292 15366 14320 15846
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 14414 14320 15302
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 14278 13968 14334 13977
rect 14278 13903 14280 13912
rect 14332 13903 14334 13912
rect 14280 13874 14332 13880
rect 14384 13326 14412 16068
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14476 14006 14504 15370
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14384 12434 14412 13262
rect 14200 12406 14320 12434
rect 14384 12406 14504 12434
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14200 10742 14228 12106
rect 14292 12102 14320 12406
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14384 12102 14412 12174
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14292 10810 14320 12038
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14372 9988 14424 9994
rect 14476 9976 14504 12406
rect 14424 9948 14504 9976
rect 14372 9930 14424 9936
rect 14568 9674 14596 16546
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14660 14618 14688 14826
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14660 13326 14688 14554
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14752 13190 14780 19306
rect 14936 18766 14964 20896
rect 15108 20800 15160 20806
rect 15160 20748 15240 20754
rect 15108 20742 15240 20748
rect 15120 20726 15240 20742
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15016 19780 15068 19786
rect 15016 19722 15068 19728
rect 15028 18766 15056 19722
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 15016 18760 15068 18766
rect 15016 18702 15068 18708
rect 15014 18048 15070 18057
rect 15014 17983 15070 17992
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14660 12238 14688 12582
rect 14752 12238 14780 13126
rect 14844 12850 14872 17614
rect 15028 17202 15056 17983
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15014 16688 15070 16697
rect 15014 16623 15070 16632
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14936 16250 14964 16458
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15028 16114 15056 16623
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14618 14964 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15028 14482 15056 15438
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15120 14362 15148 20470
rect 15028 14334 15148 14362
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 10742 14688 12038
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14200 9646 14596 9674
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14108 3534 14136 4558
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14016 2106 14044 2246
rect 14004 2100 14056 2106
rect 14004 2042 14056 2048
rect 14200 2009 14228 9646
rect 14372 8968 14424 8974
rect 14370 8936 14372 8945
rect 14424 8936 14426 8945
rect 14370 8871 14426 8880
rect 14660 8498 14688 10678
rect 14752 8498 14780 10678
rect 14844 8838 14872 12786
rect 14936 12073 14964 13670
rect 14922 12064 14978 12073
rect 14922 11999 14978 12008
rect 14936 11762 14964 11999
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14922 9072 14978 9081
rect 14922 9007 14978 9016
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14660 7410 14688 8434
rect 14752 7478 14780 8434
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 5370 14412 7278
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14476 5914 14504 7142
rect 14738 5944 14794 5953
rect 14464 5908 14516 5914
rect 14738 5879 14740 5888
rect 14464 5850 14516 5856
rect 14792 5879 14794 5888
rect 14740 5850 14792 5856
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14370 4720 14426 4729
rect 14370 4655 14372 4664
rect 14424 4655 14426 4664
rect 14372 4626 14424 4632
rect 14384 4146 14412 4626
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3194 14320 3470
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14476 2514 14504 4762
rect 14568 4554 14596 4966
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14752 4282 14780 5850
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14844 3534 14872 8774
rect 14936 5914 14964 9007
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14936 5166 14964 5646
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14936 5001 14964 5102
rect 14922 4992 14978 5001
rect 14922 4927 14978 4936
rect 14924 4616 14976 4622
rect 14922 4584 14924 4593
rect 14976 4584 14978 4593
rect 14922 4519 14978 4528
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14372 2440 14424 2446
rect 14278 2408 14334 2417
rect 14372 2382 14424 2388
rect 14278 2343 14334 2352
rect 14186 2000 14242 2009
rect 14292 1970 14320 2343
rect 14186 1935 14242 1944
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14004 1828 14056 1834
rect 14004 1770 14056 1776
rect 14016 1358 14044 1770
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 13912 1352 13964 1358
rect 13912 1294 13964 1300
rect 14004 1352 14056 1358
rect 14004 1294 14056 1300
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 14016 160 14044 1158
rect 14292 160 14320 1702
rect 14384 610 14412 2382
rect 15028 1902 15056 14334
rect 15212 13433 15240 20726
rect 15304 17678 15332 21134
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15396 20602 15424 20946
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15396 16538 15424 19926
rect 15488 16572 15516 21490
rect 15580 18714 15608 26438
rect 15936 26386 15988 26392
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15672 26042 15700 26318
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15856 25922 15884 26250
rect 15948 26042 15976 26386
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 16040 26042 16068 26250
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16028 26036 16080 26042
rect 16028 25978 16080 25984
rect 15934 25936 15990 25945
rect 15856 25894 15934 25922
rect 15934 25871 15990 25880
rect 15785 25596 16093 25605
rect 15785 25594 15791 25596
rect 15847 25594 15871 25596
rect 15927 25594 15951 25596
rect 16007 25594 16031 25596
rect 16087 25594 16093 25596
rect 15847 25542 15849 25594
rect 16029 25542 16031 25594
rect 15785 25540 15791 25542
rect 15847 25540 15871 25542
rect 15927 25540 15951 25542
rect 16007 25540 16031 25542
rect 16087 25540 16093 25542
rect 15785 25531 16093 25540
rect 15934 25256 15990 25265
rect 16132 25242 16160 28494
rect 16224 27577 16252 28902
rect 16210 27568 16266 27577
rect 16210 27503 16212 27512
rect 16264 27503 16266 27512
rect 16212 27474 16264 27480
rect 15990 25214 16160 25242
rect 15934 25191 15990 25200
rect 16118 25120 16174 25129
rect 16118 25055 16174 25064
rect 15785 24508 16093 24517
rect 15785 24506 15791 24508
rect 15847 24506 15871 24508
rect 15927 24506 15951 24508
rect 16007 24506 16031 24508
rect 16087 24506 16093 24508
rect 15847 24454 15849 24506
rect 16029 24454 16031 24506
rect 15785 24452 15791 24454
rect 15847 24452 15871 24454
rect 15927 24452 15951 24454
rect 16007 24452 16031 24454
rect 16087 24452 16093 24454
rect 15785 24443 16093 24452
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 15672 23866 15700 24210
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15948 23866 15976 24142
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15785 23420 16093 23429
rect 15785 23418 15791 23420
rect 15847 23418 15871 23420
rect 15927 23418 15951 23420
rect 16007 23418 16031 23420
rect 16087 23418 16093 23420
rect 15847 23366 15849 23418
rect 16029 23366 16031 23418
rect 15785 23364 15791 23366
rect 15847 23364 15871 23366
rect 15927 23364 15951 23366
rect 16007 23364 16031 23366
rect 16087 23364 16093 23366
rect 15785 23355 16093 23364
rect 15660 22432 15712 22438
rect 15660 22374 15712 22380
rect 15672 22216 15700 22374
rect 15785 22332 16093 22341
rect 15785 22330 15791 22332
rect 15847 22330 15871 22332
rect 15927 22330 15951 22332
rect 16007 22330 16031 22332
rect 16087 22330 16093 22332
rect 15847 22278 15849 22330
rect 16029 22278 16031 22330
rect 15785 22276 15791 22278
rect 15847 22276 15871 22278
rect 15927 22276 15951 22278
rect 16007 22276 16031 22278
rect 16087 22276 16093 22278
rect 15785 22267 16093 22276
rect 15672 22188 15884 22216
rect 15750 22128 15806 22137
rect 15750 22063 15806 22072
rect 15764 21332 15792 22063
rect 15856 21554 15884 22188
rect 16132 22094 16160 25055
rect 16132 22066 16252 22094
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16132 21622 16160 21966
rect 16120 21616 16172 21622
rect 16120 21558 16172 21564
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15672 21304 15792 21332
rect 16120 21344 16172 21350
rect 15672 21026 15700 21304
rect 16120 21286 16172 21292
rect 15785 21244 16093 21253
rect 15785 21242 15791 21244
rect 15847 21242 15871 21244
rect 15927 21242 15951 21244
rect 16007 21242 16031 21244
rect 16087 21242 16093 21244
rect 15847 21190 15849 21242
rect 16029 21190 16031 21242
rect 15785 21188 15791 21190
rect 15847 21188 15871 21190
rect 15927 21188 15951 21190
rect 16007 21188 16031 21190
rect 16087 21188 16093 21190
rect 15785 21179 16093 21188
rect 15672 21010 15792 21026
rect 16132 21010 16160 21286
rect 15672 21004 15804 21010
rect 15672 20998 15752 21004
rect 15752 20946 15804 20952
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 15785 20156 16093 20165
rect 15785 20154 15791 20156
rect 15847 20154 15871 20156
rect 15927 20154 15951 20156
rect 16007 20154 16031 20156
rect 16087 20154 16093 20156
rect 15847 20102 15849 20154
rect 16029 20102 16031 20154
rect 15785 20100 15791 20102
rect 15847 20100 15871 20102
rect 15927 20100 15951 20102
rect 16007 20100 16031 20102
rect 16087 20100 16093 20102
rect 15785 20091 16093 20100
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16132 19174 16160 19994
rect 16224 19417 16252 22066
rect 16316 20040 16344 41958
rect 16960 41721 16988 42026
rect 16946 41712 17002 41721
rect 16946 41647 17002 41656
rect 17052 41585 17080 42162
rect 17316 42084 17368 42090
rect 17316 42026 17368 42032
rect 17328 41857 17356 42026
rect 17314 41848 17370 41857
rect 17314 41783 17370 41792
rect 17038 41576 17094 41585
rect 17038 41511 17094 41520
rect 16396 41064 16448 41070
rect 16396 41006 16448 41012
rect 16408 40730 16436 41006
rect 16396 40724 16448 40730
rect 16396 40666 16448 40672
rect 17420 40458 17448 43250
rect 17512 43110 17540 43590
rect 17604 43330 17632 44463
rect 17880 43466 17908 44463
rect 18156 43858 18184 44463
rect 18144 43852 18196 43858
rect 18144 43794 18196 43800
rect 18432 43738 18460 44463
rect 18616 44418 18644 44503
rect 18694 44463 18750 44623
rect 18970 44463 19026 44623
rect 19246 44463 19302 44623
rect 19522 44463 19578 44623
rect 19798 44463 19854 44623
rect 20074 44463 20130 44623
rect 20350 44463 20406 44623
rect 20626 44463 20682 44623
rect 20902 44463 20958 44623
rect 21178 44463 21234 44623
rect 21454 44463 21510 44623
rect 21730 44463 21786 44623
rect 22006 44463 22062 44623
rect 22282 44463 22338 44623
rect 22558 44463 22614 44623
rect 22834 44463 22890 44623
rect 23110 44463 23166 44623
rect 23386 44463 23442 44623
rect 23662 44463 23718 44623
rect 23938 44463 23994 44623
rect 24214 44463 24270 44623
rect 24490 44463 24546 44623
rect 24766 44463 24822 44623
rect 25042 44463 25098 44623
rect 25318 44463 25374 44623
rect 25594 44463 25650 44623
rect 18708 44418 18736 44463
rect 18616 44390 18736 44418
rect 18432 43722 18552 43738
rect 18432 43716 18564 43722
rect 18432 43710 18512 43716
rect 18984 43704 19012 44463
rect 18984 43676 19196 43704
rect 18512 43658 18564 43664
rect 18752 43548 19060 43557
rect 18752 43546 18758 43548
rect 18814 43546 18838 43548
rect 18894 43546 18918 43548
rect 18974 43546 18998 43548
rect 19054 43546 19060 43548
rect 18814 43494 18816 43546
rect 18996 43494 18998 43546
rect 18752 43492 18758 43494
rect 18814 43492 18838 43494
rect 18894 43492 18918 43494
rect 18974 43492 18998 43494
rect 19054 43492 19060 43494
rect 18752 43483 19060 43492
rect 17880 43450 18184 43466
rect 17880 43444 18196 43450
rect 17880 43438 18144 43444
rect 18144 43386 18196 43392
rect 18236 43376 18288 43382
rect 17604 43324 18236 43330
rect 17604 43318 18288 43324
rect 17604 43302 18276 43318
rect 18328 43172 18380 43178
rect 18328 43114 18380 43120
rect 17500 43104 17552 43110
rect 17500 43046 17552 43052
rect 17592 43104 17644 43110
rect 17592 43046 17644 43052
rect 17684 43104 17736 43110
rect 17684 43046 17736 43052
rect 18144 43104 18196 43110
rect 18144 43046 18196 43052
rect 17604 42702 17632 43046
rect 17696 42906 17724 43046
rect 18156 42906 18184 43046
rect 17684 42900 17736 42906
rect 17684 42842 17736 42848
rect 18144 42900 18196 42906
rect 18144 42842 18196 42848
rect 18052 42832 18104 42838
rect 18052 42774 18104 42780
rect 17592 42696 17644 42702
rect 17592 42638 17644 42644
rect 17776 42560 17828 42566
rect 17776 42502 17828 42508
rect 17788 42362 17816 42502
rect 17776 42356 17828 42362
rect 17776 42298 17828 42304
rect 18064 42294 18092 42774
rect 18340 42702 18368 43114
rect 18420 43104 18472 43110
rect 18420 43046 18472 43052
rect 18512 43104 18564 43110
rect 18512 43046 18564 43052
rect 18432 42770 18460 43046
rect 18420 42764 18472 42770
rect 18420 42706 18472 42712
rect 18328 42696 18380 42702
rect 18328 42638 18380 42644
rect 18418 42664 18474 42673
rect 18418 42599 18474 42608
rect 18236 42560 18288 42566
rect 18236 42502 18288 42508
rect 18328 42560 18380 42566
rect 18328 42502 18380 42508
rect 18052 42288 18104 42294
rect 18052 42230 18104 42236
rect 17684 42084 17736 42090
rect 17684 42026 17736 42032
rect 18052 42084 18104 42090
rect 18052 42026 18104 42032
rect 17696 41721 17724 42026
rect 17868 41812 17920 41818
rect 17868 41754 17920 41760
rect 17682 41712 17738 41721
rect 17682 41647 17738 41656
rect 17408 40452 17460 40458
rect 17408 40394 17460 40400
rect 16672 38820 16724 38826
rect 16672 38762 16724 38768
rect 16684 36786 16712 38762
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 17132 36576 17184 36582
rect 17132 36518 17184 36524
rect 17408 36576 17460 36582
rect 17408 36518 17460 36524
rect 17144 36378 17172 36518
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 17224 36168 17276 36174
rect 17224 36110 17276 36116
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 16408 32298 16436 34954
rect 16684 34678 16712 35158
rect 16672 34672 16724 34678
rect 16672 34614 16724 34620
rect 16764 34672 16816 34678
rect 16764 34614 16816 34620
rect 16776 34218 16804 34614
rect 16592 34190 16804 34218
rect 16592 33590 16620 34190
rect 16764 34128 16816 34134
rect 16764 34070 16816 34076
rect 16776 33658 16804 34070
rect 16868 33998 16896 35634
rect 17132 35216 17184 35222
rect 17132 35158 17184 35164
rect 17144 34678 17172 35158
rect 17132 34672 17184 34678
rect 17132 34614 17184 34620
rect 17236 34474 17264 36110
rect 17420 36106 17448 36518
rect 17880 36174 17908 41754
rect 17960 41744 18012 41750
rect 17960 41686 18012 41692
rect 17972 41546 18000 41686
rect 17960 41540 18012 41546
rect 17960 41482 18012 41488
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 17408 36100 17460 36106
rect 17408 36042 17460 36048
rect 17776 36100 17828 36106
rect 17776 36042 17828 36048
rect 17592 35624 17644 35630
rect 17592 35566 17644 35572
rect 17604 35222 17632 35566
rect 17592 35216 17644 35222
rect 17592 35158 17644 35164
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17224 34468 17276 34474
rect 17224 34410 17276 34416
rect 16856 33992 16908 33998
rect 16856 33934 16908 33940
rect 17038 33960 17094 33969
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 16580 33584 16632 33590
rect 16580 33526 16632 33532
rect 16868 32842 16896 33934
rect 17038 33895 17040 33904
rect 17092 33895 17094 33904
rect 17040 33866 17092 33872
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16672 32360 16724 32366
rect 16672 32302 16724 32308
rect 16396 32292 16448 32298
rect 16396 32234 16448 32240
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16592 31906 16620 32166
rect 16500 31878 16620 31906
rect 16500 31822 16528 31878
rect 16488 31816 16540 31822
rect 16488 31758 16540 31764
rect 16684 31754 16712 32302
rect 16960 31890 16988 33798
rect 17236 33522 17264 34410
rect 17512 34202 17540 34546
rect 17500 34196 17552 34202
rect 17500 34138 17552 34144
rect 17316 34060 17368 34066
rect 17316 34002 17368 34008
rect 17328 33522 17356 34002
rect 17500 33992 17552 33998
rect 17500 33934 17552 33940
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 17316 33516 17368 33522
rect 17316 33458 17368 33464
rect 17040 32224 17092 32230
rect 17040 32166 17092 32172
rect 16948 31884 17000 31890
rect 16948 31826 17000 31832
rect 16592 31726 16712 31754
rect 16488 31340 16540 31346
rect 16488 31282 16540 31288
rect 16396 30592 16448 30598
rect 16396 30534 16448 30540
rect 16408 20262 16436 30534
rect 16500 30258 16528 31282
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 16500 27418 16528 30194
rect 16592 29646 16620 31726
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16592 27713 16620 29582
rect 16684 29510 16712 30670
rect 16960 29714 16988 31826
rect 16948 29708 17000 29714
rect 16948 29650 17000 29656
rect 16762 29608 16818 29617
rect 17052 29594 17080 32166
rect 17144 31890 17172 33458
rect 17328 32978 17356 33458
rect 17316 32972 17368 32978
rect 17316 32914 17368 32920
rect 17408 32904 17460 32910
rect 17328 32852 17408 32858
rect 17328 32846 17460 32852
rect 17328 32830 17448 32846
rect 17132 31884 17184 31890
rect 17132 31826 17184 31832
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17132 31136 17184 31142
rect 17132 31078 17184 31084
rect 17144 29714 17172 31078
rect 17132 29708 17184 29714
rect 17132 29650 17184 29656
rect 16762 29543 16818 29552
rect 16960 29566 17080 29594
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16672 28620 16724 28626
rect 16672 28562 16724 28568
rect 16684 28218 16712 28562
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16672 27940 16724 27946
rect 16672 27882 16724 27888
rect 16578 27704 16634 27713
rect 16578 27639 16634 27648
rect 16500 27390 16620 27418
rect 16488 27328 16540 27334
rect 16486 27296 16488 27305
rect 16540 27296 16542 27305
rect 16486 27231 16542 27240
rect 16500 26042 16528 27231
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16486 25936 16542 25945
rect 16592 25922 16620 27390
rect 16542 25894 16620 25922
rect 16486 25871 16542 25880
rect 16684 25344 16712 27882
rect 16776 26994 16804 29543
rect 16854 29472 16910 29481
rect 16854 29407 16910 29416
rect 16868 29170 16896 29407
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16960 28558 16988 29566
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16856 26920 16908 26926
rect 16856 26862 16908 26868
rect 16868 26246 16896 26862
rect 16856 26240 16908 26246
rect 16856 26182 16908 26188
rect 16868 25378 16896 26182
rect 16776 25362 16896 25378
rect 16592 25316 16712 25344
rect 16764 25356 16896 25362
rect 16592 24818 16620 25316
rect 16816 25350 16896 25356
rect 16764 25298 16816 25304
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16500 22030 16528 23734
rect 16592 22642 16620 24754
rect 16684 22710 16712 25162
rect 16764 24880 16816 24886
rect 16764 24822 16816 24828
rect 16776 24138 16804 24822
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16776 23322 16804 24074
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16672 22704 16724 22710
rect 16672 22646 16724 22652
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16500 21593 16528 21966
rect 16486 21584 16542 21593
rect 16486 21519 16542 21528
rect 16592 21536 16620 22578
rect 16684 22148 16712 22646
rect 16776 22574 16804 23054
rect 16764 22568 16816 22574
rect 16764 22510 16816 22516
rect 16960 22438 16988 28494
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16684 22120 16988 22148
rect 16960 22012 16988 22120
rect 17052 22080 17080 29446
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17144 27985 17172 28494
rect 17130 27976 17186 27985
rect 17130 27911 17186 27920
rect 17144 22982 17172 27911
rect 17236 27470 17264 31418
rect 17328 27946 17356 32830
rect 17408 31136 17460 31142
rect 17408 31078 17460 31084
rect 17420 30938 17448 31078
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17512 29850 17540 33934
rect 17604 32978 17632 35158
rect 17788 34105 17816 36042
rect 17972 35086 18000 36518
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17774 34096 17830 34105
rect 17774 34031 17830 34040
rect 17592 32972 17644 32978
rect 17592 32914 17644 32920
rect 17604 30190 17632 32914
rect 17684 32428 17736 32434
rect 17684 32370 17736 32376
rect 17696 30802 17724 32370
rect 17788 31346 17816 34031
rect 17880 32910 17908 34546
rect 17958 33280 18014 33289
rect 17958 33215 18014 33224
rect 17868 32904 17920 32910
rect 17868 32846 17920 32852
rect 17972 31482 18000 33215
rect 17960 31476 18012 31482
rect 17960 31418 18012 31424
rect 17776 31340 17828 31346
rect 17776 31282 17828 31288
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17972 30938 18000 31282
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17592 30184 17644 30190
rect 17592 30126 17644 30132
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17590 29336 17646 29345
rect 17590 29271 17646 29280
rect 17408 28960 17460 28966
rect 17408 28902 17460 28908
rect 17420 28626 17448 28902
rect 17408 28620 17460 28626
rect 17408 28562 17460 28568
rect 17498 28112 17554 28121
rect 17498 28047 17554 28056
rect 17316 27940 17368 27946
rect 17316 27882 17368 27888
rect 17314 27568 17370 27577
rect 17314 27503 17316 27512
rect 17368 27503 17370 27512
rect 17316 27474 17368 27480
rect 17224 27464 17276 27470
rect 17222 27432 17224 27441
rect 17276 27432 17278 27441
rect 17222 27367 17278 27376
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 17236 26926 17264 27270
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17328 26761 17356 27474
rect 17408 26784 17460 26790
rect 17314 26752 17370 26761
rect 17408 26726 17460 26732
rect 17314 26687 17370 26696
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17052 22052 17172 22080
rect 16960 21984 17080 22012
rect 16854 21856 16910 21865
rect 16854 21791 16910 21800
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16592 21508 16712 21536
rect 16486 21448 16542 21457
rect 16542 21406 16620 21434
rect 16486 21383 16542 21392
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16592 20058 16620 21406
rect 16684 20942 16712 21508
rect 16776 21010 16804 21558
rect 16868 21486 16896 21791
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16764 21004 16816 21010
rect 16764 20946 16816 20952
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 16868 20788 16896 21422
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16776 20760 16896 20788
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16580 20052 16632 20058
rect 16316 20012 16528 20040
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16210 19408 16266 19417
rect 16210 19343 16266 19352
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 15785 19068 16093 19077
rect 15785 19066 15791 19068
rect 15847 19066 15871 19068
rect 15927 19066 15951 19068
rect 16007 19066 16031 19068
rect 16087 19066 16093 19068
rect 15847 19014 15849 19066
rect 16029 19014 16031 19066
rect 15785 19012 15791 19014
rect 15847 19012 15871 19014
rect 15927 19012 15951 19014
rect 16007 19012 16031 19014
rect 16087 19012 16093 19014
rect 15785 19003 16093 19012
rect 16132 18970 16160 19110
rect 16316 18970 16344 19858
rect 16408 19378 16436 19858
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16212 18760 16264 18766
rect 16210 18728 16212 18737
rect 16264 18728 16266 18737
rect 15580 18686 15700 18714
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18057 15608 18566
rect 15566 18048 15622 18057
rect 15566 17983 15622 17992
rect 15672 16776 15700 18686
rect 15752 18692 15804 18698
rect 16210 18663 16266 18672
rect 15752 18634 15804 18640
rect 15764 18290 15792 18634
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15785 17980 16093 17989
rect 15785 17978 15791 17980
rect 15847 17978 15871 17980
rect 15927 17978 15951 17980
rect 16007 17978 16031 17980
rect 16087 17978 16093 17980
rect 15847 17926 15849 17978
rect 16029 17926 16031 17978
rect 15785 17924 15791 17926
rect 15847 17924 15871 17926
rect 15927 17924 15951 17926
rect 16007 17924 16031 17926
rect 16087 17924 16093 17926
rect 15785 17915 16093 17924
rect 15785 16892 16093 16901
rect 15785 16890 15791 16892
rect 15847 16890 15871 16892
rect 15927 16890 15951 16892
rect 16007 16890 16031 16892
rect 16087 16890 16093 16892
rect 15847 16838 15849 16890
rect 16029 16838 16031 16890
rect 15785 16836 15791 16838
rect 15847 16836 15871 16838
rect 15927 16836 15951 16838
rect 16007 16836 16031 16838
rect 16087 16836 16093 16838
rect 15785 16827 16093 16836
rect 16132 16794 16160 18022
rect 16302 17912 16358 17921
rect 16302 17847 16358 17856
rect 16316 17678 16344 17847
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16304 17196 16356 17202
rect 16356 17156 16436 17184
rect 16304 17138 16356 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16120 16788 16172 16794
rect 15672 16748 15792 16776
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15568 16584 15620 16590
rect 15488 16544 15568 16572
rect 15304 16510 15424 16538
rect 15568 16526 15620 16532
rect 15304 15026 15332 16510
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15304 14521 15332 14554
rect 15290 14512 15346 14521
rect 15290 14447 15346 14456
rect 15198 13424 15254 13433
rect 15198 13359 15254 13368
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 15120 10742 15148 12038
rect 15304 11880 15332 13262
rect 15396 12238 15424 16390
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 14074 15516 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 12442 15516 13670
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15212 11852 15332 11880
rect 15384 11892 15436 11898
rect 15212 11762 15240 11852
rect 15384 11834 15436 11840
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15212 10305 15240 11698
rect 15304 11014 15332 11698
rect 15396 11354 15424 11834
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15396 10962 15424 11018
rect 15488 10962 15516 12174
rect 15396 10934 15516 10962
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15120 9450 15148 9658
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 8634 15148 8774
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 6322 15148 6598
rect 15212 6322 15240 10231
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 7041 15332 9658
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15290 7032 15346 7041
rect 15290 6967 15346 6976
rect 15396 6866 15424 7822
rect 15488 6934 15516 10934
rect 15580 8430 15608 16526
rect 15672 9625 15700 16594
rect 15764 15910 15792 16748
rect 16120 16730 16172 16736
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16040 16561 16068 16594
rect 16026 16552 16082 16561
rect 16026 16487 16082 16496
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15785 15804 16093 15813
rect 15785 15802 15791 15804
rect 15847 15802 15871 15804
rect 15927 15802 15951 15804
rect 16007 15802 16031 15804
rect 16087 15802 16093 15804
rect 15847 15750 15849 15802
rect 16029 15750 16031 15802
rect 15785 15748 15791 15750
rect 15847 15748 15871 15750
rect 15927 15748 15951 15750
rect 16007 15748 16031 15750
rect 16087 15748 16093 15750
rect 15785 15739 16093 15748
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 15785 14716 16093 14725
rect 15785 14714 15791 14716
rect 15847 14714 15871 14716
rect 15927 14714 15951 14716
rect 16007 14714 16031 14716
rect 16087 14714 16093 14716
rect 15847 14662 15849 14714
rect 16029 14662 16031 14714
rect 15785 14660 15791 14662
rect 15847 14660 15871 14662
rect 15927 14660 15951 14662
rect 16007 14660 16031 14662
rect 16087 14660 16093 14662
rect 15785 14651 16093 14660
rect 16224 14657 16252 14826
rect 16210 14648 16266 14657
rect 16210 14583 16266 14592
rect 16224 14550 16252 14583
rect 16212 14544 16264 14550
rect 16026 14512 16082 14521
rect 16316 14521 16344 16730
rect 16212 14486 16264 14492
rect 16302 14512 16358 14521
rect 16026 14447 16028 14456
rect 16080 14447 16082 14456
rect 16028 14418 16080 14424
rect 16040 13734 16068 14418
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15785 13628 16093 13637
rect 15785 13626 15791 13628
rect 15847 13626 15871 13628
rect 15927 13626 15951 13628
rect 16007 13626 16031 13628
rect 16087 13626 16093 13628
rect 15847 13574 15849 13626
rect 16029 13574 16031 13626
rect 15785 13572 15791 13574
rect 15847 13572 15871 13574
rect 15927 13572 15951 13574
rect 16007 13572 16031 13574
rect 16087 13572 16093 13574
rect 15785 13563 16093 13572
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 15785 12540 16093 12549
rect 15785 12538 15791 12540
rect 15847 12538 15871 12540
rect 15927 12538 15951 12540
rect 16007 12538 16031 12540
rect 16087 12538 16093 12540
rect 15847 12486 15849 12538
rect 16029 12486 16031 12538
rect 15785 12484 15791 12486
rect 15847 12484 15871 12486
rect 15927 12484 15951 12486
rect 16007 12484 16031 12486
rect 16087 12484 16093 12486
rect 15785 12475 16093 12484
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15842 12064 15898 12073
rect 15764 11694 15792 12038
rect 15842 11999 15898 12008
rect 15856 11694 15884 11999
rect 16132 11694 16160 12718
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15785 11452 16093 11461
rect 15785 11450 15791 11452
rect 15847 11450 15871 11452
rect 15927 11450 15951 11452
rect 16007 11450 16031 11452
rect 16087 11450 16093 11452
rect 15847 11398 15849 11450
rect 16029 11398 16031 11450
rect 15785 11396 15791 11398
rect 15847 11396 15871 11398
rect 15927 11396 15951 11398
rect 16007 11396 16031 11398
rect 16087 11396 16093 11398
rect 15785 11387 16093 11396
rect 16224 11218 16252 14486
rect 16302 14447 16358 14456
rect 16408 14362 16436 17156
rect 16500 15178 16528 20012
rect 16580 19994 16632 20000
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16592 15609 16620 18566
rect 16578 15600 16634 15609
rect 16578 15535 16634 15544
rect 16500 15150 16620 15178
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16316 14334 16436 14362
rect 16316 11762 16344 14334
rect 16500 12238 16528 14418
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15785 10364 16093 10373
rect 15785 10362 15791 10364
rect 15847 10362 15871 10364
rect 15927 10362 15951 10364
rect 16007 10362 16031 10364
rect 16087 10362 16093 10364
rect 15847 10310 15849 10362
rect 16029 10310 16031 10362
rect 15785 10308 15791 10310
rect 15847 10308 15871 10310
rect 15927 10308 15951 10310
rect 16007 10308 16031 10310
rect 16087 10308 16093 10310
rect 15785 10299 16093 10308
rect 15658 9616 15714 9625
rect 15658 9551 15714 9560
rect 15672 8566 15700 9551
rect 15785 9276 16093 9285
rect 15785 9274 15791 9276
rect 15847 9274 15871 9276
rect 15927 9274 15951 9276
rect 16007 9274 16031 9276
rect 16087 9274 16093 9276
rect 15847 9222 15849 9274
rect 16029 9222 16031 9274
rect 15785 9220 15791 9222
rect 15847 9220 15871 9222
rect 15927 9220 15951 9222
rect 16007 9220 16031 9222
rect 16087 9220 16093 9222
rect 15785 9211 16093 9220
rect 15750 9072 15806 9081
rect 16132 9058 16160 11086
rect 16224 10810 16252 11154
rect 16592 11098 16620 15150
rect 16684 14890 16712 20538
rect 16776 16794 16804 20760
rect 16960 20466 16988 20946
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16868 19514 16896 19790
rect 16960 19718 16988 20402
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 17052 18222 17080 21984
rect 17144 21350 17172 22052
rect 17236 22030 17264 25978
rect 17420 25362 17448 26726
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17408 25356 17460 25362
rect 17408 25298 17460 25304
rect 17328 24954 17356 25298
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17316 24200 17368 24206
rect 17314 24168 17316 24177
rect 17368 24168 17370 24177
rect 17314 24103 17370 24112
rect 17420 23118 17448 25298
rect 17512 25140 17540 28047
rect 17604 26926 17632 29271
rect 17696 28014 17724 30738
rect 17960 30320 18012 30326
rect 17960 30262 18012 30268
rect 17868 30184 17920 30190
rect 17868 30126 17920 30132
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17788 29782 17816 29990
rect 17776 29776 17828 29782
rect 17776 29718 17828 29724
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17592 26920 17644 26926
rect 17592 26862 17644 26868
rect 17604 25673 17632 26862
rect 17696 26382 17724 27950
rect 17788 27418 17816 29582
rect 17880 29510 17908 30126
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17880 29170 17908 29446
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17972 29034 18000 30262
rect 17960 29028 18012 29034
rect 17960 28970 18012 28976
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17972 28082 18000 28494
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17788 27390 18000 27418
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17880 26994 17908 27270
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17590 25664 17646 25673
rect 17590 25599 17646 25608
rect 17592 25288 17644 25294
rect 17590 25256 17592 25265
rect 17644 25256 17646 25265
rect 17590 25191 17646 25200
rect 17512 25112 17632 25140
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17316 22500 17368 22506
rect 17316 22442 17368 22448
rect 17328 22234 17356 22442
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17328 21604 17356 22170
rect 17234 21576 17356 21604
rect 17234 21536 17262 21576
rect 17234 21508 17264 21536
rect 17236 21468 17264 21508
rect 17316 21480 17368 21486
rect 17236 21440 17316 21468
rect 17316 21422 17368 21428
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17144 20602 17172 21286
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 17144 17746 17172 18702
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 17052 17202 17080 17274
rect 17144 17270 17172 17682
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16868 16794 16896 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16776 16658 16804 16730
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16868 16538 16896 16730
rect 16776 16510 16896 16538
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16776 14521 16804 16510
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15706 16896 15846
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16762 14512 16818 14521
rect 16762 14447 16818 14456
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16762 14240 16818 14249
rect 16762 14175 16818 14184
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16684 13138 16712 13942
rect 16776 13734 16804 14175
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13326 16804 13670
rect 16868 13530 16896 14418
rect 16960 13938 16988 15098
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16684 13110 16896 13138
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11354 16804 12174
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 16408 11070 16620 11098
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16316 9722 16344 10950
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16132 9030 16252 9058
rect 15750 9007 15806 9016
rect 15764 8974 15792 9007
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15580 7954 15608 8366
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15672 7886 15700 8502
rect 15785 8188 16093 8197
rect 15785 8186 15791 8188
rect 15847 8186 15871 8188
rect 15927 8186 15951 8188
rect 16007 8186 16031 8188
rect 16087 8186 16093 8188
rect 15847 8134 15849 8186
rect 16029 8134 16031 8186
rect 15785 8132 15791 8134
rect 15847 8132 15871 8134
rect 15927 8132 15951 8134
rect 16007 8132 16031 8134
rect 16087 8132 16093 8134
rect 15785 8123 16093 8132
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15658 7712 15714 7721
rect 15658 7647 15714 7656
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15120 4690 15148 6258
rect 15396 5914 15424 6802
rect 15488 6798 15516 6870
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5137 15240 5510
rect 15304 5370 15332 5714
rect 15396 5642 15424 5714
rect 15488 5710 15516 6394
rect 15566 6352 15622 6361
rect 15566 6287 15622 6296
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15396 5166 15424 5578
rect 15384 5160 15436 5166
rect 15198 5128 15254 5137
rect 15384 5102 15436 5108
rect 15198 5063 15254 5072
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15304 4282 15332 5034
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15580 4078 15608 6287
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15672 3058 15700 7647
rect 15785 7100 16093 7109
rect 15785 7098 15791 7100
rect 15847 7098 15871 7100
rect 15927 7098 15951 7100
rect 16007 7098 16031 7100
rect 16087 7098 16093 7100
rect 15847 7046 15849 7098
rect 16029 7046 16031 7098
rect 15785 7044 15791 7046
rect 15847 7044 15871 7046
rect 15927 7044 15951 7046
rect 16007 7044 16031 7046
rect 16087 7044 16093 7046
rect 15785 7035 16093 7044
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15764 5234 15792 5306
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 16132 4622 16160 8774
rect 16224 7993 16252 9030
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16210 7984 16266 7993
rect 16210 7919 16266 7928
rect 16224 7886 16252 7919
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16224 5794 16252 7822
rect 16316 7274 16344 8570
rect 16408 7562 16436 11070
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8090 16528 8774
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16408 7534 16528 7562
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16304 6112 16356 6118
rect 16304 6054 16356 6060
rect 16316 5914 16344 6054
rect 16408 5914 16436 6258
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16224 5778 16344 5794
rect 16224 5772 16356 5778
rect 16224 5766 16304 5772
rect 16304 5714 16356 5720
rect 16316 5370 16344 5714
rect 16394 5672 16450 5681
rect 16394 5607 16450 5616
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16408 5250 16436 5607
rect 16224 5222 16436 5250
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16224 4162 16252 5222
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16316 4826 16344 5034
rect 16408 4826 16436 5102
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16316 4282 16344 4762
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16132 4134 16252 4162
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15476 2848 15528 2854
rect 15528 2808 15608 2836
rect 15476 2790 15528 2796
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15396 2446 15424 2586
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 15120 2106 15148 2314
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 15016 1896 15068 1902
rect 15016 1838 15068 1844
rect 15200 1828 15252 1834
rect 15200 1770 15252 1776
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14372 604 14424 610
rect 14372 546 14424 552
rect 10414 54 10548 82
rect 10414 0 10470 54
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11242 0 11298 160
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 82 14610 160
rect 14752 82 14780 1702
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 14936 626 14964 1498
rect 15108 1488 15160 1494
rect 15108 1430 15160 1436
rect 14844 598 14964 626
rect 14844 160 14872 598
rect 15120 160 15148 1430
rect 15212 1358 15240 1770
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15396 160 15424 1770
rect 15488 1358 15516 2246
rect 15580 2038 15608 2808
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15785 2683 16093 2692
rect 16132 2650 16160 4134
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16224 2446 16252 4014
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16316 2689 16344 3470
rect 16302 2680 16358 2689
rect 16302 2615 16358 2624
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 15568 2032 15620 2038
rect 15568 1974 15620 1980
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15476 1352 15528 1358
rect 15476 1294 15528 1300
rect 15672 160 15700 1702
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16316 1562 16344 1838
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16396 1556 16448 1562
rect 16396 1498 16448 1504
rect 16408 626 16436 1498
rect 16500 1358 16528 7534
rect 16592 1902 16620 9658
rect 16776 8072 16804 11290
rect 16868 8242 16896 13110
rect 17052 12850 17080 17138
rect 17236 15502 17264 21286
rect 17314 21176 17370 21185
rect 17314 21111 17370 21120
rect 17328 16794 17356 21111
rect 17420 18222 17448 22918
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17420 16454 17448 18158
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17144 14929 17172 15370
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17236 15026 17264 15302
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17408 15020 17460 15026
rect 17512 15008 17540 24006
rect 17460 14980 17540 15008
rect 17408 14962 17460 14968
rect 17130 14920 17186 14929
rect 17130 14855 17186 14864
rect 17144 14600 17172 14855
rect 17110 14572 17172 14600
rect 17110 14498 17138 14572
rect 17222 14512 17278 14521
rect 17110 14482 17172 14498
rect 17110 14476 17184 14482
rect 17110 14470 17132 14476
rect 17222 14447 17224 14456
rect 17132 14418 17184 14424
rect 17276 14447 17278 14456
rect 17224 14418 17276 14424
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17420 14074 17448 14350
rect 17512 14278 17540 14980
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11898 17080 12242
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11082 16988 11494
rect 17040 11280 17092 11286
rect 17038 11248 17040 11257
rect 17092 11248 17094 11257
rect 17038 11183 17094 11192
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 17144 8922 17172 13330
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17236 9178 17264 11018
rect 17328 10169 17356 12174
rect 17420 11150 17448 13874
rect 17604 12434 17632 25112
rect 17696 24342 17724 26318
rect 17788 24614 17816 26862
rect 17972 26330 18000 27390
rect 17880 26302 18000 26330
rect 17880 24818 17908 26302
rect 17960 26240 18012 26246
rect 17960 26182 18012 26188
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17788 22642 17816 24550
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17880 23730 17908 24278
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17696 19922 17724 21830
rect 17774 21584 17830 21593
rect 17774 21519 17776 21528
rect 17828 21519 17830 21528
rect 17776 21490 17828 21496
rect 17788 21350 17816 21490
rect 17880 21486 17908 22510
rect 17972 21729 18000 26182
rect 17958 21720 18014 21729
rect 17958 21655 18014 21664
rect 17868 21480 17920 21486
rect 18064 21434 18092 42026
rect 18248 41818 18276 42502
rect 18340 42362 18368 42502
rect 18328 42356 18380 42362
rect 18328 42298 18380 42304
rect 18432 42294 18460 42599
rect 18420 42288 18472 42294
rect 18420 42230 18472 42236
rect 18524 42106 18552 43046
rect 18880 42900 18932 42906
rect 18880 42842 18932 42848
rect 18972 42900 19024 42906
rect 19168 42888 19196 43676
rect 19260 43081 19288 44463
rect 19340 43308 19392 43314
rect 19392 43268 19472 43296
rect 19340 43250 19392 43256
rect 19246 43072 19302 43081
rect 19246 43007 19302 43016
rect 19168 42860 19334 42888
rect 18972 42842 19024 42848
rect 18892 42673 18920 42842
rect 18984 42702 19012 42842
rect 19306 42820 19334 42860
rect 19306 42792 19380 42820
rect 18972 42696 19024 42702
rect 18878 42664 18934 42673
rect 19248 42696 19300 42702
rect 18972 42638 19024 42644
rect 19168 42644 19248 42650
rect 19168 42638 19300 42644
rect 18878 42599 18934 42608
rect 19168 42622 19288 42638
rect 18604 42560 18656 42566
rect 18604 42502 18656 42508
rect 18616 42294 18644 42502
rect 18752 42460 19060 42469
rect 18752 42458 18758 42460
rect 18814 42458 18838 42460
rect 18894 42458 18918 42460
rect 18974 42458 18998 42460
rect 19054 42458 19060 42460
rect 18814 42406 18816 42458
rect 18996 42406 18998 42458
rect 18752 42404 18758 42406
rect 18814 42404 18838 42406
rect 18894 42404 18918 42406
rect 18974 42404 18998 42406
rect 19054 42404 19060 42406
rect 18752 42395 19060 42404
rect 18604 42288 18656 42294
rect 18604 42230 18656 42236
rect 18970 42256 19026 42265
rect 18970 42191 19026 42200
rect 18432 42078 18552 42106
rect 18328 42016 18380 42022
rect 18328 41958 18380 41964
rect 18236 41812 18288 41818
rect 18236 41754 18288 41760
rect 18340 41721 18368 41958
rect 18326 41712 18382 41721
rect 18326 41647 18382 41656
rect 18432 41614 18460 42078
rect 18512 42016 18564 42022
rect 18512 41958 18564 41964
rect 18236 41608 18288 41614
rect 18234 41576 18236 41585
rect 18420 41608 18472 41614
rect 18288 41576 18290 41585
rect 18420 41550 18472 41556
rect 18234 41511 18290 41520
rect 18144 41472 18196 41478
rect 18420 41472 18472 41478
rect 18144 41414 18196 41420
rect 18418 41440 18420 41449
rect 18472 41440 18474 41449
rect 18156 21457 18184 41414
rect 18418 41375 18474 41384
rect 18418 41168 18474 41177
rect 18418 41103 18474 41112
rect 18326 35864 18382 35873
rect 18326 35799 18382 35808
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 18248 35086 18276 35702
rect 18236 35080 18288 35086
rect 18236 35022 18288 35028
rect 18236 33856 18288 33862
rect 18236 33798 18288 33804
rect 18248 33658 18276 33798
rect 18236 33652 18288 33658
rect 18236 33594 18288 33600
rect 18236 30048 18288 30054
rect 18236 29990 18288 29996
rect 18248 25498 18276 29990
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 17868 21422 17920 21428
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17880 21146 17908 21422
rect 17972 21406 18092 21434
rect 18142 21448 18198 21457
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17696 17134 17724 18090
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16794 17724 16934
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 13394 17724 15438
rect 17788 15434 17816 19926
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 17882 17908 18090
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17338 17908 17478
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17880 16250 17908 16390
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17880 15366 17908 15982
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 12850 17724 13194
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17512 12406 17632 12434
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17512 10554 17540 12406
rect 17788 12322 17816 12582
rect 17604 12306 17816 12322
rect 17592 12300 17816 12306
rect 17644 12294 17816 12300
rect 17592 12242 17644 12248
rect 17880 12220 17908 14962
rect 17788 12192 17908 12220
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17420 10526 17540 10554
rect 17314 10160 17370 10169
rect 17314 10095 17370 10104
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17052 8894 17172 8922
rect 17052 8634 17080 8894
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16868 8214 17080 8242
rect 16856 8084 16908 8090
rect 16776 8044 16856 8072
rect 16670 6896 16726 6905
rect 16670 6831 16726 6840
rect 16684 2650 16712 6831
rect 16776 6458 16804 8044
rect 16856 8026 16908 8032
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 17052 5250 17080 8214
rect 17144 7954 17172 8774
rect 17328 8566 17356 10095
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 6662 17264 7686
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5370 17172 5714
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17222 5264 17278 5273
rect 17052 5222 17222 5250
rect 17222 5199 17278 5208
rect 17038 4856 17094 4865
rect 17038 4791 17094 4800
rect 16764 4208 16816 4214
rect 16764 4150 16816 4156
rect 16776 2650 16804 4150
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17052 2514 17080 4791
rect 17222 3904 17278 3913
rect 17222 3839 17278 3848
rect 17236 3534 17264 3839
rect 17328 3534 17356 8502
rect 17420 5545 17448 10526
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10266 17540 10406
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17604 10033 17632 11018
rect 17590 10024 17646 10033
rect 17590 9959 17646 9968
rect 17500 6384 17552 6390
rect 17500 6326 17552 6332
rect 17512 5817 17540 6326
rect 17498 5808 17554 5817
rect 17498 5743 17554 5752
rect 17512 5710 17540 5743
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17406 5536 17462 5545
rect 17406 5471 17462 5480
rect 17604 5302 17632 9959
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17696 6458 17724 9114
rect 17788 7818 17816 12192
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17880 11286 17908 11766
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17972 9722 18000 21406
rect 18142 21383 18198 21392
rect 18248 20534 18276 24754
rect 18340 21978 18368 35799
rect 18432 33289 18460 41103
rect 18418 33280 18474 33289
rect 18418 33215 18474 33224
rect 18524 33130 18552 41958
rect 18984 41614 19012 42191
rect 19168 41818 19196 42622
rect 19246 42256 19302 42265
rect 19246 42191 19302 42200
rect 19156 41812 19208 41818
rect 19156 41754 19208 41760
rect 18972 41608 19024 41614
rect 18972 41550 19024 41556
rect 18752 41372 19060 41381
rect 18752 41370 18758 41372
rect 18814 41370 18838 41372
rect 18894 41370 18918 41372
rect 18974 41370 18998 41372
rect 19054 41370 19060 41372
rect 18814 41318 18816 41370
rect 18996 41318 18998 41370
rect 18752 41316 18758 41318
rect 18814 41316 18838 41318
rect 18894 41316 18918 41318
rect 18974 41316 18998 41318
rect 19054 41316 19060 41318
rect 18752 41307 19060 41316
rect 19064 40928 19116 40934
rect 19064 40870 19116 40876
rect 19076 40730 19104 40870
rect 19064 40724 19116 40730
rect 19064 40666 19116 40672
rect 19260 40594 19288 42191
rect 19352 41478 19380 42792
rect 19444 41818 19472 43268
rect 19536 43194 19564 44463
rect 19536 43166 19656 43194
rect 19524 43104 19576 43110
rect 19524 43046 19576 43052
rect 19536 42294 19564 43046
rect 19524 42288 19576 42294
rect 19524 42230 19576 42236
rect 19524 42084 19576 42090
rect 19524 42026 19576 42032
rect 19432 41812 19484 41818
rect 19432 41754 19484 41760
rect 19536 41721 19564 42026
rect 19522 41712 19578 41721
rect 19522 41647 19578 41656
rect 19432 41540 19484 41546
rect 19432 41482 19484 41488
rect 19340 41472 19392 41478
rect 19340 41414 19392 41420
rect 19248 40588 19300 40594
rect 19248 40530 19300 40536
rect 19444 40526 19472 41482
rect 19628 41414 19656 43166
rect 19708 42016 19760 42022
rect 19708 41958 19760 41964
rect 19720 41818 19748 41958
rect 19708 41812 19760 41818
rect 19708 41754 19760 41760
rect 19706 41576 19762 41585
rect 19812 41562 19840 44463
rect 19892 43308 19944 43314
rect 19892 43250 19944 43256
rect 19904 42090 19932 43250
rect 19984 43240 20036 43246
rect 19984 43182 20036 43188
rect 19892 42084 19944 42090
rect 19892 42026 19944 42032
rect 19762 41534 19840 41562
rect 19706 41511 19762 41520
rect 19628 41386 19748 41414
rect 19720 41138 19748 41386
rect 19798 41304 19854 41313
rect 19798 41239 19800 41248
rect 19852 41239 19854 41248
rect 19800 41210 19852 41216
rect 19708 41132 19760 41138
rect 19708 41074 19760 41080
rect 19892 41132 19944 41138
rect 19892 41074 19944 41080
rect 19708 40656 19760 40662
rect 19708 40598 19760 40604
rect 19432 40520 19484 40526
rect 19432 40462 19484 40468
rect 19616 40384 19668 40390
rect 19616 40326 19668 40332
rect 18752 40284 19060 40293
rect 18752 40282 18758 40284
rect 18814 40282 18838 40284
rect 18894 40282 18918 40284
rect 18974 40282 18998 40284
rect 19054 40282 19060 40284
rect 18814 40230 18816 40282
rect 18996 40230 18998 40282
rect 18752 40228 18758 40230
rect 18814 40228 18838 40230
rect 18894 40228 18918 40230
rect 18974 40228 18998 40230
rect 19054 40228 19060 40230
rect 18752 40219 19060 40228
rect 19628 40186 19656 40326
rect 19616 40180 19668 40186
rect 19616 40122 19668 40128
rect 19432 39908 19484 39914
rect 19432 39850 19484 39856
rect 18752 39196 19060 39205
rect 18752 39194 18758 39196
rect 18814 39194 18838 39196
rect 18894 39194 18918 39196
rect 18974 39194 18998 39196
rect 19054 39194 19060 39196
rect 18814 39142 18816 39194
rect 18996 39142 18998 39194
rect 18752 39140 18758 39142
rect 18814 39140 18838 39142
rect 18894 39140 18918 39142
rect 18974 39140 18998 39142
rect 19054 39140 19060 39142
rect 18752 39131 19060 39140
rect 18604 38752 18656 38758
rect 19444 38729 19472 39850
rect 18604 38694 18656 38700
rect 19430 38720 19486 38729
rect 18616 33538 18644 38694
rect 19430 38655 19486 38664
rect 18752 38108 19060 38117
rect 18752 38106 18758 38108
rect 18814 38106 18838 38108
rect 18894 38106 18918 38108
rect 18974 38106 18998 38108
rect 19054 38106 19060 38108
rect 18814 38054 18816 38106
rect 18996 38054 18998 38106
rect 18752 38052 18758 38054
rect 18814 38052 18838 38054
rect 18894 38052 18918 38054
rect 18974 38052 18998 38054
rect 19054 38052 19060 38054
rect 18752 38043 19060 38052
rect 19524 37800 19576 37806
rect 19524 37742 19576 37748
rect 18752 37020 19060 37029
rect 18752 37018 18758 37020
rect 18814 37018 18838 37020
rect 18894 37018 18918 37020
rect 18974 37018 18998 37020
rect 19054 37018 19060 37020
rect 18814 36966 18816 37018
rect 18996 36966 18998 37018
rect 18752 36964 18758 36966
rect 18814 36964 18838 36966
rect 18894 36964 18918 36966
rect 18974 36964 18998 36966
rect 19054 36964 19060 36966
rect 18752 36955 19060 36964
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 18752 35932 19060 35941
rect 18752 35930 18758 35932
rect 18814 35930 18838 35932
rect 18894 35930 18918 35932
rect 18974 35930 18998 35932
rect 19054 35930 19060 35932
rect 18814 35878 18816 35930
rect 18996 35878 18998 35930
rect 18752 35876 18758 35878
rect 18814 35876 18838 35878
rect 18894 35876 18918 35878
rect 18974 35876 18998 35878
rect 19054 35876 19060 35878
rect 18752 35867 19060 35876
rect 19064 35488 19116 35494
rect 19064 35430 19116 35436
rect 19076 35290 19104 35430
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 19260 35018 19288 36722
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19352 35834 19380 35974
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19248 35012 19300 35018
rect 19248 34954 19300 34960
rect 18752 34844 19060 34853
rect 18752 34842 18758 34844
rect 18814 34842 18838 34844
rect 18894 34842 18918 34844
rect 18974 34842 18998 34844
rect 19054 34842 19060 34844
rect 18814 34790 18816 34842
rect 18996 34790 18998 34842
rect 18752 34788 18758 34790
rect 18814 34788 18838 34790
rect 18894 34788 18918 34790
rect 18974 34788 18998 34790
rect 19054 34788 19060 34790
rect 18752 34779 19060 34788
rect 18972 34604 19024 34610
rect 18972 34546 19024 34552
rect 18984 34513 19012 34546
rect 19064 34536 19116 34542
rect 18970 34504 19026 34513
rect 19064 34478 19116 34484
rect 18970 34439 19026 34448
rect 19076 33844 19104 34478
rect 19076 33816 19196 33844
rect 18752 33756 19060 33765
rect 18752 33754 18758 33756
rect 18814 33754 18838 33756
rect 18894 33754 18918 33756
rect 18974 33754 18998 33756
rect 19054 33754 19060 33756
rect 18814 33702 18816 33754
rect 18996 33702 18998 33754
rect 18752 33700 18758 33702
rect 18814 33700 18838 33702
rect 18894 33700 18918 33702
rect 18974 33700 18998 33702
rect 19054 33700 19060 33702
rect 18752 33691 19060 33700
rect 18972 33584 19024 33590
rect 18970 33552 18972 33561
rect 19024 33552 19026 33561
rect 18616 33510 18736 33538
rect 18604 33448 18656 33454
rect 18604 33390 18656 33396
rect 18432 33102 18552 33130
rect 18616 33114 18644 33390
rect 18604 33108 18656 33114
rect 18432 22137 18460 33102
rect 18604 33050 18656 33056
rect 18708 32994 18736 33510
rect 19168 33522 19196 33816
rect 18970 33487 19026 33496
rect 19156 33516 19208 33522
rect 19156 33458 19208 33464
rect 18524 32966 18736 32994
rect 18524 26874 18552 32966
rect 18752 32668 19060 32677
rect 18752 32666 18758 32668
rect 18814 32666 18838 32668
rect 18894 32666 18918 32668
rect 18974 32666 18998 32668
rect 19054 32666 19060 32668
rect 18814 32614 18816 32666
rect 18996 32614 18998 32666
rect 18752 32612 18758 32614
rect 18814 32612 18838 32614
rect 18894 32612 18918 32614
rect 18974 32612 18998 32614
rect 19054 32612 19060 32614
rect 18752 32603 19060 32612
rect 19168 32434 19196 33458
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19260 32314 19288 34954
rect 19352 34678 19380 35022
rect 19432 35012 19484 35018
rect 19432 34954 19484 34960
rect 19444 34746 19472 34954
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 19340 34672 19392 34678
rect 19340 34614 19392 34620
rect 19536 33930 19564 37742
rect 19616 34944 19668 34950
rect 19616 34886 19668 34892
rect 19628 34678 19656 34886
rect 19616 34672 19668 34678
rect 19616 34614 19668 34620
rect 19524 33924 19576 33930
rect 19524 33866 19576 33872
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19338 33416 19394 33425
rect 19444 33386 19472 33458
rect 19338 33351 19394 33360
rect 19432 33380 19484 33386
rect 19352 32502 19380 33351
rect 19432 33322 19484 33328
rect 19340 32496 19392 32502
rect 19340 32438 19392 32444
rect 19168 32286 19288 32314
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18616 31464 18644 32166
rect 18752 31580 19060 31589
rect 18752 31578 18758 31580
rect 18814 31578 18838 31580
rect 18894 31578 18918 31580
rect 18974 31578 18998 31580
rect 19054 31578 19060 31580
rect 18814 31526 18816 31578
rect 18996 31526 18998 31578
rect 18752 31524 18758 31526
rect 18814 31524 18838 31526
rect 18894 31524 18918 31526
rect 18974 31524 18998 31526
rect 19054 31524 19060 31526
rect 18752 31515 19060 31524
rect 18616 31436 18736 31464
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18616 30938 18644 31078
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 18708 30818 18736 31436
rect 18616 30790 18736 30818
rect 18616 29170 18644 30790
rect 18752 30492 19060 30501
rect 18752 30490 18758 30492
rect 18814 30490 18838 30492
rect 18894 30490 18918 30492
rect 18974 30490 18998 30492
rect 19054 30490 19060 30492
rect 18814 30438 18816 30490
rect 18996 30438 18998 30490
rect 18752 30436 18758 30438
rect 18814 30436 18838 30438
rect 18894 30436 18918 30438
rect 18974 30436 18998 30438
rect 19054 30436 19060 30438
rect 18752 30427 19060 30436
rect 19064 30252 19116 30258
rect 19168 30240 19196 32286
rect 19352 31958 19380 32438
rect 19340 31952 19392 31958
rect 19340 31894 19392 31900
rect 19536 31754 19564 33866
rect 19720 33153 19748 40598
rect 19800 39908 19852 39914
rect 19800 39850 19852 39856
rect 19812 39137 19840 39850
rect 19798 39128 19854 39137
rect 19798 39063 19854 39072
rect 19800 36032 19852 36038
rect 19800 35974 19852 35980
rect 19812 34406 19840 35974
rect 19904 35306 19932 41074
rect 19996 40372 20024 43182
rect 20088 42265 20116 44463
rect 20364 43450 20392 44463
rect 20640 43450 20668 44463
rect 20720 43784 20772 43790
rect 20720 43726 20772 43732
rect 20352 43444 20404 43450
rect 20352 43386 20404 43392
rect 20628 43444 20680 43450
rect 20628 43386 20680 43392
rect 20536 43376 20588 43382
rect 20456 43336 20536 43364
rect 20456 42378 20484 43336
rect 20536 43318 20588 43324
rect 20628 43308 20680 43314
rect 20628 43250 20680 43256
rect 20536 42560 20588 42566
rect 20536 42502 20588 42508
rect 20364 42350 20484 42378
rect 20074 42256 20130 42265
rect 20074 42191 20130 42200
rect 20260 42152 20312 42158
rect 20260 42094 20312 42100
rect 20272 41478 20300 42094
rect 20260 41472 20312 41478
rect 20260 41414 20312 41420
rect 20364 41274 20392 42350
rect 20548 41750 20576 42502
rect 20640 42362 20668 43250
rect 20732 43178 20760 43726
rect 20916 43178 20944 44463
rect 20996 43716 21048 43722
rect 20996 43658 21048 43664
rect 20720 43172 20772 43178
rect 20720 43114 20772 43120
rect 20904 43172 20956 43178
rect 20904 43114 20956 43120
rect 20812 42900 20864 42906
rect 20812 42842 20864 42848
rect 20824 42362 20852 42842
rect 20628 42356 20680 42362
rect 20628 42298 20680 42304
rect 20812 42356 20864 42362
rect 20812 42298 20864 42304
rect 20626 42256 20682 42265
rect 21008 42226 21036 43658
rect 21192 43450 21220 44463
rect 21272 43852 21324 43858
rect 21272 43794 21324 43800
rect 21180 43444 21232 43450
rect 21180 43386 21232 43392
rect 21284 42702 21312 43794
rect 21468 43364 21496 44463
rect 21744 43858 21772 44463
rect 21732 43852 21784 43858
rect 21732 43794 21784 43800
rect 21548 43376 21600 43382
rect 21468 43336 21548 43364
rect 21548 43318 21600 43324
rect 21640 43308 21692 43314
rect 21640 43250 21692 43256
rect 21364 42764 21416 42770
rect 21364 42706 21416 42712
rect 21272 42696 21324 42702
rect 21272 42638 21324 42644
rect 21180 42560 21232 42566
rect 21180 42502 21232 42508
rect 20626 42191 20682 42200
rect 20996 42220 21048 42226
rect 20640 41834 20668 42191
rect 20996 42162 21048 42168
rect 20904 42152 20956 42158
rect 20904 42094 20956 42100
rect 20640 41818 20760 41834
rect 20640 41812 20772 41818
rect 20640 41806 20720 41812
rect 20720 41754 20772 41760
rect 20812 41812 20864 41818
rect 20812 41754 20864 41760
rect 20444 41744 20496 41750
rect 20444 41686 20496 41692
rect 20536 41744 20588 41750
rect 20536 41686 20588 41692
rect 20352 41268 20404 41274
rect 20352 41210 20404 41216
rect 20456 41070 20484 41686
rect 20718 41440 20774 41449
rect 20640 41386 20718 41414
rect 20640 41274 20668 41386
rect 20718 41375 20774 41384
rect 20628 41268 20680 41274
rect 20628 41210 20680 41216
rect 20536 41132 20588 41138
rect 20536 41074 20588 41080
rect 20628 41132 20680 41138
rect 20628 41074 20680 41080
rect 20444 41064 20496 41070
rect 20444 41006 20496 41012
rect 20444 40928 20496 40934
rect 20444 40870 20496 40876
rect 20456 40662 20484 40870
rect 20260 40656 20312 40662
rect 20260 40598 20312 40604
rect 20444 40656 20496 40662
rect 20444 40598 20496 40604
rect 20168 40520 20220 40526
rect 20168 40462 20220 40468
rect 20076 40384 20128 40390
rect 19996 40344 20076 40372
rect 20076 40326 20128 40332
rect 19984 40044 20036 40050
rect 19984 39986 20036 39992
rect 19996 39642 20024 39986
rect 20074 39944 20130 39953
rect 20074 39879 20076 39888
rect 20128 39879 20130 39888
rect 20076 39850 20128 39856
rect 19984 39636 20036 39642
rect 19984 39578 20036 39584
rect 19984 39024 20036 39030
rect 19984 38966 20036 38972
rect 19996 37346 20024 38966
rect 20076 38344 20128 38350
rect 20076 38286 20128 38292
rect 20088 37466 20116 38286
rect 20180 37738 20208 40462
rect 20272 40361 20300 40598
rect 20258 40352 20314 40361
rect 20258 40287 20314 40296
rect 20168 37732 20220 37738
rect 20168 37674 20220 37680
rect 20076 37460 20128 37466
rect 20076 37402 20128 37408
rect 19996 37318 20116 37346
rect 19904 35290 20024 35306
rect 19904 35284 20036 35290
rect 19904 35278 19984 35284
rect 19800 34400 19852 34406
rect 19800 34342 19852 34348
rect 19904 34388 19932 35278
rect 19984 35226 20036 35232
rect 19984 34400 20036 34406
rect 19904 34360 19984 34388
rect 19812 33998 19840 34342
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19904 33862 19932 34360
rect 19984 34342 20036 34348
rect 19892 33856 19944 33862
rect 19892 33798 19944 33804
rect 19706 33144 19762 33153
rect 19706 33079 19762 33088
rect 19708 32836 19760 32842
rect 19708 32778 19760 32784
rect 19720 32434 19748 32778
rect 19708 32428 19760 32434
rect 19708 32370 19760 32376
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19352 31726 19564 31754
rect 19352 31278 19380 31726
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19340 31272 19392 31278
rect 19340 31214 19392 31220
rect 19444 31226 19472 31282
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19260 30394 19288 30534
rect 19248 30388 19300 30394
rect 19248 30330 19300 30336
rect 19116 30212 19196 30240
rect 19064 30194 19116 30200
rect 18752 29404 19060 29413
rect 18752 29402 18758 29404
rect 18814 29402 18838 29404
rect 18894 29402 18918 29404
rect 18974 29402 18998 29404
rect 19054 29402 19060 29404
rect 18814 29350 18816 29402
rect 18996 29350 18998 29402
rect 18752 29348 18758 29350
rect 18814 29348 18838 29350
rect 18894 29348 18918 29350
rect 18974 29348 18998 29350
rect 19054 29348 19060 29350
rect 18752 29339 19060 29348
rect 18604 29164 18656 29170
rect 18604 29106 18656 29112
rect 18604 29028 18656 29034
rect 18604 28970 18656 28976
rect 18616 27062 18644 28970
rect 19156 28552 19208 28558
rect 19156 28494 19208 28500
rect 18752 28316 19060 28325
rect 18752 28314 18758 28316
rect 18814 28314 18838 28316
rect 18894 28314 18918 28316
rect 18974 28314 18998 28316
rect 19054 28314 19060 28316
rect 18814 28262 18816 28314
rect 18996 28262 18998 28314
rect 18752 28260 18758 28262
rect 18814 28260 18838 28262
rect 18894 28260 18918 28262
rect 18974 28260 18998 28262
rect 19054 28260 19060 28262
rect 18752 28251 19060 28260
rect 19168 28218 19196 28494
rect 19156 28212 19208 28218
rect 19156 28154 19208 28160
rect 18752 27228 19060 27237
rect 18752 27226 18758 27228
rect 18814 27226 18838 27228
rect 18894 27226 18918 27228
rect 18974 27226 18998 27228
rect 19054 27226 19060 27228
rect 18814 27174 18816 27226
rect 18996 27174 18998 27226
rect 18752 27172 18758 27174
rect 18814 27172 18838 27174
rect 18894 27172 18918 27174
rect 18974 27172 18998 27174
rect 19054 27172 19060 27174
rect 18752 27163 19060 27172
rect 18604 27056 18656 27062
rect 18604 26998 18656 27004
rect 18524 26846 19196 26874
rect 18694 26480 18750 26489
rect 18694 26415 18696 26424
rect 18748 26415 18750 26424
rect 18696 26386 18748 26392
rect 18752 26140 19060 26149
rect 18752 26138 18758 26140
rect 18814 26138 18838 26140
rect 18894 26138 18918 26140
rect 18974 26138 18998 26140
rect 19054 26138 19060 26140
rect 18814 26086 18816 26138
rect 18996 26086 18998 26138
rect 18752 26084 18758 26086
rect 18814 26084 18838 26086
rect 18894 26084 18918 26086
rect 18974 26084 18998 26086
rect 19054 26084 19060 26086
rect 18752 26075 19060 26084
rect 18696 25968 18748 25974
rect 18616 25928 18696 25956
rect 18512 25356 18564 25362
rect 18512 25298 18564 25304
rect 18524 24614 18552 25298
rect 18616 24886 18644 25928
rect 18696 25910 18748 25916
rect 18752 25052 19060 25061
rect 18752 25050 18758 25052
rect 18814 25050 18838 25052
rect 18894 25050 18918 25052
rect 18974 25050 18998 25052
rect 19054 25050 19060 25052
rect 18814 24998 18816 25050
rect 18996 24998 18998 25050
rect 18752 24996 18758 24998
rect 18814 24996 18838 24998
rect 18894 24996 18918 24998
rect 18974 24996 18998 24998
rect 19054 24996 19060 24998
rect 18752 24987 19060 24996
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18708 24342 18736 24754
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18752 23964 19060 23973
rect 18752 23962 18758 23964
rect 18814 23962 18838 23964
rect 18894 23962 18918 23964
rect 18974 23962 18998 23964
rect 19054 23962 19060 23964
rect 18814 23910 18816 23962
rect 18996 23910 18998 23962
rect 18752 23908 18758 23910
rect 18814 23908 18838 23910
rect 18894 23908 18918 23910
rect 18974 23908 18998 23910
rect 19054 23908 19060 23910
rect 18752 23899 19060 23908
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18524 23118 18552 23666
rect 18512 23112 18564 23118
rect 18512 23054 18564 23060
rect 18752 22876 19060 22885
rect 18752 22874 18758 22876
rect 18814 22874 18838 22876
rect 18894 22874 18918 22876
rect 18974 22874 18998 22876
rect 19054 22874 19060 22876
rect 18814 22822 18816 22874
rect 18996 22822 18998 22874
rect 18752 22820 18758 22822
rect 18814 22820 18838 22822
rect 18894 22820 18918 22822
rect 18974 22820 18998 22822
rect 19054 22820 19060 22822
rect 18752 22811 19060 22820
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18524 22234 18552 22374
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18418 22128 18474 22137
rect 18418 22063 18474 22072
rect 18340 21950 18460 21978
rect 18432 21944 18460 21950
rect 18432 21916 18552 21944
rect 18418 21856 18474 21865
rect 18418 21791 18474 21800
rect 18326 21720 18382 21729
rect 18326 21655 18382 21664
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 17814 18092 18158
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18064 14074 18092 17546
rect 18156 16182 18184 19654
rect 18340 18714 18368 21655
rect 18248 18686 18368 18714
rect 18248 17241 18276 18686
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18290 18368 18566
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18234 17232 18290 17241
rect 18234 17167 18290 17176
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16590 18276 16934
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18144 16176 18196 16182
rect 18144 16118 18196 16124
rect 18156 15502 18184 16118
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 15094 18184 15302
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18052 14068 18104 14074
rect 18104 14028 18184 14056
rect 18052 14010 18104 14016
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17960 9716 18012 9722
rect 17960 9658 18012 9664
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17972 8838 18000 9386
rect 17960 8832 18012 8838
rect 17960 8774 18012 8780
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17788 7002 17816 7754
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17880 6866 17908 8434
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17592 5296 17644 5302
rect 17592 5238 17644 5244
rect 17788 5030 17816 6734
rect 17880 6458 17908 6802
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18064 5250 18092 13126
rect 18156 9654 18184 14028
rect 18248 13258 18276 16526
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18340 13734 18368 15506
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18340 12646 18368 13670
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18340 12306 18368 12582
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 18326 12200 18382 12209
rect 18326 12135 18382 12144
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11801 18276 12038
rect 18340 11830 18368 12135
rect 18328 11824 18380 11830
rect 18234 11792 18290 11801
rect 18328 11766 18380 11772
rect 18234 11727 18290 11736
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18156 8090 18184 8366
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18248 6458 18276 11290
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18340 9586 18368 10610
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18326 8528 18382 8537
rect 18326 8463 18328 8472
rect 18380 8463 18382 8472
rect 18328 8434 18380 8440
rect 18432 8378 18460 21791
rect 18524 21468 18552 21916
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21622 18644 21830
rect 18752 21788 19060 21797
rect 18752 21786 18758 21788
rect 18814 21786 18838 21788
rect 18894 21786 18918 21788
rect 18974 21786 18998 21788
rect 19054 21786 19060 21788
rect 18814 21734 18816 21786
rect 18996 21734 18998 21786
rect 18752 21732 18758 21734
rect 18814 21732 18838 21734
rect 18894 21732 18918 21734
rect 18974 21732 18998 21734
rect 19054 21732 19060 21734
rect 18752 21723 19060 21732
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18524 21440 18644 21468
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18524 15042 18552 20198
rect 18616 15144 18644 21440
rect 19064 21412 19116 21418
rect 19064 21354 19116 21360
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18800 21010 18828 21286
rect 19076 21010 19104 21354
rect 19168 21185 19196 26846
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19260 25294 19288 26182
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19260 24886 19288 25094
rect 19248 24880 19300 24886
rect 19248 24822 19300 24828
rect 19260 24410 19288 24822
rect 19248 24404 19300 24410
rect 19248 24346 19300 24352
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 22098 19288 22374
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19154 21176 19210 21185
rect 19154 21111 19210 21120
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 18752 20700 19060 20709
rect 18752 20698 18758 20700
rect 18814 20698 18838 20700
rect 18894 20698 18918 20700
rect 18974 20698 18998 20700
rect 19054 20698 19060 20700
rect 18814 20646 18816 20698
rect 18996 20646 18998 20698
rect 18752 20644 18758 20646
rect 18814 20644 18838 20646
rect 18894 20644 18918 20646
rect 18974 20644 18998 20646
rect 19054 20644 19060 20646
rect 18752 20635 19060 20644
rect 19168 20602 19196 20878
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19260 19922 19288 22034
rect 19352 21146 19380 31214
rect 19444 31198 19564 31226
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19444 28082 19472 30126
rect 19536 28694 19564 31198
rect 19616 29096 19668 29102
rect 19616 29038 19668 29044
rect 19708 29096 19760 29102
rect 19708 29038 19760 29044
rect 19628 28966 19656 29038
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19524 28688 19576 28694
rect 19524 28630 19576 28636
rect 19536 28218 19564 28630
rect 19628 28558 19656 28902
rect 19720 28762 19748 29038
rect 19708 28756 19760 28762
rect 19708 28698 19760 28704
rect 19616 28552 19668 28558
rect 19616 28494 19668 28500
rect 19524 28212 19576 28218
rect 19524 28154 19576 28160
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19708 28076 19760 28082
rect 19708 28018 19760 28024
rect 19444 27538 19472 28018
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19720 27470 19748 28018
rect 19708 27464 19760 27470
rect 19708 27406 19760 27412
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19444 26382 19472 26726
rect 19524 26512 19576 26518
rect 19524 26454 19576 26460
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19536 25430 19564 26454
rect 19524 25424 19576 25430
rect 19524 25366 19576 25372
rect 19628 24585 19656 26998
rect 19708 25356 19760 25362
rect 19708 25298 19760 25304
rect 19614 24576 19670 24585
rect 19614 24511 19670 24520
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19444 24206 19472 24346
rect 19720 24290 19748 25298
rect 19536 24262 19748 24290
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19536 23730 19564 24262
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 19524 23724 19576 23730
rect 19524 23666 19576 23672
rect 19522 23624 19578 23633
rect 19522 23559 19578 23568
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19444 22778 19472 22986
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19352 20856 19380 21082
rect 19352 20828 19472 20856
rect 19338 20768 19394 20777
rect 19338 20703 19394 20712
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 18752 19612 19060 19621
rect 18752 19610 18758 19612
rect 18814 19610 18838 19612
rect 18894 19610 18918 19612
rect 18974 19610 18998 19612
rect 19054 19610 19060 19612
rect 18814 19558 18816 19610
rect 18996 19558 18998 19610
rect 18752 19556 18758 19558
rect 18814 19556 18838 19558
rect 18894 19556 18918 19558
rect 18974 19556 18998 19558
rect 19054 19556 19060 19558
rect 18752 19547 19060 19556
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19076 18612 19104 19314
rect 19168 18834 19196 19654
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19076 18584 19196 18612
rect 18752 18524 19060 18533
rect 18752 18522 18758 18524
rect 18814 18522 18838 18524
rect 18894 18522 18918 18524
rect 18974 18522 18998 18524
rect 19054 18522 19060 18524
rect 18814 18470 18816 18522
rect 18996 18470 18998 18522
rect 18752 18468 18758 18470
rect 18814 18468 18838 18470
rect 18894 18468 18918 18470
rect 18974 18468 18998 18470
rect 19054 18468 19060 18470
rect 18752 18459 19060 18468
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17678 19012 18022
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18752 17436 19060 17445
rect 18752 17434 18758 17436
rect 18814 17434 18838 17436
rect 18894 17434 18918 17436
rect 18974 17434 18998 17436
rect 19054 17434 19060 17436
rect 18814 17382 18816 17434
rect 18996 17382 18998 17434
rect 18752 17380 18758 17382
rect 18814 17380 18838 17382
rect 18894 17380 18918 17382
rect 18974 17380 18998 17382
rect 19054 17380 19060 17382
rect 18752 17371 19060 17380
rect 19168 17320 19196 18584
rect 19260 18290 19288 19450
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19076 17292 19196 17320
rect 19076 16538 19104 17292
rect 19154 17232 19210 17241
rect 19210 17190 19288 17218
rect 19154 17167 19210 17176
rect 19076 16510 19196 16538
rect 18752 16348 19060 16357
rect 18752 16346 18758 16348
rect 18814 16346 18838 16348
rect 18894 16346 18918 16348
rect 18974 16346 18998 16348
rect 19054 16346 19060 16348
rect 18814 16294 18816 16346
rect 18996 16294 18998 16346
rect 18752 16292 18758 16294
rect 18814 16292 18838 16294
rect 18894 16292 18918 16294
rect 18974 16292 18998 16294
rect 19054 16292 19060 16294
rect 18752 16283 19060 16292
rect 19168 15570 19196 16510
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 18752 15260 19060 15269
rect 18752 15258 18758 15260
rect 18814 15258 18838 15260
rect 18894 15258 18918 15260
rect 18974 15258 18998 15260
rect 19054 15258 19060 15260
rect 18814 15206 18816 15258
rect 18996 15206 18998 15258
rect 18752 15204 18758 15206
rect 18814 15204 18838 15206
rect 18894 15204 18918 15206
rect 18974 15204 18998 15206
rect 19054 15204 19060 15206
rect 18752 15195 19060 15204
rect 18616 15116 18736 15144
rect 18524 15014 18644 15042
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14618 18552 14758
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 13530 18552 14214
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18616 12434 18644 15014
rect 18708 14822 18736 15116
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 18752 14172 19060 14181
rect 18752 14170 18758 14172
rect 18814 14170 18838 14172
rect 18894 14170 18918 14172
rect 18974 14170 18998 14172
rect 19054 14170 19060 14172
rect 18814 14118 18816 14170
rect 18996 14118 18998 14170
rect 18752 14116 18758 14118
rect 18814 14116 18838 14118
rect 18894 14116 18918 14118
rect 18974 14116 18998 14118
rect 19054 14116 19060 14118
rect 18752 14107 19060 14116
rect 19168 14074 19196 14214
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 19076 13734 19104 13874
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 19076 13326 19104 13670
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 18752 13084 19060 13093
rect 18752 13082 18758 13084
rect 18814 13082 18838 13084
rect 18894 13082 18918 13084
rect 18974 13082 18998 13084
rect 19054 13082 19060 13084
rect 18814 13030 18816 13082
rect 18996 13030 18998 13082
rect 18752 13028 18758 13030
rect 18814 13028 18838 13030
rect 18894 13028 18918 13030
rect 18974 13028 18998 13030
rect 19054 13028 19060 13030
rect 18752 13019 19060 13028
rect 19168 12918 19196 13738
rect 19260 13274 19288 17190
rect 19352 16561 19380 20703
rect 19444 20602 19472 20828
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19430 19408 19486 19417
rect 19430 19343 19432 19352
rect 19484 19343 19486 19352
rect 19432 19314 19484 19320
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19444 17338 19472 17546
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19536 17218 19564 23559
rect 19628 23526 19656 24142
rect 19720 23866 19748 24142
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19812 23746 19840 31962
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19892 29776 19944 29782
rect 19892 29718 19944 29724
rect 19904 24614 19932 29718
rect 19996 29510 20024 29990
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19996 28626 20024 29446
rect 20088 29073 20116 37318
rect 20548 37262 20576 41074
rect 20640 39930 20668 41074
rect 20720 41064 20772 41070
rect 20720 41006 20772 41012
rect 20732 40050 20760 41006
rect 20720 40044 20772 40050
rect 20720 39986 20772 39992
rect 20640 39902 20760 39930
rect 20628 38956 20680 38962
rect 20628 38898 20680 38904
rect 20640 38554 20668 38898
rect 20628 38548 20680 38554
rect 20628 38490 20680 38496
rect 20732 38418 20760 39902
rect 20720 38412 20772 38418
rect 20720 38354 20772 38360
rect 20260 37256 20312 37262
rect 20260 37198 20312 37204
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20272 36786 20300 37198
rect 20732 36922 20760 37198
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20260 36780 20312 36786
rect 20260 36722 20312 36728
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20720 36780 20772 36786
rect 20720 36722 20772 36728
rect 20272 36310 20300 36722
rect 20260 36304 20312 36310
rect 20260 36246 20312 36252
rect 20548 36242 20576 36722
rect 20732 36582 20760 36722
rect 20720 36576 20772 36582
rect 20720 36518 20772 36524
rect 20824 36394 20852 41754
rect 20916 41414 20944 42094
rect 20996 42084 21048 42090
rect 20996 42026 21048 42032
rect 21008 41585 21036 42026
rect 21088 41812 21140 41818
rect 21088 41754 21140 41760
rect 20994 41576 21050 41585
rect 20994 41511 21050 41520
rect 20916 41386 21036 41414
rect 20902 41032 20958 41041
rect 20902 40967 20958 40976
rect 20916 40050 20944 40967
rect 20904 40044 20956 40050
rect 20904 39986 20956 39992
rect 20904 39840 20956 39846
rect 20904 39782 20956 39788
rect 20916 39522 20944 39782
rect 21008 39642 21036 41386
rect 21100 40730 21128 41754
rect 21192 41274 21220 42502
rect 21272 42220 21324 42226
rect 21272 42162 21324 42168
rect 21284 41274 21312 42162
rect 21180 41268 21232 41274
rect 21180 41210 21232 41216
rect 21272 41268 21324 41274
rect 21272 41210 21324 41216
rect 21180 41132 21232 41138
rect 21180 41074 21232 41080
rect 21272 41132 21324 41138
rect 21272 41074 21324 41080
rect 21088 40724 21140 40730
rect 21088 40666 21140 40672
rect 21088 40520 21140 40526
rect 21088 40462 21140 40468
rect 21100 39642 21128 40462
rect 20996 39636 21048 39642
rect 20996 39578 21048 39584
rect 21088 39636 21140 39642
rect 21088 39578 21140 39584
rect 20916 39494 21036 39522
rect 20904 39432 20956 39438
rect 20904 39374 20956 39380
rect 20916 39098 20944 39374
rect 20904 39092 20956 39098
rect 20904 39034 20956 39040
rect 21008 38962 21036 39494
rect 21088 39432 21140 39438
rect 21086 39400 21088 39409
rect 21140 39400 21142 39409
rect 21086 39335 21142 39344
rect 20996 38956 21048 38962
rect 20996 38898 21048 38904
rect 21192 38554 21220 41074
rect 21284 40730 21312 41074
rect 21272 40724 21324 40730
rect 21272 40666 21324 40672
rect 21376 40610 21404 42706
rect 21548 42628 21600 42634
rect 21548 42570 21600 42576
rect 21456 41472 21508 41478
rect 21456 41414 21508 41420
rect 21560 41414 21588 42570
rect 21652 42362 21680 43250
rect 22020 43194 22048 44463
rect 22192 43240 22244 43246
rect 22020 43166 22140 43194
rect 22192 43182 22244 43188
rect 21719 43004 22027 43013
rect 21719 43002 21725 43004
rect 21781 43002 21805 43004
rect 21861 43002 21885 43004
rect 21941 43002 21965 43004
rect 22021 43002 22027 43004
rect 21781 42950 21783 43002
rect 21963 42950 21965 43002
rect 21719 42948 21725 42950
rect 21781 42948 21805 42950
rect 21861 42948 21885 42950
rect 21941 42948 21965 42950
rect 22021 42948 22027 42950
rect 21719 42939 22027 42948
rect 22112 42786 22140 43166
rect 21928 42758 22140 42786
rect 21928 42702 21956 42758
rect 21916 42696 21968 42702
rect 21916 42638 21968 42644
rect 21640 42356 21692 42362
rect 21640 42298 21692 42304
rect 21719 41916 22027 41925
rect 21719 41914 21725 41916
rect 21781 41914 21805 41916
rect 21861 41914 21885 41916
rect 21941 41914 21965 41916
rect 22021 41914 22027 41916
rect 21781 41862 21783 41914
rect 21963 41862 21965 41914
rect 21719 41860 21725 41862
rect 21781 41860 21805 41862
rect 21861 41860 21885 41862
rect 21941 41860 21965 41862
rect 22021 41860 22027 41862
rect 21719 41851 22027 41860
rect 21640 41744 21692 41750
rect 21640 41686 21692 41692
rect 21824 41744 21876 41750
rect 21824 41686 21876 41692
rect 21652 41614 21680 41686
rect 21640 41608 21692 41614
rect 21640 41550 21692 41556
rect 21836 41449 21864 41686
rect 22008 41472 22060 41478
rect 21822 41440 21878 41449
rect 21468 41290 21496 41414
rect 21560 41386 21772 41414
rect 21468 41262 21588 41290
rect 21454 41032 21510 41041
rect 21454 40967 21510 40976
rect 21468 40934 21496 40967
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 21284 40582 21404 40610
rect 21284 40390 21312 40582
rect 21456 40520 21508 40526
rect 21456 40462 21508 40468
rect 21272 40384 21324 40390
rect 21272 40326 21324 40332
rect 21272 40044 21324 40050
rect 21272 39986 21324 39992
rect 21364 40044 21416 40050
rect 21364 39986 21416 39992
rect 21284 39846 21312 39986
rect 21272 39840 21324 39846
rect 21272 39782 21324 39788
rect 21272 39432 21324 39438
rect 21272 39374 21324 39380
rect 21284 39098 21312 39374
rect 21376 39273 21404 39986
rect 21362 39264 21418 39273
rect 21362 39199 21418 39208
rect 21272 39092 21324 39098
rect 21272 39034 21324 39040
rect 21364 39092 21416 39098
rect 21364 39034 21416 39040
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 21088 36576 21140 36582
rect 21088 36518 21140 36524
rect 20732 36366 20852 36394
rect 21100 36378 21128 36518
rect 21088 36372 21140 36378
rect 20536 36236 20588 36242
rect 20536 36178 20588 36184
rect 20628 35216 20680 35222
rect 20628 35158 20680 35164
rect 20640 35018 20668 35158
rect 20628 35012 20680 35018
rect 20628 34954 20680 34960
rect 20444 34672 20496 34678
rect 20732 34649 20760 36366
rect 21088 36314 21140 36320
rect 20812 36304 20864 36310
rect 20812 36246 20864 36252
rect 20824 35850 20852 36246
rect 20824 35822 21128 35850
rect 20994 35728 21050 35737
rect 20994 35663 21050 35672
rect 20444 34614 20496 34620
rect 20718 34640 20774 34649
rect 20456 34406 20484 34614
rect 20718 34575 20774 34584
rect 20444 34400 20496 34406
rect 20444 34342 20496 34348
rect 20812 34400 20864 34406
rect 20812 34342 20864 34348
rect 20824 34202 20852 34342
rect 20536 34196 20588 34202
rect 20812 34196 20864 34202
rect 20588 34156 20668 34184
rect 20536 34138 20588 34144
rect 20536 32224 20588 32230
rect 20536 32166 20588 32172
rect 20548 32026 20576 32166
rect 20640 32042 20668 34156
rect 20812 34138 20864 34144
rect 21008 34082 21036 35663
rect 21100 35034 21128 35822
rect 21272 35692 21324 35698
rect 21272 35634 21324 35640
rect 21180 35488 21232 35494
rect 21180 35430 21232 35436
rect 21192 35154 21220 35430
rect 21180 35148 21232 35154
rect 21180 35090 21232 35096
rect 21284 35057 21312 35634
rect 21270 35048 21326 35057
rect 21100 35006 21220 35034
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21100 34202 21128 34478
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 21008 34054 21128 34082
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21008 33318 21036 33458
rect 20996 33312 21048 33318
rect 20996 33254 21048 33260
rect 20536 32020 20588 32026
rect 20536 31962 20588 31968
rect 20640 32014 20944 32042
rect 20640 31754 20668 32014
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 20456 31726 20668 31754
rect 20732 31754 20760 31894
rect 20916 31822 20944 32014
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 21100 31754 21128 34054
rect 20732 31726 20852 31754
rect 20074 29064 20130 29073
rect 20074 28999 20130 29008
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20364 28762 20392 28902
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20456 28642 20484 31726
rect 20628 31204 20680 31210
rect 20628 31146 20680 31152
rect 20640 30938 20668 31146
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20824 30734 20852 31726
rect 21008 31726 21128 31754
rect 21008 31634 21036 31726
rect 20916 31606 21036 31634
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20536 30252 20588 30258
rect 20536 30194 20588 30200
rect 20548 29850 20576 30194
rect 20536 29844 20588 29850
rect 20536 29786 20588 29792
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 19984 28620 20036 28626
rect 19984 28562 20036 28568
rect 20364 28614 20484 28642
rect 19996 26926 20024 28562
rect 20364 28558 20392 28614
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20444 28484 20496 28490
rect 20444 28426 20496 28432
rect 20074 27024 20130 27033
rect 20130 26982 20208 27010
rect 20074 26959 20130 26968
rect 19984 26920 20036 26926
rect 19984 26862 20036 26868
rect 19996 26042 20024 26862
rect 19984 26036 20036 26042
rect 19984 25978 20036 25984
rect 19996 25362 20024 25978
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 20088 25498 20116 25638
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19892 24608 19944 24614
rect 19892 24550 19944 24556
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19720 23718 19840 23746
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19628 23118 19656 23462
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19720 22012 19748 23718
rect 19904 23322 19932 24006
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19996 23118 20024 24754
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19700 21984 19748 22012
rect 19616 21956 19668 21962
rect 19616 21898 19668 21904
rect 19628 21622 19656 21898
rect 19700 21876 19728 21984
rect 19700 21848 19748 21876
rect 19616 21616 19668 21622
rect 19616 21558 19668 21564
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19628 21146 19656 21286
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 19444 17190 19564 17218
rect 19338 16552 19394 16561
rect 19338 16487 19394 16496
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19352 15706 19380 16050
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 15026 19380 15370
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19260 13246 19380 13274
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19352 12594 19380 13246
rect 18340 8350 18460 8378
rect 18524 12406 18644 12434
rect 19168 12566 19380 12594
rect 19168 12434 19196 12566
rect 19444 12434 19472 17190
rect 19628 16658 19656 20538
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19536 15026 19564 15846
rect 19628 15502 19656 16594
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19616 15088 19668 15094
rect 19616 15030 19668 15036
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19628 14074 19656 15030
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13394 19564 13670
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19168 12406 19288 12434
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5370 18184 6122
rect 18248 5914 18276 6258
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18248 5370 18276 5850
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18340 5250 18368 8350
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18432 7546 18460 8230
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18432 5370 18460 6190
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 17960 5228 18012 5234
rect 18064 5222 18184 5250
rect 17960 5170 18012 5176
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17880 4146 17908 4490
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17972 4078 18000 5170
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17682 3904 17738 3913
rect 17682 3839 17738 3848
rect 17958 3904 18014 3913
rect 17958 3839 18014 3848
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 16580 1896 16632 1902
rect 16580 1838 16632 1844
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 16580 1488 16632 1494
rect 16580 1430 16632 1436
rect 16488 1352 16540 1358
rect 16488 1294 16540 1300
rect 16592 1204 16620 1430
rect 16672 1420 16724 1426
rect 16672 1362 16724 1368
rect 15948 598 16436 626
rect 16500 1176 16620 1204
rect 15948 160 15976 598
rect 16500 490 16528 1176
rect 16408 462 16528 490
rect 14554 54 14780 82
rect 14554 0 14610 54
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 82 16266 160
rect 16408 82 16436 462
rect 16684 218 16712 1362
rect 16500 190 16712 218
rect 16500 160 16528 190
rect 16210 54 16436 82
rect 16210 0 16266 54
rect 16486 0 16542 160
rect 16762 82 16818 160
rect 16868 82 16896 1702
rect 17052 1358 17080 2246
rect 17040 1352 17092 1358
rect 17040 1294 17092 1300
rect 17144 1170 17172 2246
rect 17236 1358 17264 2790
rect 17420 1850 17448 3334
rect 17590 3088 17646 3097
rect 17696 3058 17724 3839
rect 17972 3534 18000 3839
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 17590 3023 17592 3032
rect 17644 3023 17646 3032
rect 17684 3052 17736 3058
rect 17592 2994 17644 3000
rect 17788 3040 17816 3334
rect 17788 3012 17908 3040
rect 17684 2994 17736 3000
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17512 2038 17540 2790
rect 17684 2440 17736 2446
rect 17682 2408 17684 2417
rect 17736 2408 17738 2417
rect 17592 2372 17644 2378
rect 17682 2343 17738 2352
rect 17592 2314 17644 2320
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17604 1850 17632 2314
rect 17788 2106 17816 2790
rect 17880 2446 17908 3012
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17776 2100 17828 2106
rect 17776 2042 17828 2048
rect 17420 1822 17540 1850
rect 17604 1822 17724 1850
rect 17408 1760 17460 1766
rect 17408 1702 17460 1708
rect 17224 1352 17276 1358
rect 17224 1294 17276 1300
rect 17052 1142 17172 1170
rect 17052 160 17080 1142
rect 16762 54 16896 82
rect 16762 0 16818 54
rect 17038 0 17094 160
rect 17314 82 17370 160
rect 17420 82 17448 1702
rect 17512 1358 17540 1822
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17500 1352 17552 1358
rect 17500 1294 17552 1300
rect 17604 160 17632 1702
rect 17696 1290 17724 1822
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 17972 1408 18000 1498
rect 17880 1380 18000 1408
rect 17684 1284 17736 1290
rect 17684 1226 17736 1232
rect 17880 160 17908 1380
rect 18064 1018 18092 3334
rect 18156 1834 18184 5222
rect 18248 5222 18368 5250
rect 18248 3126 18276 5222
rect 18524 4604 18552 12406
rect 19154 12336 19210 12345
rect 18604 12300 18656 12306
rect 19154 12271 19210 12280
rect 18604 12242 18656 12248
rect 18616 11830 18644 12242
rect 18752 11996 19060 12005
rect 18752 11994 18758 11996
rect 18814 11994 18838 11996
rect 18894 11994 18918 11996
rect 18974 11994 18998 11996
rect 19054 11994 19060 11996
rect 18814 11942 18816 11994
rect 18996 11942 18998 11994
rect 18752 11940 18758 11942
rect 18814 11940 18838 11942
rect 18894 11940 18918 11942
rect 18974 11940 18998 11942
rect 19054 11940 19060 11942
rect 18752 11931 19060 11940
rect 18604 11824 18656 11830
rect 18604 11766 18656 11772
rect 18616 11354 18644 11766
rect 19168 11626 19196 12271
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11354 19104 11494
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 10266 18644 11086
rect 18752 10908 19060 10917
rect 18752 10906 18758 10908
rect 18814 10906 18838 10908
rect 18894 10906 18918 10908
rect 18974 10906 18998 10908
rect 19054 10906 19060 10908
rect 18814 10854 18816 10906
rect 18996 10854 18998 10906
rect 18752 10852 18758 10854
rect 18814 10852 18838 10854
rect 18894 10852 18918 10854
rect 18974 10852 18998 10854
rect 19054 10852 19060 10854
rect 18752 10843 19060 10852
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19168 10266 19196 10406
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 18752 9820 19060 9829
rect 18752 9818 18758 9820
rect 18814 9818 18838 9820
rect 18894 9818 18918 9820
rect 18974 9818 18998 9820
rect 19054 9818 19060 9820
rect 18814 9766 18816 9818
rect 18996 9766 18998 9818
rect 18752 9764 18758 9766
rect 18814 9764 18838 9766
rect 18894 9764 18918 9766
rect 18974 9764 18998 9766
rect 19054 9764 19060 9766
rect 18752 9755 19060 9764
rect 19156 8968 19208 8974
rect 19156 8910 19208 8916
rect 18752 8732 19060 8741
rect 18752 8730 18758 8732
rect 18814 8730 18838 8732
rect 18894 8730 18918 8732
rect 18974 8730 18998 8732
rect 19054 8730 19060 8732
rect 18814 8678 18816 8730
rect 18996 8678 18998 8730
rect 18752 8676 18758 8678
rect 18814 8676 18838 8678
rect 18894 8676 18918 8678
rect 18974 8676 18998 8678
rect 19054 8676 19060 8678
rect 18752 8667 19060 8676
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18616 8090 18644 8502
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18616 7002 18644 7822
rect 18708 7750 18736 8230
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18752 7644 19060 7653
rect 18752 7642 18758 7644
rect 18814 7642 18838 7644
rect 18894 7642 18918 7644
rect 18974 7642 18998 7644
rect 19054 7642 19060 7644
rect 18814 7590 18816 7642
rect 18996 7590 18998 7642
rect 18752 7588 18758 7590
rect 18814 7588 18838 7590
rect 18894 7588 18918 7590
rect 18974 7588 18998 7590
rect 19054 7588 19060 7590
rect 18752 7579 19060 7588
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18800 6798 18828 7346
rect 18788 6792 18840 6798
rect 19168 6746 19196 8910
rect 18788 6734 18840 6740
rect 18892 6718 19196 6746
rect 18892 6644 18920 6718
rect 18616 6616 18920 6644
rect 19156 6656 19208 6662
rect 18616 4706 18644 6616
rect 19156 6598 19208 6604
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 19076 5778 19104 6394
rect 19168 5914 19196 6598
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 19260 5794 19288 12406
rect 19352 12406 19472 12434
rect 19352 9602 19380 12406
rect 19536 11218 19564 13194
rect 19628 12850 19656 14010
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10062 19472 11086
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19536 10674 19564 10950
rect 19628 10674 19656 12786
rect 19720 11665 19748 21848
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19812 19446 19840 21354
rect 19800 19440 19852 19446
rect 19800 19382 19852 19388
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 15026 19840 15302
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19904 14906 19932 22714
rect 19984 22500 20036 22506
rect 19984 22442 20036 22448
rect 19996 21622 20024 22442
rect 20180 22094 20208 26982
rect 20456 26586 20484 28426
rect 20260 26580 20312 26586
rect 20260 26522 20312 26528
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20088 22066 20208 22094
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19982 21176 20038 21185
rect 19982 21111 20038 21120
rect 19996 19514 20024 21111
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 20088 16017 20116 22066
rect 20272 22030 20300 26522
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20352 22092 20404 22098
rect 20456 22094 20484 24346
rect 20548 23730 20576 28902
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20732 28529 20760 28630
rect 20718 28520 20774 28529
rect 20718 28455 20774 28464
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 20640 27674 20668 27950
rect 20628 27668 20680 27674
rect 20628 27610 20680 27616
rect 20732 27282 20760 28154
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 27470 20852 27814
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20732 27254 20852 27282
rect 20824 27130 20852 27254
rect 20720 27124 20772 27130
rect 20720 27066 20772 27072
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20640 25498 20668 25842
rect 20628 25492 20680 25498
rect 20628 25434 20680 25440
rect 20628 25288 20680 25294
rect 20626 25256 20628 25265
rect 20680 25256 20682 25265
rect 20626 25191 20682 25200
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20640 24070 20668 24550
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20640 22438 20668 23054
rect 20732 23050 20760 27066
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20732 22778 20760 22986
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20916 22114 20944 31606
rect 21088 31204 21140 31210
rect 21088 31146 21140 31152
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 21008 28218 21036 28358
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 20994 22128 21050 22137
rect 20456 22066 20576 22094
rect 20916 22086 20994 22114
rect 20352 22034 20404 22040
rect 20260 22024 20312 22030
rect 20260 21966 20312 21972
rect 20364 21690 20392 22034
rect 20444 21956 20496 21962
rect 20444 21898 20496 21904
rect 20352 21684 20404 21690
rect 20352 21626 20404 21632
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20272 21321 20300 21490
rect 20258 21312 20314 21321
rect 20258 21247 20314 21256
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 17082 20208 20810
rect 20456 20602 20484 21898
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18970 20300 19110
rect 20456 18970 20484 19382
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20352 17128 20404 17134
rect 20180 17054 20300 17082
rect 20352 17070 20404 17076
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16794 20208 16934
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20074 16008 20130 16017
rect 20074 15943 20130 15952
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 19984 15904 20036 15910
rect 20180 15858 20208 15914
rect 19984 15846 20036 15852
rect 19996 15026 20024 15846
rect 20088 15830 20208 15858
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19904 14878 20024 14906
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19798 13560 19854 13569
rect 19798 13495 19854 13504
rect 19706 11656 19762 11665
rect 19706 11591 19762 11600
rect 19812 11082 19840 13495
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19352 9574 19472 9602
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 8498 19380 9454
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19444 7290 19472 9574
rect 19536 9518 19564 10610
rect 19628 9518 19656 10610
rect 19800 9648 19852 9654
rect 19800 9590 19852 9596
rect 19524 9512 19576 9518
rect 19524 9454 19576 9460
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 8498 19564 9318
rect 19628 9042 19656 9454
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19536 7886 19564 8434
rect 19720 8362 19748 9318
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19812 7392 19840 9590
rect 19904 8401 19932 14758
rect 19996 14006 20024 14878
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19996 13462 20024 13806
rect 19984 13456 20036 13462
rect 19984 13398 20036 13404
rect 19982 13288 20038 13297
rect 19982 13223 20038 13232
rect 19996 13190 20024 13223
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 12918 20024 13126
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 20088 12434 20116 15830
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20180 12986 20208 13194
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20088 12406 20208 12434
rect 20180 12238 20208 12406
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20272 11234 20300 17054
rect 20364 15094 20392 17070
rect 20456 16250 20484 17274
rect 20548 17202 20576 22066
rect 20994 22063 21050 22072
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 21078 20760 21898
rect 20824 21690 20852 21966
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20916 21078 20944 21830
rect 21008 21690 21036 21830
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20720 21072 20772 21078
rect 20904 21072 20956 21078
rect 20720 21014 20772 21020
rect 20810 21040 20866 21049
rect 20904 21014 20956 21020
rect 20810 20975 20866 20984
rect 20824 20890 20852 20975
rect 20824 20862 20944 20890
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20824 19854 20852 20742
rect 20916 20058 20944 20862
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 18766 20668 19654
rect 20916 19334 20944 19994
rect 21100 19938 21128 31146
rect 21192 28966 21220 35006
rect 21270 34983 21326 34992
rect 21272 32564 21324 32570
rect 21272 32506 21324 32512
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 21192 25362 21220 27406
rect 21284 27033 21312 32506
rect 21270 27024 21326 27033
rect 21270 26959 21326 26968
rect 21376 26874 21404 39034
rect 21468 39030 21496 40462
rect 21560 39420 21588 41262
rect 21640 40996 21692 41002
rect 21640 40938 21692 40944
rect 21652 40594 21680 40938
rect 21744 40934 21772 41386
rect 22008 41414 22060 41420
rect 21822 41375 21878 41384
rect 22020 41274 22048 41414
rect 22008 41268 22060 41274
rect 22204 41256 22232 43182
rect 22296 42566 22324 44463
rect 22572 43790 22600 44463
rect 22560 43784 22612 43790
rect 22560 43726 22612 43732
rect 22376 43648 22428 43654
rect 22376 43590 22428 43596
rect 22388 42702 22416 43590
rect 22848 43466 22876 44463
rect 22928 43852 22980 43858
rect 22928 43794 22980 43800
rect 22756 43438 22876 43466
rect 22940 43450 22968 43794
rect 23124 43450 23152 44463
rect 22928 43444 22980 43450
rect 22468 43308 22520 43314
rect 22468 43250 22520 43256
rect 22376 42696 22428 42702
rect 22376 42638 22428 42644
rect 22284 42560 22336 42566
rect 22284 42502 22336 42508
rect 22376 42152 22428 42158
rect 22376 42094 22428 42100
rect 22284 42016 22336 42022
rect 22284 41958 22336 41964
rect 22296 41682 22324 41958
rect 22284 41676 22336 41682
rect 22284 41618 22336 41624
rect 22388 41546 22416 42094
rect 22376 41540 22428 41546
rect 22376 41482 22428 41488
rect 22480 41274 22508 43250
rect 22652 43240 22704 43246
rect 22652 43182 22704 43188
rect 22558 41576 22614 41585
rect 22664 41546 22692 43182
rect 22756 42294 22784 43438
rect 22928 43386 22980 43392
rect 23112 43444 23164 43450
rect 23112 43386 23164 43392
rect 23020 43376 23072 43382
rect 23020 43318 23072 43324
rect 23202 43344 23258 43353
rect 22928 43308 22980 43314
rect 22928 43250 22980 43256
rect 22940 43217 22968 43250
rect 22926 43208 22982 43217
rect 22926 43143 22982 43152
rect 22744 42288 22796 42294
rect 22744 42230 22796 42236
rect 22836 42220 22888 42226
rect 22836 42162 22888 42168
rect 22558 41511 22614 41520
rect 22652 41540 22704 41546
rect 22572 41478 22600 41511
rect 22652 41482 22704 41488
rect 22560 41472 22612 41478
rect 22560 41414 22612 41420
rect 22008 41210 22060 41216
rect 22112 41228 22232 41256
rect 22468 41268 22520 41274
rect 21822 41168 21878 41177
rect 21822 41103 21824 41112
rect 21876 41103 21878 41112
rect 21824 41074 21876 41080
rect 22112 40934 22140 41228
rect 22468 41210 22520 41216
rect 22192 41132 22244 41138
rect 22468 41132 22520 41138
rect 22244 41092 22416 41120
rect 22192 41074 22244 41080
rect 22190 41032 22246 41041
rect 22190 40967 22246 40976
rect 21732 40928 21784 40934
rect 21732 40870 21784 40876
rect 22100 40928 22152 40934
rect 22100 40870 22152 40876
rect 21719 40828 22027 40837
rect 21719 40826 21725 40828
rect 21781 40826 21805 40828
rect 21861 40826 21885 40828
rect 21941 40826 21965 40828
rect 22021 40826 22027 40828
rect 21781 40774 21783 40826
rect 21963 40774 21965 40826
rect 21719 40772 21725 40774
rect 21781 40772 21805 40774
rect 21861 40772 21885 40774
rect 21941 40772 21965 40774
rect 22021 40772 22027 40774
rect 21719 40763 22027 40772
rect 22098 40760 22154 40769
rect 21732 40724 21784 40730
rect 22204 40730 22232 40967
rect 22098 40695 22154 40704
rect 22192 40724 22244 40730
rect 21732 40666 21784 40672
rect 21640 40588 21692 40594
rect 21640 40530 21692 40536
rect 21638 40488 21694 40497
rect 21638 40423 21694 40432
rect 21652 40050 21680 40423
rect 21640 40044 21692 40050
rect 21640 39986 21692 39992
rect 21744 39846 21772 40666
rect 22008 40656 22060 40662
rect 22112 40644 22140 40695
rect 22192 40666 22244 40672
rect 22060 40616 22140 40644
rect 22008 40598 22060 40604
rect 22284 40588 22336 40594
rect 22284 40530 22336 40536
rect 22100 40520 22152 40526
rect 22098 40488 22100 40497
rect 22152 40488 22154 40497
rect 22098 40423 22154 40432
rect 21822 40216 21878 40225
rect 21822 40151 21824 40160
rect 21876 40151 21878 40160
rect 21916 40180 21968 40186
rect 21824 40122 21876 40128
rect 22192 40180 22244 40186
rect 21968 40140 22192 40168
rect 21916 40122 21968 40128
rect 22192 40122 22244 40128
rect 21914 40080 21970 40089
rect 21914 40015 21970 40024
rect 22008 40044 22060 40050
rect 21928 39930 21956 40015
rect 22192 40044 22244 40050
rect 22060 40004 22140 40032
rect 22008 39986 22060 39992
rect 21836 39914 21956 39930
rect 21824 39908 21956 39914
rect 21876 39902 21956 39908
rect 21824 39850 21876 39856
rect 21732 39840 21784 39846
rect 21732 39782 21784 39788
rect 21719 39740 22027 39749
rect 21719 39738 21725 39740
rect 21781 39738 21805 39740
rect 21861 39738 21885 39740
rect 21941 39738 21965 39740
rect 22021 39738 22027 39740
rect 21781 39686 21783 39738
rect 21963 39686 21965 39738
rect 21719 39684 21725 39686
rect 21781 39684 21805 39686
rect 21861 39684 21885 39686
rect 21941 39684 21965 39686
rect 22021 39684 22027 39686
rect 21719 39675 22027 39684
rect 21732 39432 21784 39438
rect 21560 39392 21732 39420
rect 21732 39374 21784 39380
rect 22008 39432 22060 39438
rect 22008 39374 22060 39380
rect 22020 39098 22048 39374
rect 22008 39092 22060 39098
rect 22008 39034 22060 39040
rect 21456 39024 21508 39030
rect 21456 38966 21508 38972
rect 21548 38888 21600 38894
rect 22112 38876 22140 40004
rect 22192 39986 22244 39992
rect 22204 39522 22232 39986
rect 22296 39846 22324 40530
rect 22284 39840 22336 39846
rect 22284 39782 22336 39788
rect 22284 39636 22336 39642
rect 22388 39624 22416 41092
rect 22468 41074 22520 41080
rect 22480 41041 22508 41074
rect 22744 41064 22796 41070
rect 22466 41032 22522 41041
rect 22744 41006 22796 41012
rect 22466 40967 22522 40976
rect 22466 40760 22522 40769
rect 22756 40730 22784 41006
rect 22466 40695 22468 40704
rect 22520 40695 22522 40704
rect 22744 40724 22796 40730
rect 22468 40666 22520 40672
rect 22744 40666 22796 40672
rect 22650 40624 22706 40633
rect 22650 40559 22706 40568
rect 22664 40526 22692 40559
rect 22560 40520 22612 40526
rect 22560 40462 22612 40468
rect 22652 40520 22704 40526
rect 22652 40462 22704 40468
rect 22572 39642 22600 40462
rect 22652 40112 22704 40118
rect 22650 40080 22652 40089
rect 22704 40080 22706 40089
rect 22650 40015 22706 40024
rect 22744 40044 22796 40050
rect 22744 39986 22796 39992
rect 22336 39596 22416 39624
rect 22560 39636 22612 39642
rect 22284 39578 22336 39584
rect 22560 39578 22612 39584
rect 22204 39494 22416 39522
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 22112 38848 22232 38876
rect 21548 38830 21600 38836
rect 21560 33454 21588 38830
rect 22204 38758 22232 38848
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 22192 38752 22244 38758
rect 22192 38694 22244 38700
rect 21719 38652 22027 38661
rect 21719 38650 21725 38652
rect 21781 38650 21805 38652
rect 21861 38650 21885 38652
rect 21941 38650 21965 38652
rect 22021 38650 22027 38652
rect 21781 38598 21783 38650
rect 21963 38598 21965 38650
rect 21719 38596 21725 38598
rect 21781 38596 21805 38598
rect 21861 38596 21885 38598
rect 21941 38596 21965 38598
rect 22021 38596 22027 38598
rect 21719 38587 22027 38596
rect 22112 38350 22140 38694
rect 22100 38344 22152 38350
rect 22100 38286 22152 38292
rect 22192 38208 22244 38214
rect 22192 38150 22244 38156
rect 22204 38010 22232 38150
rect 22100 38004 22152 38010
rect 22100 37946 22152 37952
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 22112 37890 22140 37946
rect 22296 37890 22324 39374
rect 22112 37862 22324 37890
rect 21719 37564 22027 37573
rect 21719 37562 21725 37564
rect 21781 37562 21805 37564
rect 21861 37562 21885 37564
rect 21941 37562 21965 37564
rect 22021 37562 22027 37564
rect 21781 37510 21783 37562
rect 21963 37510 21965 37562
rect 21719 37508 21725 37510
rect 21781 37508 21805 37510
rect 21861 37508 21885 37510
rect 21941 37508 21965 37510
rect 22021 37508 22027 37510
rect 21719 37499 22027 37508
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 21836 36922 21864 37198
rect 21916 37188 21968 37194
rect 21916 37130 21968 37136
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 21928 36922 21956 37130
rect 21824 36916 21876 36922
rect 21824 36858 21876 36864
rect 21916 36916 21968 36922
rect 21916 36858 21968 36864
rect 21719 36476 22027 36485
rect 21719 36474 21725 36476
rect 21781 36474 21805 36476
rect 21861 36474 21885 36476
rect 21941 36474 21965 36476
rect 22021 36474 22027 36476
rect 21781 36422 21783 36474
rect 21963 36422 21965 36474
rect 21719 36420 21725 36422
rect 21781 36420 21805 36422
rect 21861 36420 21885 36422
rect 21941 36420 21965 36422
rect 22021 36420 22027 36422
rect 21719 36411 22027 36420
rect 21719 35388 22027 35397
rect 21719 35386 21725 35388
rect 21781 35386 21805 35388
rect 21861 35386 21885 35388
rect 21941 35386 21965 35388
rect 22021 35386 22027 35388
rect 21781 35334 21783 35386
rect 21963 35334 21965 35386
rect 21719 35332 21725 35334
rect 21781 35332 21805 35334
rect 21861 35332 21885 35334
rect 21941 35332 21965 35334
rect 22021 35332 22027 35334
rect 21719 35323 22027 35332
rect 22204 34610 22232 37130
rect 22388 36802 22416 39494
rect 22560 39432 22612 39438
rect 22560 39374 22612 39380
rect 22468 37936 22520 37942
rect 22468 37878 22520 37884
rect 22296 36774 22416 36802
rect 22296 35290 22324 36774
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22388 36378 22416 36654
rect 22376 36372 22428 36378
rect 22376 36314 22428 36320
rect 22376 35624 22428 35630
rect 22376 35566 22428 35572
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22284 35148 22336 35154
rect 22284 35090 22336 35096
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 21719 34300 22027 34309
rect 21719 34298 21725 34300
rect 21781 34298 21805 34300
rect 21861 34298 21885 34300
rect 21941 34298 21965 34300
rect 22021 34298 22027 34300
rect 21781 34246 21783 34298
rect 21963 34246 21965 34298
rect 21719 34244 21725 34246
rect 21781 34244 21805 34246
rect 21861 34244 21885 34246
rect 21941 34244 21965 34246
rect 22021 34244 22027 34246
rect 21719 34235 22027 34244
rect 21640 33856 21692 33862
rect 21640 33798 21692 33804
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21548 31748 21600 31754
rect 21548 31690 21600 31696
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21468 30938 21496 31282
rect 21560 31278 21588 31690
rect 21548 31272 21600 31278
rect 21548 31214 21600 31220
rect 21456 30932 21508 30938
rect 21456 30874 21508 30880
rect 21456 28212 21508 28218
rect 21456 28154 21508 28160
rect 21468 27674 21496 28154
rect 21548 27940 21600 27946
rect 21548 27882 21600 27888
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21560 27402 21588 27882
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21284 26846 21404 26874
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21180 25356 21232 25362
rect 21180 25298 21232 25304
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 21192 20874 21220 25094
rect 21284 21690 21312 26846
rect 21560 26024 21588 26862
rect 21652 26217 21680 33798
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 21719 33212 22027 33221
rect 21719 33210 21725 33212
rect 21781 33210 21805 33212
rect 21861 33210 21885 33212
rect 21941 33210 21965 33212
rect 22021 33210 22027 33212
rect 21781 33158 21783 33210
rect 21963 33158 21965 33210
rect 21719 33156 21725 33158
rect 21781 33156 21805 33158
rect 21861 33156 21885 33158
rect 21941 33156 21965 33158
rect 22021 33156 22027 33158
rect 21719 33147 22027 33156
rect 22204 32910 22232 33254
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 21719 32124 22027 32133
rect 21719 32122 21725 32124
rect 21781 32122 21805 32124
rect 21861 32122 21885 32124
rect 21941 32122 21965 32124
rect 22021 32122 22027 32124
rect 21781 32070 21783 32122
rect 21963 32070 21965 32122
rect 21719 32068 21725 32070
rect 21781 32068 21805 32070
rect 21861 32068 21885 32070
rect 21941 32068 21965 32070
rect 22021 32068 22027 32070
rect 21719 32059 22027 32068
rect 22192 31748 22244 31754
rect 22192 31690 22244 31696
rect 22100 31680 22152 31686
rect 22100 31622 22152 31628
rect 22112 31278 22140 31622
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21719 31036 22027 31045
rect 21719 31034 21725 31036
rect 21781 31034 21805 31036
rect 21861 31034 21885 31036
rect 21941 31034 21965 31036
rect 22021 31034 22027 31036
rect 21781 30982 21783 31034
rect 21963 30982 21965 31034
rect 21719 30980 21725 30982
rect 21781 30980 21805 30982
rect 21861 30980 21885 30982
rect 21941 30980 21965 30982
rect 22021 30980 22027 30982
rect 21719 30971 22027 30980
rect 22112 30258 22140 31214
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 21719 29948 22027 29957
rect 21719 29946 21725 29948
rect 21781 29946 21805 29948
rect 21861 29946 21885 29948
rect 21941 29946 21965 29948
rect 22021 29946 22027 29948
rect 21781 29894 21783 29946
rect 21963 29894 21965 29946
rect 21719 29892 21725 29894
rect 21781 29892 21805 29894
rect 21861 29892 21885 29894
rect 21941 29892 21965 29894
rect 22021 29892 22027 29894
rect 21719 29883 22027 29892
rect 22098 29744 22154 29753
rect 22098 29679 22154 29688
rect 21719 28860 22027 28869
rect 21719 28858 21725 28860
rect 21781 28858 21805 28860
rect 21861 28858 21885 28860
rect 21941 28858 21965 28860
rect 22021 28858 22027 28860
rect 21781 28806 21783 28858
rect 21963 28806 21965 28858
rect 21719 28804 21725 28806
rect 21781 28804 21805 28806
rect 21861 28804 21885 28806
rect 21941 28804 21965 28806
rect 22021 28804 22027 28806
rect 21719 28795 22027 28804
rect 21719 27772 22027 27781
rect 21719 27770 21725 27772
rect 21781 27770 21805 27772
rect 21861 27770 21885 27772
rect 21941 27770 21965 27772
rect 22021 27770 22027 27772
rect 21781 27718 21783 27770
rect 21963 27718 21965 27770
rect 21719 27716 21725 27718
rect 21781 27716 21805 27718
rect 21861 27716 21885 27718
rect 21941 27716 21965 27718
rect 22021 27716 22027 27718
rect 21719 27707 22027 27716
rect 22112 26874 22140 29679
rect 22204 26994 22232 31690
rect 22296 30954 22324 35090
rect 22388 31754 22416 35566
rect 22480 34762 22508 37878
rect 22572 37670 22600 39374
rect 22652 38344 22704 38350
rect 22652 38286 22704 38292
rect 22560 37664 22612 37670
rect 22560 37606 22612 37612
rect 22664 37466 22692 38286
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 22756 37346 22784 39986
rect 22848 39914 22876 42162
rect 22928 41812 22980 41818
rect 22928 41754 22980 41760
rect 22940 41546 22968 41754
rect 22928 41540 22980 41546
rect 22928 41482 22980 41488
rect 22926 41304 22982 41313
rect 22926 41239 22982 41248
rect 22940 40526 22968 41239
rect 23032 40730 23060 43318
rect 23202 43279 23258 43288
rect 23216 42362 23244 43279
rect 23204 42356 23256 42362
rect 23204 42298 23256 42304
rect 23202 41440 23258 41449
rect 23202 41375 23258 41384
rect 23112 41132 23164 41138
rect 23112 41074 23164 41080
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 23020 40452 23072 40458
rect 23020 40394 23072 40400
rect 22928 40384 22980 40390
rect 22928 40326 22980 40332
rect 22836 39908 22888 39914
rect 22836 39850 22888 39856
rect 22940 39846 22968 40326
rect 22928 39840 22980 39846
rect 22928 39782 22980 39788
rect 23032 39137 23060 40394
rect 23124 40089 23152 41074
rect 23110 40080 23166 40089
rect 23110 40015 23166 40024
rect 23112 39296 23164 39302
rect 23110 39264 23112 39273
rect 23164 39264 23166 39273
rect 23110 39199 23166 39208
rect 23018 39128 23074 39137
rect 23018 39063 23074 39072
rect 23216 38570 23244 41375
rect 23400 41274 23428 44463
rect 23676 43058 23704 44463
rect 23492 43030 23704 43058
rect 23492 42022 23520 43030
rect 23952 42786 23980 44463
rect 24124 43104 24176 43110
rect 24124 43046 24176 43052
rect 23676 42758 23980 42786
rect 23572 42084 23624 42090
rect 23572 42026 23624 42032
rect 23480 42016 23532 42022
rect 23480 41958 23532 41964
rect 23388 41268 23440 41274
rect 23388 41210 23440 41216
rect 23480 41200 23532 41206
rect 23480 41142 23532 41148
rect 23296 41064 23348 41070
rect 23296 41006 23348 41012
rect 23308 40526 23336 41006
rect 23492 40594 23520 41142
rect 23480 40588 23532 40594
rect 23480 40530 23532 40536
rect 23296 40520 23348 40526
rect 23296 40462 23348 40468
rect 23478 40488 23534 40497
rect 23478 40423 23534 40432
rect 23492 40390 23520 40423
rect 23480 40384 23532 40390
rect 23480 40326 23532 40332
rect 23386 39536 23442 39545
rect 23386 39471 23442 39480
rect 23400 39438 23428 39471
rect 23388 39432 23440 39438
rect 23388 39374 23440 39380
rect 23584 39080 23612 42026
rect 23676 41818 23704 42758
rect 23756 42628 23808 42634
rect 23756 42570 23808 42576
rect 23768 41970 23796 42570
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 23768 41942 23980 41970
rect 23664 41812 23716 41818
rect 23664 41754 23716 41760
rect 23848 41540 23900 41546
rect 23848 41482 23900 41488
rect 23664 40928 23716 40934
rect 23662 40896 23664 40905
rect 23716 40896 23718 40905
rect 23662 40831 23718 40840
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23676 40361 23704 40462
rect 23662 40352 23718 40361
rect 23662 40287 23718 40296
rect 23860 40186 23888 41482
rect 23952 40225 23980 41942
rect 24044 40730 24072 42162
rect 24136 41993 24164 43046
rect 24228 42702 24256 44463
rect 24216 42696 24268 42702
rect 24216 42638 24268 42644
rect 24504 42362 24532 44463
rect 24780 43738 24808 44463
rect 24596 43710 24808 43738
rect 24596 42702 24624 43710
rect 24686 43548 24994 43557
rect 24686 43546 24692 43548
rect 24748 43546 24772 43548
rect 24828 43546 24852 43548
rect 24908 43546 24932 43548
rect 24988 43546 24994 43548
rect 24748 43494 24750 43546
rect 24930 43494 24932 43546
rect 24686 43492 24692 43494
rect 24748 43492 24772 43494
rect 24828 43492 24852 43494
rect 24908 43492 24932 43494
rect 24988 43492 24994 43494
rect 24686 43483 24994 43492
rect 24584 42696 24636 42702
rect 24584 42638 24636 42644
rect 24686 42460 24994 42469
rect 24686 42458 24692 42460
rect 24748 42458 24772 42460
rect 24828 42458 24852 42460
rect 24908 42458 24932 42460
rect 24988 42458 24994 42460
rect 24748 42406 24750 42458
rect 24930 42406 24932 42458
rect 24686 42404 24692 42406
rect 24748 42404 24772 42406
rect 24828 42404 24852 42406
rect 24908 42404 24932 42406
rect 24988 42404 24994 42406
rect 24686 42395 24994 42404
rect 24492 42356 24544 42362
rect 24492 42298 24544 42304
rect 24584 42152 24636 42158
rect 24584 42094 24636 42100
rect 24216 42084 24268 42090
rect 24216 42026 24268 42032
rect 24122 41984 24178 41993
rect 24122 41919 24178 41928
rect 24032 40724 24084 40730
rect 24032 40666 24084 40672
rect 23938 40216 23994 40225
rect 23848 40180 23900 40186
rect 23938 40151 23994 40160
rect 23848 40122 23900 40128
rect 23756 40044 23808 40050
rect 23756 39986 23808 39992
rect 24124 40044 24176 40050
rect 24124 39986 24176 39992
rect 23492 39052 23612 39080
rect 23296 38752 23348 38758
rect 23296 38694 23348 38700
rect 23032 38542 23244 38570
rect 22836 38208 22888 38214
rect 22836 38150 22888 38156
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 22848 37738 22876 38150
rect 22940 38010 22968 38150
rect 22928 38004 22980 38010
rect 22928 37946 22980 37952
rect 22836 37732 22888 37738
rect 22836 37674 22888 37680
rect 22928 37664 22980 37670
rect 22928 37606 22980 37612
rect 22664 37318 22784 37346
rect 22664 35154 22692 37318
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22756 36009 22784 37198
rect 22940 37126 22968 37606
rect 22928 37120 22980 37126
rect 22928 37062 22980 37068
rect 23032 36904 23060 38542
rect 23112 38412 23164 38418
rect 23112 38354 23164 38360
rect 23124 38010 23152 38354
rect 23308 38350 23336 38694
rect 23204 38344 23256 38350
rect 23204 38286 23256 38292
rect 23296 38344 23348 38350
rect 23296 38286 23348 38292
rect 23112 38004 23164 38010
rect 23112 37946 23164 37952
rect 23216 37398 23244 38286
rect 23388 38276 23440 38282
rect 23388 38218 23440 38224
rect 23400 37466 23428 38218
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 23204 37392 23256 37398
rect 23204 37334 23256 37340
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 22940 36876 23060 36904
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 22848 36378 22876 36518
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22742 36000 22798 36009
rect 22742 35935 22798 35944
rect 22940 35714 22968 36876
rect 23124 36854 23152 37198
rect 23112 36848 23164 36854
rect 23112 36790 23164 36796
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 35834 23060 36722
rect 23492 36650 23520 39052
rect 23572 38956 23624 38962
rect 23572 38898 23624 38904
rect 23664 38956 23716 38962
rect 23664 38898 23716 38904
rect 23584 38554 23612 38898
rect 23572 38548 23624 38554
rect 23572 38490 23624 38496
rect 23676 37262 23704 38898
rect 23768 38554 23796 39986
rect 23940 39840 23992 39846
rect 23940 39782 23992 39788
rect 23952 39438 23980 39782
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 23940 39432 23992 39438
rect 24136 39409 24164 39986
rect 23940 39374 23992 39380
rect 24122 39400 24178 39409
rect 23860 39098 23888 39374
rect 24122 39335 24178 39344
rect 23940 39296 23992 39302
rect 23940 39238 23992 39244
rect 23848 39092 23900 39098
rect 23848 39034 23900 39040
rect 23848 38820 23900 38826
rect 23848 38762 23900 38768
rect 23756 38548 23808 38554
rect 23756 38490 23808 38496
rect 23860 38434 23888 38762
rect 23768 38406 23888 38434
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23664 37256 23716 37262
rect 23664 37198 23716 37204
rect 23480 36644 23532 36650
rect 23480 36586 23532 36592
rect 23584 36378 23612 37198
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23584 35834 23612 36110
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 23572 35828 23624 35834
rect 23572 35770 23624 35776
rect 23768 35714 23796 38406
rect 23952 38350 23980 39238
rect 24032 38752 24084 38758
rect 24032 38694 24084 38700
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 24044 38162 24072 38694
rect 23952 38134 24072 38162
rect 23848 37188 23900 37194
rect 23848 37130 23900 37136
rect 23860 36922 23888 37130
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 23952 36802 23980 38134
rect 24032 37868 24084 37874
rect 24032 37810 24084 37816
rect 24044 36922 24072 37810
rect 24124 37324 24176 37330
rect 24124 37266 24176 37272
rect 24136 37233 24164 37266
rect 24228 37262 24256 42026
rect 24400 39840 24452 39846
rect 24398 39808 24400 39817
rect 24452 39808 24454 39817
rect 24398 39743 24454 39752
rect 24400 38752 24452 38758
rect 24398 38720 24400 38729
rect 24452 38720 24454 38729
rect 24398 38655 24454 38664
rect 24400 37664 24452 37670
rect 24398 37632 24400 37641
rect 24452 37632 24454 37641
rect 24398 37567 24454 37576
rect 24216 37256 24268 37262
rect 24122 37224 24178 37233
rect 24216 37198 24268 37204
rect 24122 37159 24178 37168
rect 24032 36916 24084 36922
rect 24032 36858 24084 36864
rect 22940 35686 23060 35714
rect 22652 35148 22704 35154
rect 22652 35090 22704 35096
rect 22480 34734 22968 34762
rect 22560 33992 22612 33998
rect 22560 33934 22612 33940
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 22572 33289 22600 33934
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22664 33658 22692 33798
rect 22848 33658 22876 33934
rect 22652 33652 22704 33658
rect 22652 33594 22704 33600
rect 22836 33652 22888 33658
rect 22836 33594 22888 33600
rect 22742 33552 22798 33561
rect 22742 33487 22798 33496
rect 22558 33280 22614 33289
rect 22558 33215 22614 33224
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22296 30926 22508 30954
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22296 30054 22324 30670
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22112 26846 22232 26874
rect 21719 26684 22027 26693
rect 21719 26682 21725 26684
rect 21781 26682 21805 26684
rect 21861 26682 21885 26684
rect 21941 26682 21965 26684
rect 22021 26682 22027 26684
rect 21781 26630 21783 26682
rect 21963 26630 21965 26682
rect 21719 26628 21725 26630
rect 21781 26628 21805 26630
rect 21861 26628 21885 26630
rect 21941 26628 21965 26630
rect 22021 26628 22027 26630
rect 21719 26619 22027 26628
rect 21638 26208 21694 26217
rect 21638 26143 21694 26152
rect 21560 25996 21680 26024
rect 21364 25900 21416 25906
rect 21364 25842 21416 25848
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21376 25498 21404 25842
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21376 24954 21404 25434
rect 21364 24948 21416 24954
rect 21364 24890 21416 24896
rect 21468 24750 21496 25638
rect 21560 24954 21588 25842
rect 21548 24948 21600 24954
rect 21548 24890 21600 24896
rect 21652 24886 21680 25996
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 21719 25596 22027 25605
rect 21719 25594 21725 25596
rect 21781 25594 21805 25596
rect 21861 25594 21885 25596
rect 21941 25594 21965 25596
rect 22021 25594 22027 25596
rect 21781 25542 21783 25594
rect 21963 25542 21965 25594
rect 21719 25540 21725 25542
rect 21781 25540 21805 25542
rect 21861 25540 21885 25542
rect 21941 25540 21965 25542
rect 22021 25540 22027 25542
rect 21719 25531 22027 25540
rect 22112 25226 22140 25774
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 21640 24880 21692 24886
rect 22112 24857 22140 25162
rect 21640 24822 21692 24828
rect 22098 24848 22154 24857
rect 22098 24783 22154 24792
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 22100 24744 22152 24750
rect 22100 24686 22152 24692
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21468 24410 21496 24550
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21376 22216 21404 22918
rect 21376 22188 21496 22216
rect 21362 22128 21418 22137
rect 21362 22063 21418 22072
rect 21376 21894 21404 22063
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21272 21684 21324 21690
rect 21468 21672 21496 22188
rect 21272 21626 21324 21632
rect 21376 21644 21496 21672
rect 21376 21570 21404 21644
rect 21284 21542 21404 21570
rect 21456 21548 21508 21554
rect 21284 21026 21312 21542
rect 21456 21490 21508 21496
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21376 21146 21404 21286
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21284 20998 21404 21026
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 21100 19910 21220 19938
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 21100 19514 21128 19722
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 21086 19408 21142 19417
rect 21086 19343 21142 19352
rect 20916 19306 21036 19334
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20640 17338 20668 17478
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20536 17196 20588 17202
rect 20588 17156 20668 17184
rect 20536 17138 20588 17144
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20364 14414 20392 15030
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 12646 20392 13262
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20180 11206 20300 11234
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20088 10810 20116 11086
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20180 10690 20208 11206
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20088 10662 20208 10690
rect 19890 8392 19946 8401
rect 19890 8327 19946 8336
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19904 7546 19932 7822
rect 19996 7818 20024 8230
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 20088 7698 20116 10662
rect 20272 10266 20300 11086
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20180 8090 20208 8434
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20364 7970 20392 11698
rect 20456 10198 20484 15302
rect 20536 13320 20588 13326
rect 20534 13288 20536 13297
rect 20588 13288 20590 13297
rect 20534 13223 20590 13232
rect 20536 12912 20588 12918
rect 20536 12854 20588 12860
rect 20548 12238 20576 12854
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20640 11014 20668 17156
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 16114 20760 16390
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20824 15994 20852 19110
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20916 17338 20944 17546
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20902 16688 20958 16697
rect 20902 16623 20958 16632
rect 20732 15966 20852 15994
rect 20732 12594 20760 15966
rect 20812 15564 20864 15570
rect 20812 15506 20864 15512
rect 20824 15162 20852 15506
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20824 13530 20852 14554
rect 20916 13705 20944 16623
rect 21008 15366 21036 19306
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20902 13696 20958 13705
rect 20902 13631 20958 13640
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20996 12776 21048 12782
rect 20996 12718 21048 12724
rect 20732 12566 20944 12594
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20732 11286 20760 12038
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20732 10810 20760 11086
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20732 10470 20760 10610
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20732 10266 20760 10406
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9586 20576 9862
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 19996 7670 20116 7698
rect 20180 7942 20392 7970
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19812 7364 19932 7392
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 19168 5766 19288 5794
rect 19076 5574 19104 5714
rect 19064 5568 19116 5574
rect 19064 5510 19116 5516
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18708 5273 18736 5306
rect 18694 5264 18750 5273
rect 19168 5250 19196 5766
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 18694 5199 18750 5208
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 19076 5222 19196 5250
rect 18800 4758 18828 5170
rect 18984 4758 19012 5170
rect 18788 4752 18840 4758
rect 18616 4678 18736 4706
rect 18788 4694 18840 4700
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18604 4616 18656 4622
rect 18524 4576 18604 4604
rect 18604 4558 18656 4564
rect 18708 4468 18736 4678
rect 19076 4604 19104 5222
rect 19260 5098 19288 5510
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19352 4865 19380 7278
rect 19444 7262 19840 7290
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19628 6798 19656 6938
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19430 6488 19486 6497
rect 19430 6423 19486 6432
rect 19444 6225 19472 6423
rect 19430 6216 19486 6225
rect 19430 6151 19486 6160
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19536 5386 19564 5510
rect 19444 5358 19564 5386
rect 19444 5234 19472 5358
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19338 4856 19394 4865
rect 19260 4826 19338 4842
rect 19248 4820 19338 4826
rect 19300 4814 19338 4820
rect 19338 4791 19394 4800
rect 19248 4762 19300 4768
rect 19248 4616 19300 4622
rect 19076 4576 19196 4604
rect 18616 4440 18736 4468
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18328 3936 18380 3942
rect 18524 3913 18552 4082
rect 18328 3878 18380 3884
rect 18510 3904 18566 3913
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18144 1828 18196 1834
rect 18144 1770 18196 1776
rect 18052 1012 18104 1018
rect 18052 954 18104 960
rect 17314 54 17448 82
rect 17314 0 17370 54
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 82 18198 160
rect 18248 82 18276 2246
rect 18340 1358 18368 3878
rect 18510 3839 18566 3848
rect 18420 3732 18472 3738
rect 18616 3720 18644 4440
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 19064 4140 19116 4146
rect 19168 4128 19196 4576
rect 19248 4558 19300 4564
rect 19116 4100 19196 4128
rect 19064 4082 19116 4088
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18472 3692 18644 3720
rect 18420 3674 18472 3680
rect 18708 3482 18736 3878
rect 18512 3460 18564 3466
rect 18512 3402 18564 3408
rect 18616 3454 18736 3482
rect 18524 3194 18552 3402
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18616 3126 18644 3454
rect 18800 3398 18828 4082
rect 19260 4010 19288 4558
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19156 3936 19208 3942
rect 19352 3890 19380 4791
rect 19444 4622 19472 5170
rect 19536 4826 19564 5238
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19444 3890 19472 4014
rect 19156 3878 19208 3884
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 18972 2916 19024 2922
rect 18972 2858 19024 2864
rect 18788 2848 18840 2854
rect 18616 2808 18788 2836
rect 18512 2372 18564 2378
rect 18512 2314 18564 2320
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 18432 160 18460 2246
rect 18524 1426 18552 2314
rect 18512 1420 18564 1426
rect 18512 1362 18564 1368
rect 18616 898 18644 2808
rect 18788 2790 18840 2796
rect 18984 2514 19012 2858
rect 19076 2582 19104 2994
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 18788 1896 18840 1902
rect 18788 1838 18840 1844
rect 18800 1562 18828 1838
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 19064 1352 19116 1358
rect 19062 1320 19064 1329
rect 19116 1320 19118 1329
rect 19062 1255 19118 1264
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 18616 870 18736 898
rect 18708 160 18736 870
rect 18142 54 18276 82
rect 18142 0 18198 54
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 82 19026 160
rect 19168 82 19196 3878
rect 19260 3862 19472 3890
rect 19616 3936 19668 3942
rect 19616 3878 19668 3884
rect 19260 3534 19288 3862
rect 19444 3754 19472 3862
rect 19444 3726 19564 3754
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19260 160 19288 3334
rect 19352 2446 19380 3334
rect 19536 2650 19564 3726
rect 19628 2990 19656 3878
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19444 2106 19472 2586
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 19524 2372 19576 2378
rect 19524 2314 19576 2320
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19536 1766 19564 2314
rect 19628 2106 19656 2518
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19524 1760 19576 1766
rect 19524 1702 19576 1708
rect 18970 54 19196 82
rect 18970 0 19026 54
rect 19246 0 19302 160
rect 19522 82 19578 160
rect 19720 82 19748 3334
rect 19812 2990 19840 7262
rect 19904 6390 19932 7364
rect 19892 6384 19944 6390
rect 19892 6326 19944 6332
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19904 4729 19932 5306
rect 19890 4720 19946 4729
rect 19890 4655 19946 4664
rect 19996 4622 20024 7670
rect 20180 6186 20208 7942
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20272 7002 20300 7346
rect 20260 6996 20312 7002
rect 20260 6938 20312 6944
rect 20364 6934 20392 7822
rect 20456 7585 20484 8842
rect 20442 7576 20498 7585
rect 20442 7511 20498 7520
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20352 6928 20404 6934
rect 20352 6870 20404 6876
rect 20456 6798 20484 7346
rect 20548 6934 20576 9522
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7546 20668 7822
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20626 7440 20682 7449
rect 20732 7410 20760 10202
rect 20626 7375 20682 7384
rect 20720 7404 20772 7410
rect 20536 6928 20588 6934
rect 20536 6870 20588 6876
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20640 6610 20668 7375
rect 20720 7346 20772 7352
rect 20732 6730 20760 7346
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20456 6582 20668 6610
rect 20718 6624 20774 6633
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20272 6225 20300 6258
rect 20258 6216 20314 6225
rect 20168 6180 20220 6186
rect 20258 6151 20314 6160
rect 20168 6122 20220 6128
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20088 5370 20116 6054
rect 20350 5536 20406 5545
rect 20350 5471 20406 5480
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19904 4282 20024 4298
rect 20088 4282 20116 4558
rect 20180 4486 20208 5238
rect 20364 4622 20392 5471
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 19892 4276 20024 4282
rect 19944 4270 20024 4276
rect 19892 4218 19944 4224
rect 19996 4162 20024 4270
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 19892 4140 19944 4146
rect 19996 4134 20208 4162
rect 19892 4082 19944 4088
rect 19904 3534 19932 4082
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19904 3194 19932 3470
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19996 3097 20024 3402
rect 19982 3088 20038 3097
rect 19982 3023 20038 3032
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19522 54 19748 82
rect 19798 82 19854 160
rect 19996 82 20024 2790
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20088 160 20116 2586
rect 20180 2378 20208 4134
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 20168 1964 20220 1970
rect 20168 1906 20220 1912
rect 19798 54 20024 82
rect 19522 0 19578 54
rect 19798 0 19854 54
rect 20074 0 20130 160
rect 20180 82 20208 1906
rect 20272 1902 20300 4422
rect 20364 4146 20392 4422
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20456 2990 20484 6582
rect 20718 6559 20774 6568
rect 20732 6474 20760 6559
rect 20640 6446 20760 6474
rect 20640 6390 20668 6446
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5409 20576 6258
rect 20628 6180 20680 6186
rect 20628 6122 20680 6128
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20640 6089 20668 6122
rect 20626 6080 20682 6089
rect 20626 6015 20682 6024
rect 20732 5914 20760 6122
rect 20824 6100 20852 12174
rect 20916 7750 20944 12566
rect 21008 12442 21036 12718
rect 21100 12628 21128 19343
rect 21192 19258 21220 19910
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21284 19378 21312 19790
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21192 19230 21312 19258
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21192 14226 21220 18634
rect 21284 16182 21312 19230
rect 21376 18426 21404 20998
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21468 16776 21496 21490
rect 21560 18970 21588 24550
rect 21719 24508 22027 24517
rect 21719 24506 21725 24508
rect 21781 24506 21805 24508
rect 21861 24506 21885 24508
rect 21941 24506 21965 24508
rect 22021 24506 22027 24508
rect 21781 24454 21783 24506
rect 21963 24454 21965 24506
rect 21719 24452 21725 24454
rect 21781 24452 21805 24454
rect 21861 24452 21885 24454
rect 21941 24452 21965 24454
rect 22021 24452 22027 24454
rect 21719 24443 22027 24452
rect 21638 23760 21694 23769
rect 21638 23695 21640 23704
rect 21692 23695 21694 23704
rect 21640 23666 21692 23672
rect 21719 23420 22027 23429
rect 21719 23418 21725 23420
rect 21781 23418 21805 23420
rect 21861 23418 21885 23420
rect 21941 23418 21965 23420
rect 22021 23418 22027 23420
rect 21781 23366 21783 23418
rect 21963 23366 21965 23418
rect 21719 23364 21725 23366
rect 21781 23364 21805 23366
rect 21861 23364 21885 23366
rect 21941 23364 21965 23366
rect 22021 23364 22027 23366
rect 21719 23355 22027 23364
rect 21732 23112 21784 23118
rect 22112 23066 22140 24686
rect 22204 23497 22232 26846
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22388 23866 22416 24754
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22190 23488 22246 23497
rect 22190 23423 22246 23432
rect 22376 23112 22428 23118
rect 21732 23054 21784 23060
rect 21744 22778 21772 23054
rect 22020 23038 22324 23066
rect 22376 23054 22428 23060
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 22020 22642 22048 23038
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21652 22545 21680 22578
rect 21732 22568 21784 22574
rect 21638 22536 21694 22545
rect 21732 22510 21784 22516
rect 21638 22471 21694 22480
rect 21744 22420 21772 22510
rect 21652 22392 21772 22420
rect 21652 22166 21680 22392
rect 21719 22332 22027 22341
rect 21719 22330 21725 22332
rect 21781 22330 21805 22332
rect 21861 22330 21885 22332
rect 21941 22330 21965 22332
rect 22021 22330 22027 22332
rect 21781 22278 21783 22330
rect 21963 22278 21965 22330
rect 21719 22276 21725 22278
rect 21781 22276 21805 22278
rect 21861 22276 21885 22278
rect 21941 22276 21965 22278
rect 22021 22276 22027 22278
rect 21719 22267 22027 22276
rect 21640 22160 21692 22166
rect 21640 22102 21692 22108
rect 22112 22030 22140 22918
rect 22204 22234 22232 22918
rect 22296 22778 22324 23038
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22296 22098 22324 22374
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21652 17785 21680 21830
rect 22296 21690 22324 21830
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 21719 21244 22027 21253
rect 21719 21242 21725 21244
rect 21781 21242 21805 21244
rect 21861 21242 21885 21244
rect 21941 21242 21965 21244
rect 22021 21242 22027 21244
rect 21781 21190 21783 21242
rect 21963 21190 21965 21242
rect 21719 21188 21725 21190
rect 21781 21188 21805 21190
rect 21861 21188 21885 21190
rect 21941 21188 21965 21190
rect 22021 21188 22027 21190
rect 21719 21179 22027 21188
rect 22388 20942 22416 23054
rect 22480 22930 22508 30926
rect 22560 30592 22612 30598
rect 22560 30534 22612 30540
rect 22572 29646 22600 30534
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22572 25294 22600 27814
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22480 22902 22600 22930
rect 22466 22536 22522 22545
rect 22466 22471 22522 22480
rect 22480 22166 22508 22471
rect 22468 22160 22520 22166
rect 22468 22102 22520 22108
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21719 20156 22027 20165
rect 21719 20154 21725 20156
rect 21781 20154 21805 20156
rect 21861 20154 21885 20156
rect 21941 20154 21965 20156
rect 22021 20154 22027 20156
rect 21781 20102 21783 20154
rect 21963 20102 21965 20154
rect 21719 20100 21725 20102
rect 21781 20100 21805 20102
rect 21861 20100 21885 20102
rect 21941 20100 21965 20102
rect 22021 20100 22027 20102
rect 21719 20091 22027 20100
rect 22112 20058 22140 20402
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22296 20058 22324 20334
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 21719 19068 22027 19077
rect 21719 19066 21725 19068
rect 21781 19066 21805 19068
rect 21861 19066 21885 19068
rect 21941 19066 21965 19068
rect 22021 19066 22027 19068
rect 21781 19014 21783 19066
rect 21963 19014 21965 19066
rect 21719 19012 21725 19014
rect 21781 19012 21805 19014
rect 21861 19012 21885 19014
rect 21941 19012 21965 19014
rect 22021 19012 22027 19014
rect 21719 19003 22027 19012
rect 21719 17980 22027 17989
rect 21719 17978 21725 17980
rect 21781 17978 21805 17980
rect 21861 17978 21885 17980
rect 21941 17978 21965 17980
rect 22021 17978 22027 17980
rect 21781 17926 21783 17978
rect 21963 17926 21965 17978
rect 21719 17924 21725 17926
rect 21781 17924 21805 17926
rect 21861 17924 21885 17926
rect 21941 17924 21965 17926
rect 22021 17924 22027 17926
rect 21719 17915 22027 17924
rect 22204 17814 22232 19450
rect 22388 18290 22416 20878
rect 22480 20602 22508 20878
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22388 17882 22416 18226
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22192 17808 22244 17814
rect 21638 17776 21694 17785
rect 22192 17750 22244 17756
rect 21638 17711 21694 17720
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 21824 17128 21876 17134
rect 22112 17082 22140 17682
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 17338 22232 17614
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 21876 17076 22140 17082
rect 21824 17070 22140 17076
rect 21640 17060 21692 17066
rect 21836 17054 22140 17070
rect 21640 17002 21692 17008
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16794 21588 16934
rect 21376 16748 21496 16776
rect 21548 16788 21600 16794
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 21376 16130 21404 16748
rect 21548 16730 21600 16736
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21468 16250 21496 16594
rect 21652 16590 21680 17002
rect 21719 16892 22027 16901
rect 21719 16890 21725 16892
rect 21781 16890 21805 16892
rect 21861 16890 21885 16892
rect 21941 16890 21965 16892
rect 22021 16890 22027 16892
rect 21781 16838 21783 16890
rect 21963 16838 21965 16890
rect 21719 16836 21725 16838
rect 21781 16836 21805 16838
rect 21861 16836 21885 16838
rect 21941 16836 21965 16838
rect 22021 16836 22027 16838
rect 21719 16827 22027 16836
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21548 16244 21600 16250
rect 21548 16186 21600 16192
rect 21376 16102 21496 16130
rect 21192 14198 21404 14226
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21192 13784 21220 14010
rect 21192 13756 21312 13784
rect 21284 13462 21312 13756
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 21180 12640 21232 12646
rect 21100 12600 21180 12628
rect 21180 12582 21232 12588
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 21008 10810 21036 12378
rect 21284 12306 21312 13398
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21376 11744 21404 14198
rect 21192 11716 21404 11744
rect 21192 11150 21220 11716
rect 21468 11642 21496 16102
rect 21560 13938 21588 16186
rect 22112 15910 22140 17054
rect 22296 16794 22324 17478
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22190 16144 22246 16153
rect 22246 16102 22324 16130
rect 22190 16079 22246 16088
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 21719 15804 22027 15813
rect 21719 15802 21725 15804
rect 21781 15802 21805 15804
rect 21861 15802 21885 15804
rect 21941 15802 21965 15804
rect 22021 15802 22027 15804
rect 21781 15750 21783 15802
rect 21963 15750 21965 15802
rect 21719 15748 21725 15750
rect 21781 15748 21805 15750
rect 21861 15748 21885 15750
rect 21941 15748 21965 15750
rect 22021 15748 22027 15750
rect 21719 15739 22027 15748
rect 22296 15502 22324 16102
rect 22388 15570 22416 17818
rect 22480 17746 22508 19994
rect 22468 17740 22520 17746
rect 22468 17682 22520 17688
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 17338 22508 17478
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22376 15564 22428 15570
rect 22376 15506 22428 15512
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 21744 14958 21772 15438
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 22112 15162 22140 15302
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 21732 14952 21784 14958
rect 21732 14894 21784 14900
rect 21640 14816 21692 14822
rect 21640 14758 21692 14764
rect 21652 14482 21680 14758
rect 21719 14716 22027 14725
rect 21719 14714 21725 14716
rect 21781 14714 21805 14716
rect 21861 14714 21885 14716
rect 21941 14714 21965 14716
rect 22021 14714 22027 14716
rect 21781 14662 21783 14714
rect 21963 14662 21965 14714
rect 21719 14660 21725 14662
rect 21781 14660 21805 14662
rect 21861 14660 21885 14662
rect 21941 14660 21965 14662
rect 22021 14660 22027 14662
rect 21719 14651 22027 14660
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 22204 14414 22232 14962
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22100 14272 22152 14278
rect 22100 14214 22152 14220
rect 21640 14000 21692 14006
rect 22112 13977 22140 14214
rect 21640 13942 21692 13948
rect 22098 13968 22154 13977
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21560 12714 21588 13262
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11762 21588 12106
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21284 11614 21496 11642
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 21008 6610 21036 10406
rect 21100 9722 21128 10610
rect 21088 9716 21140 9722
rect 21284 9674 21312 11614
rect 21456 11008 21508 11014
rect 21456 10950 21508 10956
rect 21088 9658 21140 9664
rect 21192 9646 21312 9674
rect 21192 9058 21220 9646
rect 21100 9030 21220 9058
rect 21272 9036 21324 9042
rect 21100 8498 21128 9030
rect 21272 8978 21324 8984
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21284 7954 21312 8978
rect 21272 7948 21324 7954
rect 21272 7890 21324 7896
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 21100 7002 21128 7822
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21272 7268 21324 7274
rect 21272 7210 21324 7216
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21192 6798 21220 7142
rect 21284 7002 21312 7210
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21270 6896 21326 6905
rect 21270 6831 21326 6840
rect 21284 6798 21312 6831
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 20916 6582 21036 6610
rect 21100 6610 21128 6666
rect 21100 6582 21220 6610
rect 20916 6440 20944 6582
rect 21088 6452 21140 6458
rect 20916 6412 21036 6440
rect 20904 6112 20956 6118
rect 20824 6072 20904 6100
rect 20904 6054 20956 6060
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 21008 5794 21036 6412
rect 21088 6394 21140 6400
rect 20916 5766 21036 5794
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20534 5400 20590 5409
rect 20534 5335 20590 5344
rect 20732 5137 20760 5646
rect 20812 5160 20864 5166
rect 20718 5128 20774 5137
rect 20812 5102 20864 5108
rect 20718 5063 20774 5072
rect 20536 5024 20588 5030
rect 20588 4984 20668 5012
rect 20536 4966 20588 4972
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20548 3346 20576 4558
rect 20640 4282 20668 4984
rect 20824 4842 20852 5102
rect 20916 5098 20944 5766
rect 21100 5710 21128 6394
rect 21192 6186 21220 6582
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21180 5840 21232 5846
rect 21178 5808 21180 5817
rect 21232 5808 21234 5817
rect 21178 5743 21234 5752
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20904 5092 20956 5098
rect 20904 5034 20956 5040
rect 21008 5030 21036 5646
rect 21180 5228 21232 5234
rect 21100 5188 21180 5216
rect 20996 5024 21048 5030
rect 20996 4966 21048 4972
rect 20824 4814 21036 4842
rect 21100 4826 21128 5188
rect 21180 5170 21232 5176
rect 21180 5092 21232 5098
rect 21180 5034 21232 5040
rect 21192 4826 21220 5034
rect 20904 4752 20956 4758
rect 20904 4694 20956 4700
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3466 20668 4082
rect 20732 3534 20760 4626
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20824 3738 20852 4558
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20718 3360 20774 3369
rect 20548 3318 20718 3346
rect 20718 3295 20774 3304
rect 20916 3126 20944 4694
rect 21008 4672 21036 4814
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21088 4684 21140 4690
rect 21008 4644 21088 4672
rect 21088 4626 21140 4632
rect 21284 4593 21312 6190
rect 21270 4584 21326 4593
rect 21270 4519 21326 4528
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 21008 3602 21036 4218
rect 21086 4040 21142 4049
rect 21086 3975 21088 3984
rect 21140 3975 21142 3984
rect 21088 3946 21140 3952
rect 20996 3596 21048 3602
rect 21048 3556 21128 3584
rect 20996 3538 21048 3544
rect 20904 3120 20956 3126
rect 20904 3062 20956 3068
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20444 2984 20496 2990
rect 20732 2961 20760 2994
rect 20444 2926 20496 2932
rect 20718 2952 20774 2961
rect 20628 2916 20680 2922
rect 20718 2887 20774 2896
rect 20628 2858 20680 2864
rect 20534 2680 20590 2689
rect 20534 2615 20590 2624
rect 20260 1896 20312 1902
rect 20260 1838 20312 1844
rect 20548 1494 20576 2615
rect 20640 1850 20668 2858
rect 21100 2514 21128 3556
rect 21192 3505 21220 4422
rect 21178 3496 21234 3505
rect 21178 3431 21234 3440
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 20812 1964 20864 1970
rect 20812 1906 20864 1912
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 20718 1864 20774 1873
rect 20640 1822 20718 1850
rect 20718 1799 20774 1808
rect 20536 1488 20588 1494
rect 20536 1430 20588 1436
rect 20628 1352 20680 1358
rect 20628 1294 20680 1300
rect 20640 160 20668 1294
rect 20720 1012 20772 1018
rect 20720 954 20772 960
rect 20732 649 20760 954
rect 20718 640 20774 649
rect 20718 575 20774 584
rect 20350 82 20406 160
rect 20180 54 20406 82
rect 20350 0 20406 54
rect 20626 0 20682 160
rect 20824 82 20852 1906
rect 21100 1408 21128 1906
rect 21192 1426 21220 2382
rect 21008 1380 21128 1408
rect 21180 1420 21232 1426
rect 21008 490 21036 1380
rect 21180 1362 21232 1368
rect 21088 1284 21140 1290
rect 21088 1226 21140 1232
rect 21180 1284 21232 1290
rect 21180 1226 21232 1232
rect 21100 678 21128 1226
rect 21192 1018 21220 1226
rect 21180 1012 21232 1018
rect 21180 954 21232 960
rect 21088 672 21140 678
rect 21088 614 21140 620
rect 21008 462 21220 490
rect 21192 160 21220 462
rect 20902 82 20958 160
rect 20824 54 20958 82
rect 20902 0 20958 54
rect 21178 0 21234 160
rect 21284 82 21312 2994
rect 21376 2774 21404 7686
rect 21468 5574 21496 10950
rect 21546 7848 21602 7857
rect 21546 7783 21602 7792
rect 21560 6798 21588 7783
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21548 6112 21600 6118
rect 21546 6080 21548 6089
rect 21600 6080 21602 6089
rect 21546 6015 21602 6024
rect 21652 5930 21680 13942
rect 22098 13903 22154 13912
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 22100 13728 22152 13734
rect 22098 13696 22100 13705
rect 22152 13696 22154 13705
rect 21719 13628 22027 13637
rect 22098 13631 22154 13640
rect 21719 13626 21725 13628
rect 21781 13626 21805 13628
rect 21861 13626 21885 13628
rect 21941 13626 21965 13628
rect 22021 13626 22027 13628
rect 21781 13574 21783 13626
rect 21963 13574 21965 13626
rect 21719 13572 21725 13574
rect 21781 13572 21805 13574
rect 21861 13572 21885 13574
rect 21941 13572 21965 13574
rect 22021 13572 22027 13574
rect 21719 13563 22027 13572
rect 22204 12850 22232 13738
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21719 12540 22027 12549
rect 21719 12538 21725 12540
rect 21781 12538 21805 12540
rect 21861 12538 21885 12540
rect 21941 12538 21965 12540
rect 22021 12538 22027 12540
rect 21781 12486 21783 12538
rect 21963 12486 21965 12538
rect 21719 12484 21725 12486
rect 21781 12484 21805 12486
rect 21861 12484 21885 12486
rect 21941 12484 21965 12486
rect 22021 12484 22027 12486
rect 21719 12475 22027 12484
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11830 21864 12038
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21719 11452 22027 11461
rect 21719 11450 21725 11452
rect 21781 11450 21805 11452
rect 21861 11450 21885 11452
rect 21941 11450 21965 11452
rect 22021 11450 22027 11452
rect 21781 11398 21783 11450
rect 21963 11398 21965 11450
rect 21719 11396 21725 11398
rect 21781 11396 21805 11398
rect 21861 11396 21885 11398
rect 21941 11396 21965 11398
rect 22021 11396 22027 11398
rect 21719 11387 22027 11396
rect 21719 10364 22027 10373
rect 21719 10362 21725 10364
rect 21781 10362 21805 10364
rect 21861 10362 21885 10364
rect 21941 10362 21965 10364
rect 22021 10362 22027 10364
rect 21781 10310 21783 10362
rect 21963 10310 21965 10362
rect 21719 10308 21725 10310
rect 21781 10308 21805 10310
rect 21861 10308 21885 10310
rect 21941 10308 21965 10310
rect 22021 10308 22027 10310
rect 21719 10299 22027 10308
rect 22112 10198 22140 12582
rect 22296 11286 22324 14758
rect 22388 13462 22416 15506
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22480 14414 22508 14962
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22572 13682 22600 22902
rect 22664 22642 22692 32710
rect 22756 28626 22784 33487
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 22848 29850 22876 29990
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22940 28694 22968 34734
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22744 28212 22796 28218
rect 22744 28154 22796 28160
rect 22756 27470 22784 28154
rect 22940 28082 22968 28630
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22928 28076 22980 28082
rect 22928 28018 22980 28024
rect 22848 27674 22876 28018
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 22744 27464 22796 27470
rect 23032 27418 23060 35686
rect 23584 35686 23796 35714
rect 23860 36774 23980 36802
rect 24032 36780 24084 36786
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23296 34740 23348 34746
rect 23296 34682 23348 34688
rect 23112 34400 23164 34406
rect 23112 34342 23164 34348
rect 23124 33522 23152 34342
rect 23204 33924 23256 33930
rect 23204 33866 23256 33872
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 23216 32842 23244 33866
rect 23308 32842 23336 34682
rect 23400 34202 23428 35022
rect 23480 34944 23532 34950
rect 23480 34886 23532 34892
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23492 33998 23520 34886
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23400 33114 23428 33254
rect 23388 33108 23440 33114
rect 23388 33050 23440 33056
rect 23204 32836 23256 32842
rect 23204 32778 23256 32784
rect 23296 32836 23348 32842
rect 23296 32778 23348 32784
rect 23204 31816 23256 31822
rect 23202 31784 23204 31793
rect 23256 31784 23258 31793
rect 23202 31719 23258 31728
rect 23584 31754 23612 35686
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23676 34746 23704 35226
rect 23768 34746 23796 35430
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23756 34740 23808 34746
rect 23756 34682 23808 34688
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23676 33658 23704 33798
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 23860 31754 23888 36774
rect 24032 36722 24084 36728
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 23940 35692 23992 35698
rect 23940 35634 23992 35640
rect 23952 34678 23980 35634
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 23952 32570 23980 32846
rect 23940 32564 23992 32570
rect 23940 32506 23992 32512
rect 24044 32230 24072 36722
rect 24400 36576 24452 36582
rect 24398 36544 24400 36553
rect 24452 36544 24454 36553
rect 24398 36479 24454 36488
rect 24400 35488 24452 35494
rect 24398 35456 24400 35465
rect 24452 35456 24454 35465
rect 24398 35391 24454 35400
rect 24216 35012 24268 35018
rect 24216 34954 24268 34960
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 24136 32026 24164 32370
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24228 31754 24256 34954
rect 24400 34536 24452 34542
rect 24398 34504 24400 34513
rect 24452 34504 24454 34513
rect 24398 34439 24454 34448
rect 24400 33312 24452 33318
rect 24398 33280 24400 33289
rect 24452 33280 24454 33289
rect 24398 33215 24454 33224
rect 24400 32224 24452 32230
rect 24398 32192 24400 32201
rect 24452 32192 24454 32201
rect 24398 32127 24454 32136
rect 23584 31726 23704 31754
rect 23860 31726 24072 31754
rect 23296 31272 23348 31278
rect 23296 31214 23348 31220
rect 23308 30734 23336 31214
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23296 30252 23348 30258
rect 23296 30194 23348 30200
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 23216 29850 23244 29990
rect 23204 29844 23256 29850
rect 23204 29786 23256 29792
rect 23112 29028 23164 29034
rect 23112 28970 23164 28976
rect 22744 27406 22796 27412
rect 22836 27396 22888 27402
rect 22836 27338 22888 27344
rect 22940 27390 23060 27418
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 26790 22784 27270
rect 22848 27130 22876 27338
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 22744 26784 22796 26790
rect 22744 26726 22796 26732
rect 22940 24857 22968 27390
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23032 27130 23060 27270
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 23124 27010 23152 28970
rect 23202 28656 23258 28665
rect 23308 28642 23336 30194
rect 23258 28614 23336 28642
rect 23202 28591 23258 28600
rect 23032 26982 23152 27010
rect 22926 24848 22982 24857
rect 22926 24783 22982 24792
rect 23032 24698 23060 26982
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23124 25498 23152 25638
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23216 25378 23244 28591
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 22940 24670 23060 24698
rect 23124 25350 23244 25378
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22756 23050 22784 23666
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22652 22636 22704 22642
rect 22652 22578 22704 22584
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22664 20466 22692 20810
rect 22756 20466 22784 22646
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22848 22234 22876 22374
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22940 22094 22968 24670
rect 23124 22094 23152 25350
rect 23308 23866 23336 28494
rect 23676 27962 23704 31726
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23860 30394 23888 31282
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23952 30394 23980 31078
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23676 27934 23888 27962
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 23492 27470 23520 27814
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23584 27130 23612 27406
rect 23768 27130 23796 27814
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23756 27124 23808 27130
rect 23756 27066 23808 27072
rect 23756 26988 23808 26994
rect 23756 26930 23808 26936
rect 23768 26586 23796 26930
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23400 24410 23428 25774
rect 23492 25362 23520 26318
rect 23584 26042 23612 26318
rect 23664 26240 23716 26246
rect 23664 26182 23716 26188
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23584 25498 23612 25842
rect 23676 25498 23704 26182
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23492 24954 23520 25298
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23216 22778 23244 23666
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 22848 22066 22968 22094
rect 23032 22066 23152 22094
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22652 20324 22704 20330
rect 22652 20266 22704 20272
rect 22664 19378 22692 20266
rect 22848 20262 22876 22066
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22836 20256 22888 20262
rect 22836 20198 22888 20204
rect 22940 19378 22968 20402
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 23032 18850 23060 22066
rect 23112 22024 23164 22030
rect 23216 21978 23244 22714
rect 23308 22098 23336 23462
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23400 21978 23428 24006
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23164 21972 23244 21978
rect 23112 21966 23244 21972
rect 23124 21950 23244 21966
rect 23308 21950 23428 21978
rect 23492 21962 23520 22578
rect 23584 22234 23612 23462
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23676 22094 23704 24142
rect 23768 23118 23796 25094
rect 23860 24410 23888 27934
rect 23952 27674 23980 28018
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 23940 26784 23992 26790
rect 23940 26726 23992 26732
rect 23952 25922 23980 26726
rect 24044 26042 24072 31726
rect 24136 31726 24256 31754
rect 24032 26036 24084 26042
rect 24032 25978 24084 25984
rect 24136 25974 24164 31726
rect 24400 31136 24452 31142
rect 24398 31104 24400 31113
rect 24452 31104 24454 31113
rect 24398 31039 24454 31048
rect 24400 30048 24452 30054
rect 24398 30016 24400 30025
rect 24452 30016 24454 30025
rect 24398 29951 24454 29960
rect 24308 29572 24360 29578
rect 24308 29514 24360 29520
rect 24214 26208 24270 26217
rect 24214 26143 24270 26152
rect 24124 25968 24176 25974
rect 23952 25894 24072 25922
rect 24124 25910 24176 25916
rect 23940 25764 23992 25770
rect 23940 25706 23992 25712
rect 23848 24404 23900 24410
rect 23848 24346 23900 24352
rect 23846 24304 23902 24313
rect 23846 24239 23902 24248
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23860 22094 23888 24239
rect 23952 24206 23980 25706
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23952 23322 23980 23666
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 24044 22094 24072 25894
rect 23676 22066 23796 22094
rect 23860 22066 23980 22094
rect 24044 22066 24164 22094
rect 23480 21956 23532 21962
rect 23308 21876 23336 21950
rect 23480 21898 23532 21904
rect 23768 21894 23796 22066
rect 23124 21848 23336 21876
rect 23388 21888 23440 21894
rect 23124 19394 23152 21848
rect 23388 21830 23440 21836
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23216 19514 23244 19654
rect 23308 19514 23336 20742
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23124 19366 23244 19394
rect 22756 18822 23060 18850
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22480 13654 22600 13682
rect 22376 13456 22428 13462
rect 22376 13398 22428 13404
rect 22480 12986 22508 13654
rect 22558 13560 22614 13569
rect 22558 13495 22560 13504
rect 22612 13495 22614 13504
rect 22560 13466 22612 13472
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22468 12854 22520 12860
rect 22468 12796 22520 12802
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22296 10130 22324 11222
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22284 10124 22336 10130
rect 22284 10066 22336 10072
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22204 9586 22232 9862
rect 22296 9722 22324 9862
rect 22388 9722 22416 11154
rect 22480 10266 22508 12796
rect 22572 11558 22600 13262
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22560 10464 22612 10470
rect 22560 10406 22612 10412
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22376 9580 22428 9586
rect 22376 9522 22428 9528
rect 22204 9466 22232 9522
rect 22204 9438 22324 9466
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 21719 9276 22027 9285
rect 21719 9274 21725 9276
rect 21781 9274 21805 9276
rect 21861 9274 21885 9276
rect 21941 9274 21965 9276
rect 22021 9274 22027 9276
rect 21781 9222 21783 9274
rect 21963 9222 21965 9274
rect 21719 9220 21725 9222
rect 21781 9220 21805 9222
rect 21861 9220 21885 9222
rect 21941 9220 21965 9222
rect 22021 9220 22027 9222
rect 21719 9211 22027 9220
rect 22008 8832 22060 8838
rect 22008 8774 22060 8780
rect 22020 8514 22048 8774
rect 22112 8634 22140 9318
rect 22204 8634 22232 9318
rect 22100 8628 22152 8634
rect 22100 8570 22152 8576
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22020 8486 22232 8514
rect 22204 8242 22232 8486
rect 22296 8430 22324 9438
rect 22388 8906 22416 9522
rect 22480 9178 22508 9998
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22572 8974 22600 10406
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22376 8900 22428 8906
rect 22376 8842 22428 8848
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22204 8214 22508 8242
rect 21719 8188 22027 8197
rect 21719 8186 21725 8188
rect 21781 8186 21805 8188
rect 21861 8186 21885 8188
rect 21941 8186 21965 8188
rect 22021 8186 22027 8188
rect 21781 8134 21783 8186
rect 21963 8134 21965 8186
rect 21719 8132 21725 8134
rect 21781 8132 21805 8134
rect 21861 8132 21885 8134
rect 21941 8132 21965 8134
rect 22021 8132 22027 8134
rect 21719 8123 22027 8132
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 21719 7100 22027 7109
rect 21719 7098 21725 7100
rect 21781 7098 21805 7100
rect 21861 7098 21885 7100
rect 21941 7098 21965 7100
rect 22021 7098 22027 7100
rect 21781 7046 21783 7098
rect 21963 7046 21965 7098
rect 21719 7044 21725 7046
rect 21781 7044 21805 7046
rect 21861 7044 21885 7046
rect 21941 7044 21965 7046
rect 22021 7044 22027 7046
rect 21719 7035 22027 7044
rect 21730 6896 21786 6905
rect 21730 6831 21786 6840
rect 21744 6361 21772 6831
rect 22112 6662 22140 7686
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 21916 6656 21968 6662
rect 21916 6598 21968 6604
rect 22100 6656 22152 6662
rect 22204 6644 22232 7278
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 22204 6616 22324 6644
rect 22100 6598 22152 6604
rect 21928 6474 21956 6598
rect 21928 6458 22094 6474
rect 21928 6452 22106 6458
rect 21928 6446 22054 6452
rect 22054 6394 22106 6400
rect 21730 6352 21786 6361
rect 21730 6287 21786 6296
rect 21824 6316 21876 6322
rect 22020 6310 22140 6338
rect 22020 6304 22048 6310
rect 21876 6276 22048 6304
rect 21824 6258 21876 6264
rect 22112 6202 22140 6310
rect 22296 6202 22324 6616
rect 22112 6174 22324 6202
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 21560 5902 21680 5930
rect 21560 5828 21588 5902
rect 21560 5800 21680 5828
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21560 5386 21588 5646
rect 21468 5358 21588 5386
rect 21468 5098 21496 5358
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21456 5092 21508 5098
rect 21456 5034 21508 5040
rect 21468 4865 21496 5034
rect 21454 4856 21510 4865
rect 21560 4826 21588 5170
rect 21454 4791 21510 4800
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21652 4706 21680 5800
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21560 4678 21680 4706
rect 22006 4720 22062 4729
rect 21468 3534 21496 4626
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21376 2746 21496 2774
rect 21468 2038 21496 2746
rect 21560 2428 21588 4678
rect 22112 4706 22140 5102
rect 22062 4678 22140 4706
rect 22204 4690 22232 6174
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22192 4684 22244 4690
rect 22006 4655 22062 4664
rect 22192 4626 22244 4632
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21652 4282 21680 4558
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21836 4049 21864 4558
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 21638 4040 21694 4049
rect 21638 3975 21694 3984
rect 21822 4040 21878 4049
rect 21822 3975 21878 3984
rect 21652 3534 21680 3975
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 22112 3618 22140 4422
rect 22112 3590 22232 3618
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 22112 2650 22140 2926
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 21914 2544 21970 2553
rect 21914 2479 21970 2488
rect 21928 2446 21956 2479
rect 21732 2440 21784 2446
rect 21560 2400 21732 2428
rect 21732 2382 21784 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 22020 2400 22140 2428
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21456 2032 21508 2038
rect 21456 1974 21508 1980
rect 21652 1902 21680 2246
rect 22020 2106 22048 2400
rect 22112 2281 22140 2400
rect 22098 2272 22154 2281
rect 22098 2207 22154 2216
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 21640 1896 21692 1902
rect 21640 1838 21692 1844
rect 21640 1760 21692 1766
rect 21640 1702 21692 1708
rect 21652 1442 21680 1702
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 21652 1414 21772 1442
rect 21640 1352 21692 1358
rect 21638 1320 21640 1329
rect 21692 1320 21694 1329
rect 21364 1284 21416 1290
rect 21638 1255 21694 1264
rect 21364 1226 21416 1232
rect 21376 1193 21404 1226
rect 21362 1184 21418 1193
rect 21362 1119 21418 1128
rect 21744 160 21772 1414
rect 22204 1290 22232 3590
rect 22192 1284 22244 1290
rect 22192 1226 22244 1232
rect 22008 672 22060 678
rect 22008 614 22060 620
rect 22020 160 22048 614
rect 22296 160 22324 5170
rect 22388 4146 22416 6870
rect 22480 4842 22508 8214
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22572 7546 22600 7822
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22664 7410 22692 17478
rect 22756 15314 22784 18822
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22848 17202 22876 17818
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22940 16590 22968 18702
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23032 17338 23060 18566
rect 23124 18358 23152 18702
rect 23112 18352 23164 18358
rect 23112 18294 23164 18300
rect 23216 18170 23244 19366
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23308 18408 23336 19246
rect 23400 18766 23428 21830
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 20398 23520 21286
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23584 19514 23612 21490
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23676 19854 23704 21354
rect 23768 20602 23796 21422
rect 23848 21344 23900 21350
rect 23846 21312 23848 21321
rect 23900 21312 23902 21321
rect 23846 21247 23902 21256
rect 23756 20596 23808 20602
rect 23756 20538 23808 20544
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23860 19514 23888 20198
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 23848 19168 23900 19174
rect 23846 19136 23848 19145
rect 23900 19136 23902 19145
rect 23846 19071 23902 19080
rect 23480 18896 23532 18902
rect 23480 18838 23532 18844
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23308 18380 23428 18408
rect 23296 18284 23348 18290
rect 23296 18226 23348 18232
rect 23124 18142 23244 18170
rect 23124 17610 23152 18142
rect 23112 17604 23164 17610
rect 23112 17546 23164 17552
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 23308 16250 23336 18226
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 22756 15286 22876 15314
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22756 13938 22784 15098
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22848 12986 22876 15286
rect 23020 14952 23072 14958
rect 23020 14894 23072 14900
rect 22926 13968 22982 13977
rect 22926 13903 22982 13912
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11898 22784 12174
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22848 11898 22876 12038
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22940 11694 22968 13903
rect 23032 13802 23060 14894
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 23124 14074 23152 14214
rect 23308 14074 23336 14554
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 23216 13569 23244 13874
rect 23296 13728 23348 13734
rect 23294 13696 23296 13705
rect 23348 13696 23350 13705
rect 23294 13631 23350 13640
rect 23202 13560 23258 13569
rect 23202 13495 23258 13504
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11898 23152 12038
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23400 11744 23428 18380
rect 23492 16046 23520 18838
rect 23756 18692 23808 18698
rect 23756 18634 23808 18640
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23584 16590 23612 18022
rect 23768 17882 23796 18634
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 23584 15162 23612 15846
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23480 13932 23532 13938
rect 23480 13874 23532 13880
rect 23492 13530 23520 13874
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23480 13252 23532 13258
rect 23480 13194 23532 13200
rect 23492 11914 23520 13194
rect 23584 12986 23612 13806
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23676 12238 23704 16390
rect 23768 16250 23796 17818
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23860 16250 23888 17138
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 14482 23796 15302
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23860 12306 23888 15846
rect 23952 15586 23980 22066
rect 24030 20224 24086 20233
rect 24030 20159 24086 20168
rect 24044 20058 24072 20159
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24136 19446 24164 22066
rect 24228 21554 24256 26143
rect 24320 24818 24348 29514
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24412 28937 24440 28970
rect 24398 28928 24454 28937
rect 24398 28863 24454 28872
rect 24400 27872 24452 27878
rect 24398 27840 24400 27849
rect 24452 27840 24454 27849
rect 24398 27775 24454 27784
rect 24400 26784 24452 26790
rect 24398 26752 24400 26761
rect 24452 26752 24454 26761
rect 24398 26687 24454 26696
rect 24400 25696 24452 25702
rect 24398 25664 24400 25673
rect 24452 25664 24454 25673
rect 24398 25599 24454 25608
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 24400 24608 24452 24614
rect 24398 24576 24400 24585
rect 24452 24576 24454 24585
rect 24398 24511 24454 24520
rect 24400 23520 24452 23526
rect 24398 23488 24400 23497
rect 24452 23488 24454 23497
rect 24398 23423 24454 23432
rect 24504 23338 24532 36722
rect 24596 35290 24624 42094
rect 24686 41372 24994 41381
rect 24686 41370 24692 41372
rect 24748 41370 24772 41372
rect 24828 41370 24852 41372
rect 24908 41370 24932 41372
rect 24988 41370 24994 41372
rect 24748 41318 24750 41370
rect 24930 41318 24932 41370
rect 24686 41316 24692 41318
rect 24748 41316 24772 41318
rect 24828 41316 24852 41318
rect 24908 41316 24932 41318
rect 24988 41316 24994 41318
rect 24686 41307 24994 41316
rect 25056 41274 25084 44463
rect 25332 43160 25360 44463
rect 25240 43132 25360 43160
rect 25136 42764 25188 42770
rect 25136 42706 25188 42712
rect 25148 42537 25176 42706
rect 25134 42528 25190 42537
rect 25134 42463 25190 42472
rect 25136 42016 25188 42022
rect 25136 41958 25188 41964
rect 25148 41449 25176 41958
rect 25240 41750 25268 43132
rect 25318 43072 25374 43081
rect 25318 43007 25374 43016
rect 25332 41818 25360 43007
rect 25608 42362 25636 44463
rect 25596 42356 25648 42362
rect 25596 42298 25648 42304
rect 25320 41812 25372 41818
rect 25320 41754 25372 41760
rect 25228 41744 25280 41750
rect 25228 41686 25280 41692
rect 25504 41472 25556 41478
rect 25134 41440 25190 41449
rect 25504 41414 25556 41420
rect 25134 41375 25190 41384
rect 25044 41268 25096 41274
rect 25044 41210 25096 41216
rect 25136 40452 25188 40458
rect 25136 40394 25188 40400
rect 25148 40361 25176 40394
rect 25134 40352 25190 40361
rect 24686 40284 24994 40293
rect 25134 40287 25190 40296
rect 24686 40282 24692 40284
rect 24748 40282 24772 40284
rect 24828 40282 24852 40284
rect 24908 40282 24932 40284
rect 24988 40282 24994 40284
rect 24748 40230 24750 40282
rect 24930 40230 24932 40282
rect 24686 40228 24692 40230
rect 24748 40228 24772 40230
rect 24828 40228 24852 40230
rect 24908 40228 24932 40230
rect 24988 40228 24994 40230
rect 24686 40219 24994 40228
rect 25228 39296 25280 39302
rect 25226 39264 25228 39273
rect 25280 39264 25282 39273
rect 24686 39196 24994 39205
rect 25226 39199 25282 39208
rect 24686 39194 24692 39196
rect 24748 39194 24772 39196
rect 24828 39194 24852 39196
rect 24908 39194 24932 39196
rect 24988 39194 24994 39196
rect 24748 39142 24750 39194
rect 24930 39142 24932 39194
rect 24686 39140 24692 39142
rect 24748 39140 24772 39142
rect 24828 39140 24852 39142
rect 24908 39140 24932 39142
rect 24988 39140 24994 39142
rect 24686 39131 24994 39140
rect 25228 38208 25280 38214
rect 25226 38176 25228 38185
rect 25280 38176 25282 38185
rect 24686 38108 24994 38117
rect 25226 38111 25282 38120
rect 24686 38106 24692 38108
rect 24748 38106 24772 38108
rect 24828 38106 24852 38108
rect 24908 38106 24932 38108
rect 24988 38106 24994 38108
rect 24748 38054 24750 38106
rect 24930 38054 24932 38106
rect 24686 38052 24692 38054
rect 24748 38052 24772 38054
rect 24828 38052 24852 38054
rect 24908 38052 24932 38054
rect 24988 38052 24994 38054
rect 24686 38043 24994 38052
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 24686 37020 24994 37029
rect 24686 37018 24692 37020
rect 24748 37018 24772 37020
rect 24828 37018 24852 37020
rect 24908 37018 24932 37020
rect 24988 37018 24994 37020
rect 24748 36966 24750 37018
rect 24930 36966 24932 37018
rect 24686 36964 24692 36966
rect 24748 36964 24772 36966
rect 24828 36964 24852 36966
rect 24908 36964 24932 36966
rect 24988 36964 24994 36966
rect 24686 36955 24994 36964
rect 24686 35932 24994 35941
rect 24686 35930 24692 35932
rect 24748 35930 24772 35932
rect 24828 35930 24852 35932
rect 24908 35930 24932 35932
rect 24988 35930 24994 35932
rect 24748 35878 24750 35930
rect 24930 35878 24932 35930
rect 24686 35876 24692 35878
rect 24748 35876 24772 35878
rect 24828 35876 24852 35878
rect 24908 35876 24932 35878
rect 24988 35876 24994 35878
rect 24686 35867 24994 35876
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 24686 34844 24994 34853
rect 24686 34842 24692 34844
rect 24748 34842 24772 34844
rect 24828 34842 24852 34844
rect 24908 34842 24932 34844
rect 24988 34842 24994 34844
rect 24748 34790 24750 34842
rect 24930 34790 24932 34842
rect 24686 34788 24692 34790
rect 24748 34788 24772 34790
rect 24828 34788 24852 34790
rect 24908 34788 24932 34790
rect 24988 34788 24994 34790
rect 24686 34779 24994 34788
rect 24686 33756 24994 33765
rect 24686 33754 24692 33756
rect 24748 33754 24772 33756
rect 24828 33754 24852 33756
rect 24908 33754 24932 33756
rect 24988 33754 24994 33756
rect 24748 33702 24750 33754
rect 24930 33702 24932 33754
rect 24686 33700 24692 33702
rect 24748 33700 24772 33702
rect 24828 33700 24852 33702
rect 24908 33700 24932 33702
rect 24988 33700 24994 33702
rect 24686 33691 24994 33700
rect 24686 32668 24994 32677
rect 24686 32666 24692 32668
rect 24748 32666 24772 32668
rect 24828 32666 24852 32668
rect 24908 32666 24932 32668
rect 24988 32666 24994 32668
rect 24748 32614 24750 32666
rect 24930 32614 24932 32666
rect 24686 32612 24692 32614
rect 24748 32612 24772 32614
rect 24828 32612 24852 32614
rect 24908 32612 24932 32614
rect 24988 32612 24994 32614
rect 24686 32603 24994 32612
rect 24686 31580 24994 31589
rect 24686 31578 24692 31580
rect 24748 31578 24772 31580
rect 24828 31578 24852 31580
rect 24908 31578 24932 31580
rect 24988 31578 24994 31580
rect 24748 31526 24750 31578
rect 24930 31526 24932 31578
rect 24686 31524 24692 31526
rect 24748 31524 24772 31526
rect 24828 31524 24852 31526
rect 24908 31524 24932 31526
rect 24988 31524 24994 31526
rect 24686 31515 24994 31524
rect 24582 30832 24638 30841
rect 24582 30767 24638 30776
rect 24412 23310 24532 23338
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24228 20466 24256 20742
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24124 16992 24176 16998
rect 24122 16960 24124 16969
rect 24176 16960 24178 16969
rect 24122 16895 24178 16904
rect 24122 15872 24178 15881
rect 24122 15807 24178 15816
rect 24136 15706 24164 15807
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 23952 15558 24164 15586
rect 24032 14816 24084 14822
rect 24030 14784 24032 14793
rect 24084 14784 24086 14793
rect 24030 14719 24086 14728
rect 24136 12434 24164 15558
rect 24228 14414 24256 19722
rect 24320 15094 24348 20198
rect 24412 18222 24440 23310
rect 24490 22400 24546 22409
rect 24490 22335 24546 22344
rect 24504 21690 24532 22335
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24400 18216 24452 18222
rect 24400 18158 24452 18164
rect 24400 18080 24452 18086
rect 24398 18048 24400 18057
rect 24452 18048 24454 18057
rect 24398 17983 24454 17992
rect 24492 17536 24544 17542
rect 24492 17478 24544 17484
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16114 24440 16934
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24400 13728 24452 13734
rect 24398 13696 24400 13705
rect 24452 13696 24454 13705
rect 24398 13631 24454 13640
rect 24504 12918 24532 17478
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24216 12640 24268 12646
rect 24214 12608 24216 12617
rect 24268 12608 24270 12617
rect 24214 12543 24270 12552
rect 24136 12406 24440 12434
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23492 11886 23612 11914
rect 23584 11762 23612 11886
rect 23124 11716 23428 11744
rect 23480 11756 23532 11762
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22756 10674 22784 11154
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22744 10192 22796 10198
rect 22744 10134 22796 10140
rect 22756 10010 22784 10134
rect 22756 9982 22876 10010
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22756 7290 22784 9862
rect 22848 7970 22876 9982
rect 22940 8294 22968 11086
rect 23020 9920 23072 9926
rect 23020 9862 23072 9868
rect 23032 9382 23060 9862
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 23032 8090 23060 8434
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22848 7942 23060 7970
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 22664 7262 22784 7290
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22572 5545 22600 6598
rect 22664 6322 22692 7262
rect 22744 6792 22796 6798
rect 22744 6734 22796 6740
rect 22756 6458 22784 6734
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22558 5536 22614 5545
rect 22558 5471 22614 5480
rect 22848 5098 22876 7822
rect 22928 6928 22980 6934
rect 22928 6870 22980 6876
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 22480 4814 22692 4842
rect 22468 4616 22520 4622
rect 22520 4576 22600 4604
rect 22468 4558 22520 4564
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22468 4072 22520 4078
rect 22468 4014 22520 4020
rect 22374 3768 22430 3777
rect 22374 3703 22430 3712
rect 22388 2417 22416 3703
rect 22480 3398 22508 4014
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22572 3210 22600 4576
rect 22480 3182 22600 3210
rect 22374 2408 22430 2417
rect 22374 2343 22430 2352
rect 22480 2106 22508 3182
rect 22664 2774 22692 4814
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22572 2746 22692 2774
rect 22468 2100 22520 2106
rect 22468 2042 22520 2048
rect 22572 1562 22600 2746
rect 22560 1556 22612 1562
rect 22560 1498 22612 1504
rect 21454 82 21510 160
rect 21284 54 21510 82
rect 21454 0 21510 54
rect 21730 0 21786 160
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 82 22614 160
rect 22756 82 22784 4082
rect 22940 3534 22968 6870
rect 23032 5681 23060 7942
rect 23018 5672 23074 5681
rect 23018 5607 23074 5616
rect 23124 4622 23152 11716
rect 23480 11698 23532 11704
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23492 11354 23520 11698
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23584 11014 23612 11698
rect 23848 11552 23900 11558
rect 23846 11520 23848 11529
rect 23900 11520 23902 11529
rect 23846 11455 23902 11464
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 23204 10736 23256 10742
rect 23204 10678 23256 10684
rect 23216 10169 23244 10678
rect 23294 10432 23350 10441
rect 23294 10367 23350 10376
rect 23202 10160 23258 10169
rect 23202 10095 23258 10104
rect 23308 9178 23336 10367
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23296 9172 23348 9178
rect 23296 9114 23348 9120
rect 23572 8968 23624 8974
rect 23570 8936 23572 8945
rect 23624 8936 23626 8945
rect 23570 8871 23626 8880
rect 23676 8514 23704 9658
rect 23768 8634 23796 9862
rect 23848 9648 23900 9654
rect 23848 9590 23900 9596
rect 23860 9042 23888 9590
rect 24124 9376 24176 9382
rect 24030 9344 24086 9353
rect 24124 9318 24176 9324
rect 24030 9279 24086 9288
rect 24044 9178 24072 9279
rect 24136 9178 24164 9318
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23940 9036 23992 9042
rect 23940 8978 23992 8984
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23676 8486 23888 8514
rect 23480 8356 23532 8362
rect 23480 8298 23532 8304
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23216 6934 23244 8230
rect 23492 7546 23520 8298
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23492 7002 23520 7482
rect 23768 7478 23796 7754
rect 23756 7472 23808 7478
rect 23756 7414 23808 7420
rect 23754 7168 23810 7177
rect 23754 7103 23810 7112
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23204 6928 23256 6934
rect 23204 6870 23256 6876
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23202 6760 23258 6769
rect 23202 6695 23258 6704
rect 23216 5846 23244 6695
rect 23308 6322 23336 6802
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23216 4672 23244 5510
rect 23308 4826 23336 5850
rect 23296 4820 23348 4826
rect 23296 4762 23348 4768
rect 23216 4644 23336 4672
rect 23112 4616 23164 4622
rect 23112 4558 23164 4564
rect 23204 4548 23256 4554
rect 23204 4490 23256 4496
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22928 3392 22980 3398
rect 22928 3334 22980 3340
rect 22836 2916 22888 2922
rect 22836 2858 22888 2864
rect 22848 1834 22876 2858
rect 22940 2106 22968 3334
rect 23216 2650 23244 4490
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 22928 2100 22980 2106
rect 22928 2042 22980 2048
rect 23112 1964 23164 1970
rect 23112 1906 23164 1912
rect 22836 1828 22888 1834
rect 22836 1770 22888 1776
rect 22836 1420 22888 1426
rect 22836 1362 22888 1368
rect 22848 160 22876 1362
rect 23124 160 23152 1906
rect 23308 1222 23336 4644
rect 23400 3126 23428 6734
rect 23492 6202 23520 6734
rect 23572 6656 23624 6662
rect 23624 6616 23704 6644
rect 23572 6598 23624 6604
rect 23492 6174 23612 6202
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23388 3120 23440 3126
rect 23388 3062 23440 3068
rect 23492 2428 23520 6054
rect 23584 5914 23612 6174
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23584 4486 23612 5646
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23584 2582 23612 4422
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23572 2440 23624 2446
rect 23492 2400 23572 2428
rect 23676 2428 23704 6616
rect 23768 6322 23796 7103
rect 23860 6746 23888 8486
rect 23952 8430 23980 8978
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 24044 6866 24072 8434
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24320 7478 24348 8230
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 23860 6718 24164 6746
rect 24136 6338 24164 6718
rect 24228 6458 24256 7346
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 24032 6316 24084 6322
rect 24136 6310 24348 6338
rect 24032 6258 24084 6264
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23768 3670 23796 4150
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23754 3496 23810 3505
rect 23754 3431 23810 3440
rect 23768 3398 23796 3431
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23756 2440 23808 2446
rect 23676 2400 23756 2428
rect 23572 2382 23624 2388
rect 23756 2382 23808 2388
rect 23664 1896 23716 1902
rect 23664 1838 23716 1844
rect 23388 1352 23440 1358
rect 23388 1294 23440 1300
rect 23296 1216 23348 1222
rect 23296 1158 23348 1164
rect 23400 160 23428 1294
rect 23676 160 23704 1838
rect 23860 1562 23888 4490
rect 23952 2650 23980 5646
rect 24044 3194 24072 6258
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 24136 5914 24164 6054
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24228 5370 24256 6190
rect 24320 6066 24348 6310
rect 24412 6202 24440 12406
rect 24596 10198 24624 30767
rect 24686 30492 24994 30501
rect 24686 30490 24692 30492
rect 24748 30490 24772 30492
rect 24828 30490 24852 30492
rect 24908 30490 24932 30492
rect 24988 30490 24994 30492
rect 24748 30438 24750 30490
rect 24930 30438 24932 30490
rect 24686 30436 24692 30438
rect 24748 30436 24772 30438
rect 24828 30436 24852 30438
rect 24908 30436 24932 30438
rect 24988 30436 24994 30438
rect 24686 30427 24994 30436
rect 24686 29404 24994 29413
rect 24686 29402 24692 29404
rect 24748 29402 24772 29404
rect 24828 29402 24852 29404
rect 24908 29402 24932 29404
rect 24988 29402 24994 29404
rect 24748 29350 24750 29402
rect 24930 29350 24932 29402
rect 24686 29348 24692 29350
rect 24748 29348 24772 29350
rect 24828 29348 24852 29350
rect 24908 29348 24932 29350
rect 24988 29348 24994 29350
rect 24686 29339 24994 29348
rect 24686 28316 24994 28325
rect 24686 28314 24692 28316
rect 24748 28314 24772 28316
rect 24828 28314 24852 28316
rect 24908 28314 24932 28316
rect 24988 28314 24994 28316
rect 24748 28262 24750 28314
rect 24930 28262 24932 28314
rect 24686 28260 24692 28262
rect 24748 28260 24772 28262
rect 24828 28260 24852 28262
rect 24908 28260 24932 28262
rect 24988 28260 24994 28262
rect 24686 28251 24994 28260
rect 24686 27228 24994 27237
rect 24686 27226 24692 27228
rect 24748 27226 24772 27228
rect 24828 27226 24852 27228
rect 24908 27226 24932 27228
rect 24988 27226 24994 27228
rect 24748 27174 24750 27226
rect 24930 27174 24932 27226
rect 24686 27172 24692 27174
rect 24748 27172 24772 27174
rect 24828 27172 24852 27174
rect 24908 27172 24932 27174
rect 24988 27172 24994 27174
rect 24686 27163 24994 27172
rect 24686 26140 24994 26149
rect 24686 26138 24692 26140
rect 24748 26138 24772 26140
rect 24828 26138 24852 26140
rect 24908 26138 24932 26140
rect 24988 26138 24994 26140
rect 24748 26086 24750 26138
rect 24930 26086 24932 26138
rect 24686 26084 24692 26086
rect 24748 26084 24772 26086
rect 24828 26084 24852 26086
rect 24908 26084 24932 26086
rect 24988 26084 24994 26086
rect 24686 26075 24994 26084
rect 24686 25052 24994 25061
rect 24686 25050 24692 25052
rect 24748 25050 24772 25052
rect 24828 25050 24852 25052
rect 24908 25050 24932 25052
rect 24988 25050 24994 25052
rect 24748 24998 24750 25050
rect 24930 24998 24932 25050
rect 24686 24996 24692 24998
rect 24748 24996 24772 24998
rect 24828 24996 24852 24998
rect 24908 24996 24932 24998
rect 24988 24996 24994 24998
rect 24686 24987 24994 24996
rect 24686 23964 24994 23973
rect 24686 23962 24692 23964
rect 24748 23962 24772 23964
rect 24828 23962 24852 23964
rect 24908 23962 24932 23964
rect 24988 23962 24994 23964
rect 24748 23910 24750 23962
rect 24930 23910 24932 23962
rect 24686 23908 24692 23910
rect 24748 23908 24772 23910
rect 24828 23908 24852 23910
rect 24908 23908 24932 23910
rect 24988 23908 24994 23910
rect 24686 23899 24994 23908
rect 24686 22876 24994 22885
rect 24686 22874 24692 22876
rect 24748 22874 24772 22876
rect 24828 22874 24852 22876
rect 24908 22874 24932 22876
rect 24988 22874 24994 22876
rect 24748 22822 24750 22874
rect 24930 22822 24932 22874
rect 24686 22820 24692 22822
rect 24748 22820 24772 22822
rect 24828 22820 24852 22822
rect 24908 22820 24932 22822
rect 24988 22820 24994 22822
rect 24686 22811 24994 22820
rect 24686 21788 24994 21797
rect 24686 21786 24692 21788
rect 24748 21786 24772 21788
rect 24828 21786 24852 21788
rect 24908 21786 24932 21788
rect 24988 21786 24994 21788
rect 24748 21734 24750 21786
rect 24930 21734 24932 21786
rect 24686 21732 24692 21734
rect 24748 21732 24772 21734
rect 24828 21732 24852 21734
rect 24908 21732 24932 21734
rect 24988 21732 24994 21734
rect 24686 21723 24994 21732
rect 24686 20700 24994 20709
rect 24686 20698 24692 20700
rect 24748 20698 24772 20700
rect 24828 20698 24852 20700
rect 24908 20698 24932 20700
rect 24988 20698 24994 20700
rect 24748 20646 24750 20698
rect 24930 20646 24932 20698
rect 24686 20644 24692 20646
rect 24748 20644 24772 20646
rect 24828 20644 24852 20646
rect 24908 20644 24932 20646
rect 24988 20644 24994 20646
rect 24686 20635 24994 20644
rect 24686 19612 24994 19621
rect 24686 19610 24692 19612
rect 24748 19610 24772 19612
rect 24828 19610 24852 19612
rect 24908 19610 24932 19612
rect 24988 19610 24994 19612
rect 24748 19558 24750 19610
rect 24930 19558 24932 19610
rect 24686 19556 24692 19558
rect 24748 19556 24772 19558
rect 24828 19556 24852 19558
rect 24908 19556 24932 19558
rect 24988 19556 24994 19558
rect 24686 19547 24994 19556
rect 24686 18524 24994 18533
rect 24686 18522 24692 18524
rect 24748 18522 24772 18524
rect 24828 18522 24852 18524
rect 24908 18522 24932 18524
rect 24988 18522 24994 18524
rect 24748 18470 24750 18522
rect 24930 18470 24932 18522
rect 24686 18468 24692 18470
rect 24748 18468 24772 18470
rect 24828 18468 24852 18470
rect 24908 18468 24932 18470
rect 24988 18468 24994 18470
rect 24686 18459 24994 18468
rect 25056 17542 25084 37606
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 25148 36009 25176 36042
rect 25134 36000 25190 36009
rect 25134 35935 25190 35944
rect 25320 35760 25372 35766
rect 25320 35702 25372 35708
rect 25228 34944 25280 34950
rect 25226 34912 25228 34921
rect 25280 34912 25282 34921
rect 25226 34847 25282 34856
rect 25228 33856 25280 33862
rect 25226 33824 25228 33833
rect 25280 33824 25282 33833
rect 25226 33759 25282 33768
rect 25136 32836 25188 32842
rect 25136 32778 25188 32784
rect 25148 32314 25176 32778
rect 25228 32768 25280 32774
rect 25226 32736 25228 32745
rect 25280 32736 25282 32745
rect 25226 32671 25282 32680
rect 25148 32286 25268 32314
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 25148 31657 25176 31758
rect 25134 31648 25190 31657
rect 25134 31583 25190 31592
rect 25136 30660 25188 30666
rect 25136 30602 25188 30608
rect 25148 30569 25176 30602
rect 25134 30560 25190 30569
rect 25134 30495 25190 30504
rect 25136 29504 25188 29510
rect 25134 29472 25136 29481
rect 25188 29472 25190 29481
rect 25134 29407 25190 29416
rect 25136 28416 25188 28422
rect 25134 28384 25136 28393
rect 25188 28384 25190 28393
rect 25134 28319 25190 28328
rect 25136 27328 25188 27334
rect 25134 27296 25136 27305
rect 25188 27296 25190 27305
rect 25134 27231 25190 27240
rect 25240 26602 25268 32286
rect 25332 26722 25360 35702
rect 25412 33380 25464 33386
rect 25412 33322 25464 33328
rect 25320 26716 25372 26722
rect 25320 26658 25372 26664
rect 25240 26574 25360 26602
rect 25228 26512 25280 26518
rect 25228 26454 25280 26460
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25148 26217 25176 26250
rect 25134 26208 25190 26217
rect 25134 26143 25190 26152
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25148 25129 25176 25162
rect 25134 25120 25190 25129
rect 25134 25055 25190 25064
rect 25136 24064 25188 24070
rect 25134 24032 25136 24041
rect 25188 24032 25190 24041
rect 25134 23967 25190 23976
rect 25136 22976 25188 22982
rect 25134 22944 25136 22953
rect 25188 22944 25190 22953
rect 25134 22879 25190 22888
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25148 21865 25176 21898
rect 25134 21856 25190 21865
rect 25134 21791 25190 21800
rect 25134 20768 25190 20777
rect 25134 20703 25190 20712
rect 25148 19310 25176 20703
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25148 18601 25176 18838
rect 25134 18592 25190 18601
rect 25134 18527 25190 18536
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 25134 17504 25190 17513
rect 24686 17436 24994 17445
rect 25134 17439 25190 17448
rect 24686 17434 24692 17436
rect 24748 17434 24772 17436
rect 24828 17434 24852 17436
rect 24908 17434 24932 17436
rect 24988 17434 24994 17436
rect 24748 17382 24750 17434
rect 24930 17382 24932 17434
rect 24686 17380 24692 17382
rect 24748 17380 24772 17382
rect 24828 17380 24852 17382
rect 24908 17380 24932 17382
rect 24988 17380 24994 17382
rect 24686 17371 24994 17380
rect 25148 17338 25176 17439
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25240 17218 25268 26454
rect 25332 21978 25360 26574
rect 25424 22094 25452 33322
rect 25516 24177 25544 41414
rect 25780 40384 25832 40390
rect 25780 40326 25832 40332
rect 25594 38992 25650 39001
rect 25594 38927 25650 38936
rect 25502 24168 25558 24177
rect 25502 24103 25558 24112
rect 25424 22066 25544 22094
rect 25332 21950 25452 21978
rect 25318 19680 25374 19689
rect 25318 19615 25374 19624
rect 25332 18630 25360 19615
rect 25320 18624 25372 18630
rect 25320 18566 25372 18572
rect 25056 17190 25268 17218
rect 24686 16348 24994 16357
rect 24686 16346 24692 16348
rect 24748 16346 24772 16348
rect 24828 16346 24852 16348
rect 24908 16346 24932 16348
rect 24988 16346 24994 16348
rect 24748 16294 24750 16346
rect 24930 16294 24932 16346
rect 24686 16292 24692 16294
rect 24748 16292 24772 16294
rect 24828 16292 24852 16294
rect 24908 16292 24932 16294
rect 24988 16292 24994 16294
rect 24686 16283 24994 16292
rect 24686 15260 24994 15269
rect 24686 15258 24692 15260
rect 24748 15258 24772 15260
rect 24828 15258 24852 15260
rect 24908 15258 24932 15260
rect 24988 15258 24994 15260
rect 24748 15206 24750 15258
rect 24930 15206 24932 15258
rect 24686 15204 24692 15206
rect 24748 15204 24772 15206
rect 24828 15204 24852 15206
rect 24908 15204 24932 15206
rect 24988 15204 24994 15206
rect 24686 15195 24994 15204
rect 24686 14172 24994 14181
rect 24686 14170 24692 14172
rect 24748 14170 24772 14172
rect 24828 14170 24852 14172
rect 24908 14170 24932 14172
rect 24988 14170 24994 14172
rect 24748 14118 24750 14170
rect 24930 14118 24932 14170
rect 24686 14116 24692 14118
rect 24748 14116 24772 14118
rect 24828 14116 24852 14118
rect 24908 14116 24932 14118
rect 24988 14116 24994 14118
rect 24686 14107 24994 14116
rect 24686 13084 24994 13093
rect 24686 13082 24692 13084
rect 24748 13082 24772 13084
rect 24828 13082 24852 13084
rect 24908 13082 24932 13084
rect 24988 13082 24994 13084
rect 24748 13030 24750 13082
rect 24930 13030 24932 13082
rect 24686 13028 24692 13030
rect 24748 13028 24772 13030
rect 24828 13028 24852 13030
rect 24908 13028 24932 13030
rect 24988 13028 24994 13030
rect 24686 13019 24994 13028
rect 24686 11996 24994 12005
rect 24686 11994 24692 11996
rect 24748 11994 24772 11996
rect 24828 11994 24852 11996
rect 24908 11994 24932 11996
rect 24988 11994 24994 11996
rect 24748 11942 24750 11994
rect 24930 11942 24932 11994
rect 24686 11940 24692 11942
rect 24748 11940 24772 11942
rect 24828 11940 24852 11942
rect 24908 11940 24932 11942
rect 24988 11940 24994 11942
rect 24686 11931 24994 11940
rect 25056 11914 25084 17190
rect 25228 16516 25280 16522
rect 25228 16458 25280 16464
rect 25240 16425 25268 16458
rect 25226 16416 25282 16425
rect 25226 16351 25282 16360
rect 25318 15328 25374 15337
rect 25318 15263 25374 15272
rect 25136 14544 25188 14550
rect 25136 14486 25188 14492
rect 25148 14249 25176 14486
rect 25332 14278 25360 15263
rect 25320 14272 25372 14278
rect 25134 14240 25190 14249
rect 25320 14214 25372 14220
rect 25134 14175 25190 14184
rect 25320 14136 25372 14142
rect 25320 14078 25372 14084
rect 25134 12744 25190 12753
rect 25134 12679 25190 12688
rect 25148 12442 25176 12679
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25240 12073 25268 12310
rect 25226 12064 25282 12073
rect 25226 11999 25282 12008
rect 25056 11886 25176 11914
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24686 10908 24994 10917
rect 24686 10906 24692 10908
rect 24748 10906 24772 10908
rect 24828 10906 24852 10908
rect 24908 10906 24932 10908
rect 24988 10906 24994 10908
rect 24748 10854 24750 10906
rect 24930 10854 24932 10906
rect 24686 10852 24692 10854
rect 24748 10852 24772 10854
rect 24828 10852 24852 10854
rect 24908 10852 24932 10854
rect 24988 10852 24994 10854
rect 24686 10843 24994 10852
rect 24584 10192 24636 10198
rect 24584 10134 24636 10140
rect 24686 9820 24994 9829
rect 24686 9818 24692 9820
rect 24748 9818 24772 9820
rect 24828 9818 24852 9820
rect 24908 9818 24932 9820
rect 24988 9818 24994 9820
rect 24748 9766 24750 9818
rect 24930 9766 24932 9818
rect 24686 9764 24692 9766
rect 24748 9764 24772 9766
rect 24828 9764 24852 9766
rect 24908 9764 24932 9766
rect 24988 9764 24994 9766
rect 24686 9755 24994 9764
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24490 8256 24546 8265
rect 24490 8191 24546 8200
rect 24504 6322 24532 8191
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24412 6174 24532 6202
rect 24320 6038 24440 6066
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24228 4078 24256 5034
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24124 4004 24176 4010
rect 24124 3946 24176 3952
rect 24032 3188 24084 3194
rect 24032 3130 24084 3136
rect 24030 3088 24086 3097
rect 24030 3023 24086 3032
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 23848 1556 23900 1562
rect 23848 1498 23900 1504
rect 23952 1358 23980 2042
rect 23940 1352 23992 1358
rect 23940 1294 23992 1300
rect 23940 1216 23992 1222
rect 23940 1158 23992 1164
rect 23952 160 23980 1158
rect 24044 1034 24072 3023
rect 24136 1222 24164 3946
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24228 2514 24256 3606
rect 24320 3058 24348 5170
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24412 2938 24440 6038
rect 24504 4146 24532 6174
rect 24596 5098 24624 9454
rect 24686 8732 24994 8741
rect 24686 8730 24692 8732
rect 24748 8730 24772 8732
rect 24828 8730 24852 8732
rect 24908 8730 24932 8732
rect 24988 8730 24994 8732
rect 24748 8678 24750 8730
rect 24930 8678 24932 8730
rect 24686 8676 24692 8678
rect 24748 8676 24772 8678
rect 24828 8676 24852 8678
rect 24908 8676 24932 8678
rect 24988 8676 24994 8678
rect 24686 8667 24994 8676
rect 24686 7644 24994 7653
rect 24686 7642 24692 7644
rect 24748 7642 24772 7644
rect 24828 7642 24852 7644
rect 24908 7642 24932 7644
rect 24988 7642 24994 7644
rect 24748 7590 24750 7642
rect 24930 7590 24932 7642
rect 24686 7588 24692 7590
rect 24748 7588 24772 7590
rect 24828 7588 24852 7590
rect 24908 7588 24932 7590
rect 24988 7588 24994 7590
rect 24686 7579 24994 7588
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 25056 5817 25084 11698
rect 25148 11642 25176 11886
rect 25332 11762 25360 14078
rect 25320 11756 25372 11762
rect 25320 11698 25372 11704
rect 25148 11614 25360 11642
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25240 10985 25268 11494
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25136 10192 25188 10198
rect 25188 10140 25268 10146
rect 25136 10134 25268 10140
rect 25148 10118 25268 10134
rect 25134 9888 25190 9897
rect 25134 9823 25190 9832
rect 25148 7546 25176 9823
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25042 5808 25098 5817
rect 25042 5743 25098 5752
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 24584 5092 24636 5098
rect 24584 5034 24636 5040
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24584 4208 24636 4214
rect 24584 4150 24636 4156
rect 24492 4140 24544 4146
rect 24492 4082 24544 4088
rect 24320 2910 24440 2938
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24320 2038 24348 2910
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 24492 1828 24544 1834
rect 24492 1770 24544 1776
rect 24124 1216 24176 1222
rect 24124 1158 24176 1164
rect 24044 1006 24256 1034
rect 24228 160 24256 1006
rect 24504 160 24532 1770
rect 22558 54 22784 82
rect 22558 0 22614 54
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24596 82 24624 4150
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 24766 82 24822 160
rect 24596 54 24822 82
rect 24766 0 24822 54
rect 25042 82 25098 160
rect 25148 82 25176 3878
rect 25240 3777 25268 10118
rect 25226 3768 25282 3777
rect 25226 3703 25282 3712
rect 25332 1766 25360 11614
rect 25424 2990 25452 21950
rect 25516 19378 25544 22066
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25516 6905 25544 19178
rect 25502 6896 25558 6905
rect 25502 6831 25558 6840
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25412 2984 25464 2990
rect 25412 2926 25464 2932
rect 25320 1760 25372 1766
rect 25320 1702 25372 1708
rect 25320 1488 25372 1494
rect 25320 1430 25372 1436
rect 25332 160 25360 1430
rect 25516 1193 25544 4966
rect 25608 3641 25636 38927
rect 25688 30660 25740 30666
rect 25688 30602 25740 30608
rect 25700 22166 25728 30602
rect 25688 22160 25740 22166
rect 25688 22102 25740 22108
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 25700 9654 25728 21966
rect 25792 14074 25820 40326
rect 25872 24132 25924 24138
rect 25872 24074 25924 24080
rect 25884 14142 25912 24074
rect 25872 14136 25924 14142
rect 25872 14078 25924 14084
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25688 9648 25740 9654
rect 25688 9590 25740 9596
rect 25792 4826 25820 13806
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 25594 3632 25650 3641
rect 25594 3567 25650 3576
rect 25502 1184 25558 1193
rect 25502 1119 25558 1128
rect 25596 944 25648 950
rect 25596 886 25648 892
rect 25608 160 25636 886
rect 25042 54 25176 82
rect 25042 0 25098 54
rect 25318 0 25374 160
rect 25594 0 25650 160
<< via2 >>
rect 18602 44512 18658 44568
rect 478 41520 534 41576
rect 754 37848 810 37904
rect 754 34584 810 34640
rect 1030 36488 1086 36544
rect 1030 35808 1086 35864
rect 1030 33768 1086 33824
rect 2042 42336 2098 42392
rect 1214 39888 1270 39944
rect 1398 39344 1454 39400
rect 1214 38156 1216 38176
rect 1216 38156 1268 38176
rect 1268 38156 1270 38176
rect 1214 38120 1270 38156
rect 1306 36216 1362 36272
rect 1398 34992 1454 35048
rect 1306 33496 1362 33552
rect 1674 39364 1730 39400
rect 1674 39344 1676 39364
rect 1676 39344 1728 39364
rect 1728 39344 1730 39364
rect 1582 35400 1638 35456
rect 2226 41132 2282 41168
rect 2226 41112 2228 41132
rect 2228 41112 2280 41132
rect 2280 41112 2282 41132
rect 2870 41420 2872 41440
rect 2872 41420 2924 41440
rect 2924 41420 2926 41440
rect 2870 41384 2926 41420
rect 2226 39616 2282 39672
rect 2226 37712 2282 37768
rect 1674 34584 1730 34640
rect 1490 32952 1546 33008
rect 1306 32408 1362 32464
rect 1214 32136 1270 32192
rect 938 29688 994 29744
rect 2042 35572 2044 35592
rect 2044 35572 2096 35592
rect 2096 35572 2098 35592
rect 2042 35536 2098 35572
rect 3422 42064 3478 42120
rect 2778 38936 2834 38992
rect 3238 40024 3294 40080
rect 3054 38392 3110 38448
rect 2778 37188 2834 37224
rect 2778 37168 2780 37188
rect 2780 37168 2832 37188
rect 2832 37168 2834 37188
rect 2226 33632 2282 33688
rect 1398 31320 1454 31376
rect 1306 30776 1362 30832
rect 1122 29416 1178 29472
rect 1122 28736 1178 28792
rect 938 28600 994 28656
rect 754 28464 810 28520
rect 846 28056 902 28112
rect 754 27784 810 27840
rect 1306 30368 1362 30424
rect 2042 32816 2098 32872
rect 1490 29960 1546 30016
rect 1582 29724 1584 29744
rect 1584 29724 1636 29744
rect 1636 29724 1638 29744
rect 1582 29688 1638 29724
rect 1306 29144 1362 29200
rect 478 27104 534 27160
rect 478 26832 534 26888
rect 294 24112 350 24168
rect 386 23568 442 23624
rect 294 17584 350 17640
rect 846 23840 902 23896
rect 754 23432 810 23488
rect 846 20304 902 20360
rect 754 20168 810 20224
rect 846 19896 902 19952
rect 1490 28328 1546 28384
rect 1398 27648 1454 27704
rect 1306 26988 1362 27024
rect 1306 26968 1308 26988
rect 1308 26968 1360 26988
rect 1360 26968 1362 26988
rect 1214 26696 1270 26752
rect 1122 26424 1178 26480
rect 1306 25336 1362 25392
rect 1214 25064 1270 25120
rect 1122 24520 1178 24576
rect 1122 23024 1178 23080
rect 1030 22888 1086 22944
rect 1030 17312 1086 17368
rect 662 1808 718 1864
rect 938 10104 994 10160
rect 938 9560 994 9616
rect 1398 23976 1454 24032
rect 1306 23704 1362 23760
rect 1306 22652 1308 22672
rect 1308 22652 1360 22672
rect 1360 22652 1362 22672
rect 1306 22616 1362 22652
rect 1766 29416 1822 29472
rect 3146 36896 3202 36952
rect 3238 36760 3294 36816
rect 2962 35808 3018 35864
rect 2870 35672 2926 35728
rect 3238 36624 3294 36680
rect 3422 37848 3478 37904
rect 3422 37460 3478 37496
rect 3422 37440 3424 37460
rect 3424 37440 3476 37460
rect 3476 37440 3478 37460
rect 2134 31764 2136 31784
rect 2136 31764 2188 31784
rect 2188 31764 2190 31784
rect 2134 31728 2190 31764
rect 2410 32408 2466 32464
rect 2226 31456 2282 31512
rect 2226 30368 2282 30424
rect 2042 29028 2098 29064
rect 2042 29008 2044 29028
rect 2044 29008 2096 29028
rect 2096 29008 2098 29028
rect 1950 28192 2006 28248
rect 1858 28056 1914 28112
rect 1858 26424 1914 26480
rect 1858 26016 1914 26072
rect 2042 26288 2098 26344
rect 1674 24248 1730 24304
rect 1490 23160 1546 23216
rect 1306 21800 1362 21856
rect 1214 21528 1270 21584
rect 1490 22344 1546 22400
rect 1858 25200 1914 25256
rect 1858 24248 1914 24304
rect 1766 21528 1822 21584
rect 1214 21256 1270 21312
rect 1306 20984 1362 21040
rect 1306 20712 1362 20768
rect 1398 20440 1454 20496
rect 1306 19624 1362 19680
rect 2870 33224 2926 33280
rect 2778 32680 2834 32736
rect 3054 32952 3110 33008
rect 2778 31048 2834 31104
rect 2594 30676 2596 30696
rect 2596 30676 2648 30696
rect 2648 30676 2650 30696
rect 2594 30640 2650 30676
rect 3238 36216 3294 36272
rect 3422 35980 3424 36000
rect 3424 35980 3476 36000
rect 3476 35980 3478 36000
rect 3422 35944 3478 35980
rect 3923 43002 3979 43004
rect 4003 43002 4059 43004
rect 4083 43002 4139 43004
rect 4163 43002 4219 43004
rect 3923 42950 3969 43002
rect 3969 42950 3979 43002
rect 4003 42950 4033 43002
rect 4033 42950 4045 43002
rect 4045 42950 4059 43002
rect 4083 42950 4097 43002
rect 4097 42950 4109 43002
rect 4109 42950 4139 43002
rect 4163 42950 4173 43002
rect 4173 42950 4219 43002
rect 3923 42948 3979 42950
rect 4003 42948 4059 42950
rect 4083 42948 4139 42950
rect 4163 42948 4219 42950
rect 3974 42064 4030 42120
rect 3923 41914 3979 41916
rect 4003 41914 4059 41916
rect 4083 41914 4139 41916
rect 4163 41914 4219 41916
rect 3923 41862 3969 41914
rect 3969 41862 3979 41914
rect 4003 41862 4033 41914
rect 4033 41862 4045 41914
rect 4045 41862 4059 41914
rect 4083 41862 4097 41914
rect 4097 41862 4109 41914
rect 4109 41862 4139 41914
rect 4163 41862 4173 41914
rect 4173 41862 4219 41914
rect 3923 41860 3979 41862
rect 4003 41860 4059 41862
rect 4083 41860 4139 41862
rect 4163 41860 4219 41862
rect 3923 40826 3979 40828
rect 4003 40826 4059 40828
rect 4083 40826 4139 40828
rect 4163 40826 4219 40828
rect 3923 40774 3969 40826
rect 3969 40774 3979 40826
rect 4003 40774 4033 40826
rect 4033 40774 4045 40826
rect 4045 40774 4059 40826
rect 4083 40774 4097 40826
rect 4097 40774 4109 40826
rect 4109 40774 4139 40826
rect 4163 40774 4173 40826
rect 4173 40774 4219 40826
rect 3923 40772 3979 40774
rect 4003 40772 4059 40774
rect 4083 40772 4139 40774
rect 4163 40772 4219 40774
rect 4250 40296 4306 40352
rect 3923 39738 3979 39740
rect 4003 39738 4059 39740
rect 4083 39738 4139 39740
rect 4163 39738 4219 39740
rect 3923 39686 3969 39738
rect 3969 39686 3979 39738
rect 4003 39686 4033 39738
rect 4033 39686 4045 39738
rect 4045 39686 4059 39738
rect 4083 39686 4097 39738
rect 4097 39686 4109 39738
rect 4109 39686 4139 39738
rect 4163 39686 4173 39738
rect 4173 39686 4219 39738
rect 3923 39684 3979 39686
rect 4003 39684 4059 39686
rect 4083 39684 4139 39686
rect 4163 39684 4219 39686
rect 3790 39616 3846 39672
rect 3882 38836 3884 38856
rect 3884 38836 3936 38856
rect 3936 38836 3938 38856
rect 3882 38800 3938 38836
rect 3923 38650 3979 38652
rect 4003 38650 4059 38652
rect 4083 38650 4139 38652
rect 4163 38650 4219 38652
rect 3923 38598 3969 38650
rect 3969 38598 3979 38650
rect 4003 38598 4033 38650
rect 4033 38598 4045 38650
rect 4045 38598 4059 38650
rect 4083 38598 4097 38650
rect 4097 38598 4109 38650
rect 4109 38598 4139 38650
rect 4163 38598 4173 38650
rect 4173 38598 4219 38650
rect 3923 38596 3979 38598
rect 4003 38596 4059 38598
rect 4083 38596 4139 38598
rect 4163 38596 4219 38598
rect 4342 38800 4398 38856
rect 4710 42220 4766 42256
rect 4710 42200 4712 42220
rect 4712 42200 4764 42220
rect 4764 42200 4766 42220
rect 4434 38256 4490 38312
rect 3923 37562 3979 37564
rect 4003 37562 4059 37564
rect 4083 37562 4139 37564
rect 4163 37562 4219 37564
rect 3923 37510 3969 37562
rect 3969 37510 3979 37562
rect 4003 37510 4033 37562
rect 4033 37510 4045 37562
rect 4045 37510 4059 37562
rect 4083 37510 4097 37562
rect 4097 37510 4109 37562
rect 4109 37510 4139 37562
rect 4163 37510 4173 37562
rect 4173 37510 4219 37562
rect 3923 37508 3979 37510
rect 4003 37508 4059 37510
rect 4083 37508 4139 37510
rect 4163 37508 4219 37510
rect 3882 37032 3938 37088
rect 4066 36624 4122 36680
rect 3923 36474 3979 36476
rect 4003 36474 4059 36476
rect 4083 36474 4139 36476
rect 4163 36474 4219 36476
rect 3923 36422 3969 36474
rect 3969 36422 3979 36474
rect 4003 36422 4033 36474
rect 4033 36422 4045 36474
rect 4045 36422 4059 36474
rect 4083 36422 4097 36474
rect 4097 36422 4109 36474
rect 4109 36422 4139 36474
rect 4163 36422 4173 36474
rect 4173 36422 4219 36474
rect 3923 36420 3979 36422
rect 4003 36420 4059 36422
rect 4083 36420 4139 36422
rect 4163 36420 4219 36422
rect 3698 35808 3754 35864
rect 3330 34720 3386 34776
rect 3422 34040 3478 34096
rect 3606 32544 3662 32600
rect 3330 31864 3386 31920
rect 2502 28600 2558 28656
rect 2410 27920 2466 27976
rect 2318 27512 2374 27568
rect 3146 29144 3202 29200
rect 2686 27940 2742 27976
rect 2686 27920 2688 27940
rect 2688 27920 2740 27940
rect 2740 27920 2742 27940
rect 2594 27240 2650 27296
rect 2134 24792 2190 24848
rect 2594 26188 2596 26208
rect 2596 26188 2648 26208
rect 2648 26188 2650 26208
rect 2594 26152 2650 26188
rect 2686 25472 2742 25528
rect 2778 24928 2834 24984
rect 3054 28736 3110 28792
rect 3422 30504 3478 30560
rect 3422 30096 3478 30152
rect 2962 25336 3018 25392
rect 3146 24792 3202 24848
rect 2502 22888 2558 22944
rect 2870 23976 2926 24032
rect 2318 20984 2374 21040
rect 2042 20576 2098 20632
rect 2226 19896 2282 19952
rect 1582 19760 1638 19816
rect 1766 19352 1822 19408
rect 1398 18808 1454 18864
rect 1306 18264 1362 18320
rect 1214 17992 1270 18048
rect 1674 18536 1730 18592
rect 1490 18128 1546 18184
rect 1582 17856 1638 17912
rect 1490 17176 1546 17232
rect 1398 15272 1454 15328
rect 1306 13640 1362 13696
rect 1858 18536 1914 18592
rect 1766 17448 1822 17504
rect 2042 16904 2098 16960
rect 2042 16768 2098 16824
rect 2778 20440 2834 20496
rect 2318 16904 2374 16960
rect 4066 35944 4122 36000
rect 3923 35386 3979 35388
rect 4003 35386 4059 35388
rect 4083 35386 4139 35388
rect 4163 35386 4219 35388
rect 3923 35334 3969 35386
rect 3969 35334 3979 35386
rect 4003 35334 4033 35386
rect 4033 35334 4045 35386
rect 4045 35334 4059 35386
rect 4083 35334 4097 35386
rect 4097 35334 4109 35386
rect 4109 35334 4139 35386
rect 4163 35334 4173 35386
rect 4173 35334 4219 35386
rect 3923 35332 3979 35334
rect 4003 35332 4059 35334
rect 4083 35332 4139 35334
rect 4163 35332 4219 35334
rect 3790 35128 3846 35184
rect 4894 40568 4950 40624
rect 4618 38392 4674 38448
rect 4526 35572 4528 35592
rect 4528 35572 4580 35592
rect 4580 35572 4582 35592
rect 4526 35536 4582 35572
rect 4066 34448 4122 34504
rect 3923 34298 3979 34300
rect 4003 34298 4059 34300
rect 4083 34298 4139 34300
rect 4163 34298 4219 34300
rect 3923 34246 3969 34298
rect 3969 34246 3979 34298
rect 4003 34246 4033 34298
rect 4033 34246 4045 34298
rect 4045 34246 4059 34298
rect 4083 34246 4097 34298
rect 4097 34246 4109 34298
rect 4109 34246 4139 34298
rect 4163 34246 4173 34298
rect 4173 34246 4219 34298
rect 3923 34244 3979 34246
rect 4003 34244 4059 34246
rect 4083 34244 4139 34246
rect 4163 34244 4219 34246
rect 4066 33924 4122 33960
rect 4066 33904 4068 33924
rect 4068 33904 4120 33924
rect 4120 33904 4122 33924
rect 3923 33210 3979 33212
rect 4003 33210 4059 33212
rect 4083 33210 4139 33212
rect 4163 33210 4219 33212
rect 3923 33158 3969 33210
rect 3969 33158 3979 33210
rect 4003 33158 4033 33210
rect 4033 33158 4045 33210
rect 4045 33158 4059 33210
rect 4083 33158 4097 33210
rect 4097 33158 4109 33210
rect 4109 33158 4139 33210
rect 4163 33158 4173 33210
rect 4173 33158 4219 33210
rect 3923 33156 3979 33158
rect 4003 33156 4059 33158
rect 4083 33156 4139 33158
rect 4163 33156 4219 33158
rect 4066 32308 4068 32328
rect 4068 32308 4120 32328
rect 4120 32308 4122 32328
rect 4066 32272 4122 32308
rect 3923 32122 3979 32124
rect 4003 32122 4059 32124
rect 4083 32122 4139 32124
rect 4163 32122 4219 32124
rect 3923 32070 3969 32122
rect 3969 32070 3979 32122
rect 4003 32070 4033 32122
rect 4033 32070 4045 32122
rect 4045 32070 4059 32122
rect 4083 32070 4097 32122
rect 4097 32070 4109 32122
rect 4109 32070 4139 32122
rect 4163 32070 4173 32122
rect 4173 32070 4219 32122
rect 3923 32068 3979 32070
rect 4003 32068 4059 32070
rect 4083 32068 4139 32070
rect 4163 32068 4219 32070
rect 4342 33380 4398 33416
rect 4342 33360 4344 33380
rect 4344 33360 4396 33380
rect 4396 33360 4398 33380
rect 3790 31592 3846 31648
rect 4526 32680 4582 32736
rect 4158 31456 4214 31512
rect 4158 31356 4160 31376
rect 4160 31356 4212 31376
rect 4212 31356 4214 31376
rect 4158 31320 4214 31356
rect 3923 31034 3979 31036
rect 4003 31034 4059 31036
rect 4083 31034 4139 31036
rect 4163 31034 4219 31036
rect 3923 30982 3969 31034
rect 3969 30982 3979 31034
rect 4003 30982 4033 31034
rect 4033 30982 4045 31034
rect 4045 30982 4059 31034
rect 4083 30982 4097 31034
rect 4097 30982 4109 31034
rect 4109 30982 4139 31034
rect 4163 30982 4173 31034
rect 4173 30982 4219 31034
rect 3923 30980 3979 30982
rect 4003 30980 4059 30982
rect 4083 30980 4139 30982
rect 4163 30980 4219 30982
rect 3790 30232 3846 30288
rect 3606 29280 3662 29336
rect 3606 28872 3662 28928
rect 3514 25880 3570 25936
rect 3054 23160 3110 23216
rect 3238 22072 3294 22128
rect 4250 30368 4306 30424
rect 3923 29946 3979 29948
rect 4003 29946 4059 29948
rect 4083 29946 4139 29948
rect 4163 29946 4219 29948
rect 3923 29894 3969 29946
rect 3969 29894 3979 29946
rect 4003 29894 4033 29946
rect 4033 29894 4045 29946
rect 4045 29894 4059 29946
rect 4083 29894 4097 29946
rect 4097 29894 4109 29946
rect 4109 29894 4139 29946
rect 4163 29894 4173 29946
rect 4173 29894 4219 29946
rect 3923 29892 3979 29894
rect 4003 29892 4059 29894
rect 4083 29892 4139 29894
rect 4163 29892 4219 29894
rect 3882 29688 3938 29744
rect 3923 28858 3979 28860
rect 4003 28858 4059 28860
rect 4083 28858 4139 28860
rect 4163 28858 4219 28860
rect 3923 28806 3969 28858
rect 3969 28806 3979 28858
rect 4003 28806 4033 28858
rect 4033 28806 4045 28858
rect 4045 28806 4059 28858
rect 4083 28806 4097 28858
rect 4097 28806 4109 28858
rect 4109 28806 4139 28858
rect 4163 28806 4173 28858
rect 4173 28806 4219 28858
rect 3923 28804 3979 28806
rect 4003 28804 4059 28806
rect 4083 28804 4139 28806
rect 4163 28804 4219 28806
rect 3882 28212 3938 28248
rect 3882 28192 3884 28212
rect 3884 28192 3936 28212
rect 3936 28192 3938 28212
rect 3923 27770 3979 27772
rect 4003 27770 4059 27772
rect 4083 27770 4139 27772
rect 4163 27770 4219 27772
rect 3923 27718 3969 27770
rect 3969 27718 3979 27770
rect 4003 27718 4033 27770
rect 4033 27718 4045 27770
rect 4045 27718 4059 27770
rect 4083 27718 4097 27770
rect 4097 27718 4109 27770
rect 4109 27718 4139 27770
rect 4163 27718 4173 27770
rect 4173 27718 4219 27770
rect 3923 27716 3979 27718
rect 4003 27716 4059 27718
rect 4083 27716 4139 27718
rect 4163 27716 4219 27718
rect 3923 26682 3979 26684
rect 4003 26682 4059 26684
rect 4083 26682 4139 26684
rect 4163 26682 4219 26684
rect 3923 26630 3969 26682
rect 3969 26630 3979 26682
rect 4003 26630 4033 26682
rect 4033 26630 4045 26682
rect 4045 26630 4059 26682
rect 4083 26630 4097 26682
rect 4097 26630 4109 26682
rect 4109 26630 4139 26682
rect 4163 26630 4173 26682
rect 4173 26630 4219 26682
rect 3923 26628 3979 26630
rect 4003 26628 4059 26630
rect 4083 26628 4139 26630
rect 4163 26628 4219 26630
rect 3974 25916 3976 25936
rect 3976 25916 4028 25936
rect 4028 25916 4030 25936
rect 3974 25880 4030 25916
rect 4066 25744 4122 25800
rect 4618 31456 4674 31512
rect 3923 25594 3979 25596
rect 4003 25594 4059 25596
rect 4083 25594 4139 25596
rect 4163 25594 4219 25596
rect 3923 25542 3969 25594
rect 3969 25542 3979 25594
rect 4003 25542 4033 25594
rect 4033 25542 4045 25594
rect 4045 25542 4059 25594
rect 4083 25542 4097 25594
rect 4097 25542 4109 25594
rect 4109 25542 4139 25594
rect 4163 25542 4173 25594
rect 4173 25542 4219 25594
rect 3923 25540 3979 25542
rect 4003 25540 4059 25542
rect 4083 25540 4139 25542
rect 4163 25540 4219 25542
rect 3698 24656 3754 24712
rect 4158 24792 4214 24848
rect 3923 24506 3979 24508
rect 4003 24506 4059 24508
rect 4083 24506 4139 24508
rect 4163 24506 4219 24508
rect 3923 24454 3969 24506
rect 3969 24454 3979 24506
rect 4003 24454 4033 24506
rect 4033 24454 4045 24506
rect 4045 24454 4059 24506
rect 4083 24454 4097 24506
rect 4097 24454 4109 24506
rect 4109 24454 4139 24506
rect 4163 24454 4173 24506
rect 4173 24454 4219 24506
rect 3923 24452 3979 24454
rect 4003 24452 4059 24454
rect 4083 24452 4139 24454
rect 4163 24452 4219 24454
rect 4066 23860 4122 23896
rect 4066 23840 4068 23860
rect 4068 23840 4120 23860
rect 4120 23840 4122 23860
rect 3923 23418 3979 23420
rect 4003 23418 4059 23420
rect 4083 23418 4139 23420
rect 4163 23418 4219 23420
rect 3923 23366 3969 23418
rect 3969 23366 3979 23418
rect 4003 23366 4033 23418
rect 4033 23366 4045 23418
rect 4045 23366 4059 23418
rect 4083 23366 4097 23418
rect 4097 23366 4109 23418
rect 4109 23366 4139 23418
rect 4163 23366 4173 23418
rect 4173 23366 4219 23418
rect 3923 23364 3979 23366
rect 4003 23364 4059 23366
rect 4083 23364 4139 23366
rect 4163 23364 4219 23366
rect 3790 23160 3846 23216
rect 3923 22330 3979 22332
rect 4003 22330 4059 22332
rect 4083 22330 4139 22332
rect 4163 22330 4219 22332
rect 3923 22278 3969 22330
rect 3969 22278 3979 22330
rect 4003 22278 4033 22330
rect 4033 22278 4045 22330
rect 4045 22278 4059 22330
rect 4083 22278 4097 22330
rect 4097 22278 4109 22330
rect 4109 22278 4139 22330
rect 4163 22278 4173 22330
rect 4173 22278 4219 22330
rect 3923 22276 3979 22278
rect 4003 22276 4059 22278
rect 4083 22276 4139 22278
rect 4163 22276 4219 22278
rect 2870 19760 2926 19816
rect 2410 16496 2466 16552
rect 2318 15000 2374 15056
rect 1674 13912 1730 13968
rect 1858 14356 1860 14376
rect 1860 14356 1912 14376
rect 1912 14356 1914 14376
rect 1858 14320 1914 14356
rect 1490 13640 1546 13696
rect 1214 13096 1270 13152
rect 1582 12552 1638 12608
rect 1398 12008 1454 12064
rect 1766 13776 1822 13832
rect 1858 12960 1914 13016
rect 2134 12824 2190 12880
rect 1950 11464 2006 11520
rect 1398 9832 1454 9888
rect 1214 9016 1270 9072
rect 1306 8472 1362 8528
rect 1674 10376 1730 10432
rect 1582 9580 1638 9616
rect 1582 9560 1584 9580
rect 1584 9560 1636 9580
rect 1636 9560 1638 9580
rect 1490 8880 1546 8936
rect 2870 16632 2926 16688
rect 3330 19080 3386 19136
rect 4158 21936 4214 21992
rect 3923 21242 3979 21244
rect 4003 21242 4059 21244
rect 4083 21242 4139 21244
rect 4163 21242 4219 21244
rect 3923 21190 3969 21242
rect 3969 21190 3979 21242
rect 4003 21190 4033 21242
rect 4033 21190 4045 21242
rect 4045 21190 4059 21242
rect 4083 21190 4097 21242
rect 4097 21190 4109 21242
rect 4109 21190 4139 21242
rect 4163 21190 4173 21242
rect 4173 21190 4219 21242
rect 3923 21188 3979 21190
rect 4003 21188 4059 21190
rect 4083 21188 4139 21190
rect 4163 21188 4219 21190
rect 3974 20984 4030 21040
rect 3882 20460 3938 20496
rect 3882 20440 3884 20460
rect 3884 20440 3936 20460
rect 3936 20440 3938 20460
rect 3923 20154 3979 20156
rect 4003 20154 4059 20156
rect 4083 20154 4139 20156
rect 4163 20154 4219 20156
rect 3923 20102 3969 20154
rect 3969 20102 3979 20154
rect 4003 20102 4033 20154
rect 4033 20102 4045 20154
rect 4045 20102 4059 20154
rect 4083 20102 4097 20154
rect 4097 20102 4109 20154
rect 4109 20102 4139 20154
rect 4163 20102 4173 20154
rect 4173 20102 4219 20154
rect 3923 20100 3979 20102
rect 4003 20100 4059 20102
rect 4083 20100 4139 20102
rect 4163 20100 4219 20102
rect 3790 19216 3846 19272
rect 3606 17720 3662 17776
rect 3923 19066 3979 19068
rect 4003 19066 4059 19068
rect 4083 19066 4139 19068
rect 4163 19066 4219 19068
rect 3923 19014 3969 19066
rect 3969 19014 3979 19066
rect 4003 19014 4033 19066
rect 4033 19014 4045 19066
rect 4045 19014 4059 19066
rect 4083 19014 4097 19066
rect 4097 19014 4109 19066
rect 4109 19014 4139 19066
rect 4163 19014 4173 19066
rect 4173 19014 4219 19066
rect 3923 19012 3979 19014
rect 4003 19012 4059 19014
rect 4083 19012 4139 19014
rect 4163 19012 4219 19014
rect 3974 18808 4030 18864
rect 4158 18400 4214 18456
rect 4158 18284 4214 18320
rect 4158 18264 4160 18284
rect 4160 18264 4212 18284
rect 4212 18264 4214 18284
rect 3923 17978 3979 17980
rect 4003 17978 4059 17980
rect 4083 17978 4139 17980
rect 4163 17978 4219 17980
rect 3923 17926 3969 17978
rect 3969 17926 3979 17978
rect 4003 17926 4033 17978
rect 4033 17926 4045 17978
rect 4045 17926 4059 17978
rect 4083 17926 4097 17978
rect 4097 17926 4109 17978
rect 4109 17926 4139 17978
rect 4163 17926 4173 17978
rect 4173 17926 4219 17978
rect 3923 17924 3979 17926
rect 4003 17924 4059 17926
rect 4083 17924 4139 17926
rect 4163 17924 4219 17926
rect 3330 16224 3386 16280
rect 3054 16088 3110 16144
rect 3054 15544 3110 15600
rect 2778 14728 2834 14784
rect 2226 10920 2282 10976
rect 1766 8744 1822 8800
rect 2134 10124 2190 10160
rect 2134 10104 2136 10124
rect 2136 10104 2188 10124
rect 2188 10104 2190 10124
rect 1582 8200 1638 8256
rect 1398 7656 1454 7712
rect 1030 6568 1086 6624
rect 1214 6840 1270 6896
rect 1306 6296 1362 6352
rect 1306 5752 1362 5808
rect 1766 7384 1822 7440
rect 1582 5616 1638 5672
rect 846 1400 902 1456
rect 2318 9696 2374 9752
rect 2870 12144 2926 12200
rect 3054 11600 3110 11656
rect 3330 14456 3386 14512
rect 3238 12416 3294 12472
rect 3923 16890 3979 16892
rect 4003 16890 4059 16892
rect 4083 16890 4139 16892
rect 4163 16890 4219 16892
rect 3923 16838 3969 16890
rect 3969 16838 3979 16890
rect 4003 16838 4033 16890
rect 4033 16838 4045 16890
rect 4045 16838 4059 16890
rect 4083 16838 4097 16890
rect 4097 16838 4109 16890
rect 4109 16838 4139 16890
rect 4163 16838 4173 16890
rect 4173 16838 4219 16890
rect 3923 16836 3979 16838
rect 4003 16836 4059 16838
rect 4083 16836 4139 16838
rect 4163 16836 4219 16838
rect 3974 16396 3976 16416
rect 3976 16396 4028 16416
rect 4028 16396 4030 16416
rect 3974 16360 4030 16396
rect 3923 15802 3979 15804
rect 4003 15802 4059 15804
rect 4083 15802 4139 15804
rect 4163 15802 4219 15804
rect 3923 15750 3969 15802
rect 3969 15750 3979 15802
rect 4003 15750 4033 15802
rect 4033 15750 4045 15802
rect 4045 15750 4059 15802
rect 4083 15750 4097 15802
rect 4097 15750 4109 15802
rect 4109 15750 4139 15802
rect 4163 15750 4173 15802
rect 4173 15750 4219 15802
rect 3923 15748 3979 15750
rect 4003 15748 4059 15750
rect 4083 15748 4139 15750
rect 4163 15748 4219 15750
rect 3974 15544 4030 15600
rect 4158 15544 4214 15600
rect 4342 20984 4398 21040
rect 4618 21836 4620 21856
rect 4620 21836 4672 21856
rect 4672 21836 4674 21856
rect 4618 21800 4674 21836
rect 4894 34720 4950 34776
rect 6890 43546 6946 43548
rect 6970 43546 7026 43548
rect 7050 43546 7106 43548
rect 7130 43546 7186 43548
rect 6890 43494 6936 43546
rect 6936 43494 6946 43546
rect 6970 43494 7000 43546
rect 7000 43494 7012 43546
rect 7012 43494 7026 43546
rect 7050 43494 7064 43546
rect 7064 43494 7076 43546
rect 7076 43494 7106 43546
rect 7130 43494 7140 43546
rect 7140 43494 7186 43546
rect 6890 43492 6946 43494
rect 6970 43492 7026 43494
rect 7050 43492 7106 43494
rect 7130 43492 7186 43494
rect 5814 42336 5870 42392
rect 6274 41792 6330 41848
rect 6890 42458 6946 42460
rect 6970 42458 7026 42460
rect 7050 42458 7106 42460
rect 7130 42458 7186 42460
rect 6890 42406 6936 42458
rect 6936 42406 6946 42458
rect 6970 42406 7000 42458
rect 7000 42406 7012 42458
rect 7012 42406 7026 42458
rect 7050 42406 7064 42458
rect 7064 42406 7076 42458
rect 7076 42406 7106 42458
rect 7130 42406 7140 42458
rect 7140 42406 7186 42458
rect 6890 42404 6946 42406
rect 6970 42404 7026 42406
rect 7050 42404 7106 42406
rect 7130 42404 7186 42406
rect 7102 42064 7158 42120
rect 7470 41792 7526 41848
rect 5630 40568 5686 40624
rect 5354 40160 5410 40216
rect 5354 37440 5410 37496
rect 5538 37304 5594 37360
rect 5262 36760 5318 36816
rect 5446 36116 5448 36136
rect 5448 36116 5500 36136
rect 5500 36116 5502 36136
rect 5446 36080 5502 36116
rect 5354 35944 5410 36000
rect 5170 34584 5226 34640
rect 5354 34448 5410 34504
rect 5262 32952 5318 33008
rect 4986 31184 5042 31240
rect 4894 30776 4950 30832
rect 5262 30232 5318 30288
rect 5630 32272 5686 32328
rect 6890 41370 6946 41372
rect 6970 41370 7026 41372
rect 7050 41370 7106 41372
rect 7130 41370 7186 41372
rect 6890 41318 6936 41370
rect 6936 41318 6946 41370
rect 6970 41318 7000 41370
rect 7000 41318 7012 41370
rect 7012 41318 7026 41370
rect 7050 41318 7064 41370
rect 7064 41318 7076 41370
rect 7076 41318 7106 41370
rect 7130 41318 7140 41370
rect 7140 41318 7186 41370
rect 6890 41316 6946 41318
rect 6970 41316 7026 41318
rect 7050 41316 7106 41318
rect 7130 41316 7186 41318
rect 8206 41792 8262 41848
rect 8850 42608 8906 42664
rect 7286 40432 7342 40488
rect 6890 40282 6946 40284
rect 6970 40282 7026 40284
rect 7050 40282 7106 40284
rect 7130 40282 7186 40284
rect 6890 40230 6936 40282
rect 6936 40230 6946 40282
rect 6970 40230 7000 40282
rect 7000 40230 7012 40282
rect 7012 40230 7026 40282
rect 7050 40230 7064 40282
rect 7064 40230 7076 40282
rect 7076 40230 7106 40282
rect 7130 40230 7140 40282
rect 7140 40230 7186 40282
rect 6890 40228 6946 40230
rect 6970 40228 7026 40230
rect 7050 40228 7106 40230
rect 7130 40228 7186 40230
rect 6090 36488 6146 36544
rect 4986 29144 5042 29200
rect 5078 29008 5134 29064
rect 4894 28500 4896 28520
rect 4896 28500 4948 28520
rect 4948 28500 4950 28520
rect 4894 28464 4950 28500
rect 4986 27784 5042 27840
rect 4710 20984 4766 21040
rect 5170 24928 5226 24984
rect 5078 17720 5134 17776
rect 3698 14864 3754 14920
rect 3923 14714 3979 14716
rect 4003 14714 4059 14716
rect 4083 14714 4139 14716
rect 4163 14714 4219 14716
rect 3923 14662 3969 14714
rect 3969 14662 3979 14714
rect 4003 14662 4033 14714
rect 4033 14662 4045 14714
rect 4045 14662 4059 14714
rect 4083 14662 4097 14714
rect 4097 14662 4109 14714
rect 4109 14662 4139 14714
rect 4163 14662 4173 14714
rect 4173 14662 4219 14714
rect 3923 14660 3979 14662
rect 4003 14660 4059 14662
rect 4083 14660 4139 14662
rect 4163 14660 4219 14662
rect 3238 11736 3294 11792
rect 3422 11756 3478 11792
rect 3422 11736 3424 11756
rect 3424 11736 3476 11756
rect 3476 11736 3478 11756
rect 3330 11092 3332 11112
rect 3332 11092 3384 11112
rect 3384 11092 3386 11112
rect 3330 11056 3386 11092
rect 3054 10240 3110 10296
rect 2870 10004 2872 10024
rect 2872 10004 2924 10024
rect 2924 10004 2926 10024
rect 2870 9968 2926 10004
rect 2318 9288 2374 9344
rect 2686 9696 2742 9752
rect 2778 9444 2834 9480
rect 2778 9424 2780 9444
rect 2780 9424 2832 9444
rect 2832 9424 2834 9444
rect 2226 7828 2228 7848
rect 2228 7828 2280 7848
rect 2280 7828 2282 7848
rect 2226 7792 2282 7828
rect 2134 7112 2190 7168
rect 1950 5344 2006 5400
rect 2134 4936 2190 4992
rect 2594 6568 2650 6624
rect 2318 4120 2374 4176
rect 1858 2352 1914 2408
rect 2962 9696 3018 9752
rect 3146 9696 3202 9752
rect 3054 8880 3110 8936
rect 3698 12824 3754 12880
rect 4250 14456 4306 14512
rect 4342 13932 4398 13968
rect 4342 13912 4344 13932
rect 4344 13912 4396 13932
rect 4396 13912 4398 13932
rect 3923 13626 3979 13628
rect 4003 13626 4059 13628
rect 4083 13626 4139 13628
rect 4163 13626 4219 13628
rect 3923 13574 3969 13626
rect 3969 13574 3979 13626
rect 4003 13574 4033 13626
rect 4033 13574 4045 13626
rect 4045 13574 4059 13626
rect 4083 13574 4097 13626
rect 4097 13574 4109 13626
rect 4109 13574 4139 13626
rect 4163 13574 4173 13626
rect 4173 13574 4219 13626
rect 3923 13572 3979 13574
rect 4003 13572 4059 13574
rect 4083 13572 4139 13574
rect 4163 13572 4219 13574
rect 4066 13368 4122 13424
rect 3882 13232 3938 13288
rect 3923 12538 3979 12540
rect 4003 12538 4059 12540
rect 4083 12538 4139 12540
rect 4163 12538 4219 12540
rect 3923 12486 3969 12538
rect 3969 12486 3979 12538
rect 4003 12486 4033 12538
rect 4033 12486 4045 12538
rect 4045 12486 4059 12538
rect 4083 12486 4097 12538
rect 4097 12486 4109 12538
rect 4109 12486 4139 12538
rect 4163 12486 4173 12538
rect 4173 12486 4219 12538
rect 3923 12484 3979 12486
rect 4003 12484 4059 12486
rect 4083 12484 4139 12486
rect 4163 12484 4219 12486
rect 3790 12280 3846 12336
rect 3698 12008 3754 12064
rect 3606 9696 3662 9752
rect 1858 1264 1914 1320
rect 2502 1284 2558 1320
rect 2502 1264 2504 1284
rect 2504 1264 2556 1284
rect 2556 1264 2558 1284
rect 2962 6568 3018 6624
rect 2962 6432 3018 6488
rect 2962 6160 3018 6216
rect 2870 5208 2926 5264
rect 3146 4120 3202 4176
rect 3146 3052 3202 3088
rect 3146 3032 3148 3052
rect 3148 3032 3200 3052
rect 3200 3032 3202 3052
rect 3330 7928 3386 7984
rect 3974 12008 4030 12064
rect 3923 11450 3979 11452
rect 4003 11450 4059 11452
rect 4083 11450 4139 11452
rect 4163 11450 4219 11452
rect 3923 11398 3969 11450
rect 3969 11398 3979 11450
rect 4003 11398 4033 11450
rect 4033 11398 4045 11450
rect 4045 11398 4059 11450
rect 4083 11398 4097 11450
rect 4097 11398 4109 11450
rect 4109 11398 4139 11450
rect 4163 11398 4173 11450
rect 4173 11398 4219 11450
rect 3923 11396 3979 11398
rect 4003 11396 4059 11398
rect 4083 11396 4139 11398
rect 4163 11396 4219 11398
rect 3882 11192 3938 11248
rect 3422 5752 3478 5808
rect 3330 3984 3386 4040
rect 3606 6840 3662 6896
rect 3974 10648 4030 10704
rect 4066 10548 4068 10568
rect 4068 10548 4120 10568
rect 4120 10548 4122 10568
rect 4066 10512 4122 10548
rect 3923 10362 3979 10364
rect 4003 10362 4059 10364
rect 4083 10362 4139 10364
rect 4163 10362 4219 10364
rect 3923 10310 3969 10362
rect 3969 10310 3979 10362
rect 4003 10310 4033 10362
rect 4033 10310 4045 10362
rect 4045 10310 4059 10362
rect 4083 10310 4097 10362
rect 4097 10310 4109 10362
rect 4109 10310 4139 10362
rect 4163 10310 4173 10362
rect 4173 10310 4219 10362
rect 3923 10308 3979 10310
rect 4003 10308 4059 10310
rect 4083 10308 4139 10310
rect 4163 10308 4219 10310
rect 3974 10124 4030 10160
rect 3974 10104 3976 10124
rect 3976 10104 4028 10124
rect 4028 10104 4030 10124
rect 4158 10104 4214 10160
rect 4066 9968 4122 10024
rect 3923 9274 3979 9276
rect 4003 9274 4059 9276
rect 4083 9274 4139 9276
rect 4163 9274 4219 9276
rect 3923 9222 3969 9274
rect 3969 9222 3979 9274
rect 4003 9222 4033 9274
rect 4033 9222 4045 9274
rect 4045 9222 4059 9274
rect 4083 9222 4097 9274
rect 4097 9222 4109 9274
rect 4109 9222 4139 9274
rect 4163 9222 4173 9274
rect 4173 9222 4219 9274
rect 3923 9220 3979 9222
rect 4003 9220 4059 9222
rect 4083 9220 4139 9222
rect 4163 9220 4219 9222
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 5446 18536 5502 18592
rect 5078 15136 5134 15192
rect 4802 14356 4804 14376
rect 4804 14356 4856 14376
rect 4856 14356 4858 14376
rect 4802 14320 4858 14356
rect 4802 12552 4858 12608
rect 4618 12280 4674 12336
rect 4342 10920 4398 10976
rect 4342 9424 4398 9480
rect 4342 7248 4398 7304
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 4250 5072 4306 5128
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 3974 4564 3976 4584
rect 3976 4564 4028 4584
rect 4028 4564 4030 4584
rect 3974 4528 4030 4564
rect 4802 12180 4804 12200
rect 4804 12180 4856 12200
rect 4856 12180 4858 12200
rect 4802 12144 4858 12180
rect 5078 13776 5134 13832
rect 4986 12280 5042 12336
rect 4894 11636 4896 11656
rect 4896 11636 4948 11656
rect 4948 11636 4950 11656
rect 4894 11600 4950 11636
rect 5814 30368 5870 30424
rect 6182 34176 6238 34232
rect 6090 30504 6146 30560
rect 6090 29300 6146 29336
rect 6090 29280 6092 29300
rect 6092 29280 6144 29300
rect 6144 29280 6146 29300
rect 6090 27784 6146 27840
rect 6090 27512 6146 27568
rect 6090 26560 6146 26616
rect 5998 25744 6054 25800
rect 5630 21800 5686 21856
rect 5630 18420 5686 18456
rect 5630 18400 5632 18420
rect 5632 18400 5684 18420
rect 5684 18400 5686 18420
rect 5170 11192 5226 11248
rect 5078 9832 5134 9888
rect 4802 5480 4858 5536
rect 4618 5208 4674 5264
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 4526 4664 4582 4720
rect 5170 6160 5226 6216
rect 4894 4392 4950 4448
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 5630 16904 5686 16960
rect 5446 12552 5502 12608
rect 6890 39194 6946 39196
rect 6970 39194 7026 39196
rect 7050 39194 7106 39196
rect 7130 39194 7186 39196
rect 6890 39142 6936 39194
rect 6936 39142 6946 39194
rect 6970 39142 7000 39194
rect 7000 39142 7012 39194
rect 7012 39142 7026 39194
rect 7050 39142 7064 39194
rect 7064 39142 7076 39194
rect 7076 39142 7106 39194
rect 7130 39142 7140 39194
rect 7140 39142 7186 39194
rect 6890 39140 6946 39142
rect 6970 39140 7026 39142
rect 7050 39140 7106 39142
rect 7130 39140 7186 39142
rect 6890 38106 6946 38108
rect 6970 38106 7026 38108
rect 7050 38106 7106 38108
rect 7130 38106 7186 38108
rect 6890 38054 6936 38106
rect 6936 38054 6946 38106
rect 6970 38054 7000 38106
rect 7000 38054 7012 38106
rect 7012 38054 7026 38106
rect 7050 38054 7064 38106
rect 7064 38054 7076 38106
rect 7076 38054 7106 38106
rect 7130 38054 7140 38106
rect 7140 38054 7186 38106
rect 6890 38052 6946 38054
rect 6970 38052 7026 38054
rect 7050 38052 7106 38054
rect 7130 38052 7186 38054
rect 6642 37576 6698 37632
rect 6550 37032 6606 37088
rect 6890 37018 6946 37020
rect 6970 37018 7026 37020
rect 7050 37018 7106 37020
rect 7130 37018 7186 37020
rect 6890 36966 6936 37018
rect 6936 36966 6946 37018
rect 6970 36966 7000 37018
rect 7000 36966 7012 37018
rect 7012 36966 7026 37018
rect 7050 36966 7064 37018
rect 7064 36966 7076 37018
rect 7076 36966 7106 37018
rect 7130 36966 7140 37018
rect 7140 36966 7186 37018
rect 6890 36964 6946 36966
rect 6970 36964 7026 36966
rect 7050 36964 7106 36966
rect 7130 36964 7186 36966
rect 7746 40024 7802 40080
rect 7562 39480 7618 39536
rect 6366 32952 6422 33008
rect 6458 31456 6514 31512
rect 6890 35930 6946 35932
rect 6970 35930 7026 35932
rect 7050 35930 7106 35932
rect 7130 35930 7186 35932
rect 6890 35878 6936 35930
rect 6936 35878 6946 35930
rect 6970 35878 7000 35930
rect 7000 35878 7012 35930
rect 7012 35878 7026 35930
rect 7050 35878 7064 35930
rect 7064 35878 7076 35930
rect 7076 35878 7106 35930
rect 7130 35878 7140 35930
rect 7140 35878 7186 35930
rect 6890 35876 6946 35878
rect 6970 35876 7026 35878
rect 7050 35876 7106 35878
rect 7130 35876 7186 35878
rect 7654 36896 7710 36952
rect 7654 36624 7710 36680
rect 8206 38528 8262 38584
rect 6890 34842 6946 34844
rect 6970 34842 7026 34844
rect 7050 34842 7106 34844
rect 7130 34842 7186 34844
rect 6890 34790 6936 34842
rect 6936 34790 6946 34842
rect 6970 34790 7000 34842
rect 7000 34790 7012 34842
rect 7012 34790 7026 34842
rect 7050 34790 7064 34842
rect 7064 34790 7076 34842
rect 7076 34790 7106 34842
rect 7130 34790 7140 34842
rect 7140 34790 7186 34842
rect 6890 34788 6946 34790
rect 6970 34788 7026 34790
rect 7050 34788 7106 34790
rect 7130 34788 7186 34790
rect 6826 34060 6882 34096
rect 6826 34040 6828 34060
rect 6828 34040 6880 34060
rect 6880 34040 6882 34060
rect 6890 33754 6946 33756
rect 6970 33754 7026 33756
rect 7050 33754 7106 33756
rect 7130 33754 7186 33756
rect 6890 33702 6936 33754
rect 6936 33702 6946 33754
rect 6970 33702 7000 33754
rect 7000 33702 7012 33754
rect 7012 33702 7026 33754
rect 7050 33702 7064 33754
rect 7064 33702 7076 33754
rect 7076 33702 7106 33754
rect 7130 33702 7140 33754
rect 7140 33702 7186 33754
rect 6890 33700 6946 33702
rect 6970 33700 7026 33702
rect 7050 33700 7106 33702
rect 7130 33700 7186 33702
rect 7470 33496 7526 33552
rect 6918 32816 6974 32872
rect 7838 33496 7894 33552
rect 7654 32816 7710 32872
rect 7286 32680 7342 32736
rect 6890 32666 6946 32668
rect 6970 32666 7026 32668
rect 7050 32666 7106 32668
rect 7130 32666 7186 32668
rect 6890 32614 6936 32666
rect 6936 32614 6946 32666
rect 6970 32614 7000 32666
rect 7000 32614 7012 32666
rect 7012 32614 7026 32666
rect 7050 32614 7064 32666
rect 7064 32614 7076 32666
rect 7076 32614 7106 32666
rect 7130 32614 7140 32666
rect 7140 32614 7186 32666
rect 6890 32612 6946 32614
rect 6970 32612 7026 32614
rect 7050 32612 7106 32614
rect 7130 32612 7186 32614
rect 6642 31592 6698 31648
rect 6890 31578 6946 31580
rect 6970 31578 7026 31580
rect 7050 31578 7106 31580
rect 7130 31578 7186 31580
rect 6890 31526 6936 31578
rect 6936 31526 6946 31578
rect 6970 31526 7000 31578
rect 7000 31526 7012 31578
rect 7012 31526 7026 31578
rect 7050 31526 7064 31578
rect 7064 31526 7076 31578
rect 7076 31526 7106 31578
rect 7130 31526 7140 31578
rect 7140 31526 7186 31578
rect 6890 31524 6946 31526
rect 6970 31524 7026 31526
rect 7050 31524 7106 31526
rect 7130 31524 7186 31526
rect 6458 30232 6514 30288
rect 6550 29960 6606 30016
rect 6458 29416 6514 29472
rect 6890 30490 6946 30492
rect 6970 30490 7026 30492
rect 7050 30490 7106 30492
rect 7130 30490 7186 30492
rect 6890 30438 6936 30490
rect 6936 30438 6946 30490
rect 6970 30438 7000 30490
rect 7000 30438 7012 30490
rect 7012 30438 7026 30490
rect 7050 30438 7064 30490
rect 7064 30438 7076 30490
rect 7076 30438 7106 30490
rect 7130 30438 7140 30490
rect 7140 30438 7186 30490
rect 6890 30436 6946 30438
rect 6970 30436 7026 30438
rect 7050 30436 7106 30438
rect 7130 30436 7186 30438
rect 6734 30232 6790 30288
rect 7286 29416 7342 29472
rect 6890 29402 6946 29404
rect 6970 29402 7026 29404
rect 7050 29402 7106 29404
rect 7130 29402 7186 29404
rect 6890 29350 6936 29402
rect 6936 29350 6946 29402
rect 6970 29350 7000 29402
rect 7000 29350 7012 29402
rect 7012 29350 7026 29402
rect 7050 29350 7064 29402
rect 7064 29350 7076 29402
rect 7076 29350 7106 29402
rect 7130 29350 7140 29402
rect 7140 29350 7186 29402
rect 6890 29348 6946 29350
rect 6970 29348 7026 29350
rect 7050 29348 7106 29350
rect 7130 29348 7186 29350
rect 7194 28736 7250 28792
rect 6890 28314 6946 28316
rect 6970 28314 7026 28316
rect 7050 28314 7106 28316
rect 7130 28314 7186 28316
rect 6890 28262 6936 28314
rect 6936 28262 6946 28314
rect 6970 28262 7000 28314
rect 7000 28262 7012 28314
rect 7012 28262 7026 28314
rect 7050 28262 7064 28314
rect 7064 28262 7076 28314
rect 7076 28262 7106 28314
rect 7130 28262 7140 28314
rect 7140 28262 7186 28314
rect 6890 28260 6946 28262
rect 6970 28260 7026 28262
rect 7050 28260 7106 28262
rect 7130 28260 7186 28262
rect 6366 27240 6422 27296
rect 6090 23704 6146 23760
rect 5998 18672 6054 18728
rect 6090 18536 6146 18592
rect 5906 17312 5962 17368
rect 6890 27226 6946 27228
rect 6970 27226 7026 27228
rect 7050 27226 7106 27228
rect 7130 27226 7186 27228
rect 6890 27174 6936 27226
rect 6936 27174 6946 27226
rect 6970 27174 7000 27226
rect 7000 27174 7012 27226
rect 7012 27174 7026 27226
rect 7050 27174 7064 27226
rect 7064 27174 7076 27226
rect 7076 27174 7106 27226
rect 7130 27174 7140 27226
rect 7140 27174 7186 27226
rect 6890 27172 6946 27174
rect 6970 27172 7026 27174
rect 7050 27172 7106 27174
rect 7130 27172 7186 27174
rect 6826 26424 6882 26480
rect 6890 26138 6946 26140
rect 6970 26138 7026 26140
rect 7050 26138 7106 26140
rect 7130 26138 7186 26140
rect 6890 26086 6936 26138
rect 6936 26086 6946 26138
rect 6970 26086 7000 26138
rect 7000 26086 7012 26138
rect 7012 26086 7026 26138
rect 7050 26086 7064 26138
rect 7064 26086 7076 26138
rect 7076 26086 7106 26138
rect 7130 26086 7140 26138
rect 7140 26086 7186 26138
rect 6890 26084 6946 26086
rect 6970 26084 7026 26086
rect 7050 26084 7106 26086
rect 7130 26084 7186 26086
rect 6918 25336 6974 25392
rect 7286 25356 7342 25392
rect 7286 25336 7288 25356
rect 7288 25336 7340 25356
rect 7340 25336 7342 25356
rect 6890 25050 6946 25052
rect 6970 25050 7026 25052
rect 7050 25050 7106 25052
rect 7130 25050 7186 25052
rect 6890 24998 6936 25050
rect 6936 24998 6946 25050
rect 6970 24998 7000 25050
rect 7000 24998 7012 25050
rect 7012 24998 7026 25050
rect 7050 24998 7064 25050
rect 7064 24998 7076 25050
rect 7076 24998 7106 25050
rect 7130 24998 7140 25050
rect 7140 24998 7186 25050
rect 6890 24996 6946 24998
rect 6970 24996 7026 24998
rect 7050 24996 7106 24998
rect 7130 24996 7186 24998
rect 6890 23962 6946 23964
rect 6970 23962 7026 23964
rect 7050 23962 7106 23964
rect 7130 23962 7186 23964
rect 6890 23910 6936 23962
rect 6936 23910 6946 23962
rect 6970 23910 7000 23962
rect 7000 23910 7012 23962
rect 7012 23910 7026 23962
rect 7050 23910 7064 23962
rect 7064 23910 7076 23962
rect 7076 23910 7106 23962
rect 7130 23910 7140 23962
rect 7140 23910 7186 23962
rect 6890 23908 6946 23910
rect 6970 23908 7026 23910
rect 7050 23908 7106 23910
rect 7130 23908 7186 23910
rect 6366 20576 6422 20632
rect 6366 20168 6422 20224
rect 6550 22752 6606 22808
rect 6890 22874 6946 22876
rect 6970 22874 7026 22876
rect 7050 22874 7106 22876
rect 7130 22874 7186 22876
rect 6890 22822 6936 22874
rect 6936 22822 6946 22874
rect 6970 22822 7000 22874
rect 7000 22822 7012 22874
rect 7012 22822 7026 22874
rect 7050 22822 7064 22874
rect 7064 22822 7076 22874
rect 7076 22822 7106 22874
rect 7130 22822 7140 22874
rect 7140 22822 7186 22874
rect 6890 22820 6946 22822
rect 6970 22820 7026 22822
rect 7050 22820 7106 22822
rect 7130 22820 7186 22822
rect 7470 29688 7526 29744
rect 7838 30504 7894 30560
rect 8114 30368 8170 30424
rect 6890 21786 6946 21788
rect 6970 21786 7026 21788
rect 7050 21786 7106 21788
rect 7130 21786 7186 21788
rect 6890 21734 6936 21786
rect 6936 21734 6946 21786
rect 6970 21734 7000 21786
rect 7000 21734 7012 21786
rect 7012 21734 7026 21786
rect 7050 21734 7064 21786
rect 7064 21734 7076 21786
rect 7076 21734 7106 21786
rect 7130 21734 7140 21786
rect 7140 21734 7186 21786
rect 6890 21732 6946 21734
rect 6970 21732 7026 21734
rect 7050 21732 7106 21734
rect 7130 21732 7186 21734
rect 6550 20712 6606 20768
rect 6458 18944 6514 19000
rect 5722 12280 5778 12336
rect 5722 7656 5778 7712
rect 5722 6452 5778 6488
rect 5722 6432 5724 6452
rect 5724 6432 5776 6452
rect 5776 6432 5778 6452
rect 6458 14320 6514 14376
rect 6274 12280 6330 12336
rect 5998 9968 6054 10024
rect 5446 5616 5502 5672
rect 6366 12144 6422 12200
rect 6458 9968 6514 10024
rect 6090 7268 6146 7304
rect 6090 7248 6092 7268
rect 6092 7248 6144 7268
rect 6144 7248 6146 7268
rect 6890 20698 6946 20700
rect 6970 20698 7026 20700
rect 7050 20698 7106 20700
rect 7130 20698 7186 20700
rect 6890 20646 6936 20698
rect 6936 20646 6946 20698
rect 6970 20646 7000 20698
rect 7000 20646 7012 20698
rect 7012 20646 7026 20698
rect 7050 20646 7064 20698
rect 7064 20646 7076 20698
rect 7076 20646 7106 20698
rect 7130 20646 7140 20698
rect 7140 20646 7186 20698
rect 6890 20644 6946 20646
rect 6970 20644 7026 20646
rect 7050 20644 7106 20646
rect 7130 20644 7186 20646
rect 6826 19780 6882 19816
rect 7562 27648 7618 27704
rect 7654 26832 7710 26888
rect 7654 21564 7656 21584
rect 7656 21564 7708 21584
rect 7708 21564 7710 21584
rect 7654 21528 7710 21564
rect 7562 20712 7618 20768
rect 6826 19760 6828 19780
rect 6828 19760 6880 19780
rect 6880 19760 6882 19780
rect 6890 19610 6946 19612
rect 6970 19610 7026 19612
rect 7050 19610 7106 19612
rect 7130 19610 7186 19612
rect 6890 19558 6936 19610
rect 6936 19558 6946 19610
rect 6970 19558 7000 19610
rect 7000 19558 7012 19610
rect 7012 19558 7026 19610
rect 7050 19558 7064 19610
rect 7064 19558 7076 19610
rect 7076 19558 7106 19610
rect 7130 19558 7140 19610
rect 7140 19558 7186 19610
rect 6890 19556 6946 19558
rect 6970 19556 7026 19558
rect 7050 19556 7106 19558
rect 7130 19556 7186 19558
rect 7194 19372 7250 19408
rect 7194 19352 7196 19372
rect 7196 19352 7248 19372
rect 7248 19352 7250 19372
rect 7470 19760 7526 19816
rect 6890 18522 6946 18524
rect 6970 18522 7026 18524
rect 7050 18522 7106 18524
rect 7130 18522 7186 18524
rect 6890 18470 6936 18522
rect 6936 18470 6946 18522
rect 6970 18470 7000 18522
rect 7000 18470 7012 18522
rect 7012 18470 7026 18522
rect 7050 18470 7064 18522
rect 7064 18470 7076 18522
rect 7076 18470 7106 18522
rect 7130 18470 7140 18522
rect 7140 18470 7186 18522
rect 6890 18468 6946 18470
rect 6970 18468 7026 18470
rect 7050 18468 7106 18470
rect 7130 18468 7186 18470
rect 6918 18128 6974 18184
rect 7286 17584 7342 17640
rect 6890 17434 6946 17436
rect 6970 17434 7026 17436
rect 7050 17434 7106 17436
rect 7130 17434 7186 17436
rect 6890 17382 6936 17434
rect 6936 17382 6946 17434
rect 6970 17382 7000 17434
rect 7000 17382 7012 17434
rect 7012 17382 7026 17434
rect 7050 17382 7064 17434
rect 7064 17382 7076 17434
rect 7076 17382 7106 17434
rect 7130 17382 7140 17434
rect 7140 17382 7186 17434
rect 6890 17380 6946 17382
rect 6970 17380 7026 17382
rect 7050 17380 7106 17382
rect 7130 17380 7186 17382
rect 6642 17212 6644 17232
rect 6644 17212 6696 17232
rect 6696 17212 6698 17232
rect 6642 17176 6698 17212
rect 6826 17040 6882 17096
rect 7194 16904 7250 16960
rect 8206 29280 8262 29336
rect 8298 24248 8354 24304
rect 8574 32544 8630 32600
rect 8482 31728 8538 31784
rect 8482 25880 8538 25936
rect 7930 22888 7986 22944
rect 8022 20712 8078 20768
rect 7930 18400 7986 18456
rect 7838 17992 7894 18048
rect 6826 16668 6828 16688
rect 6828 16668 6880 16688
rect 6880 16668 6882 16688
rect 6826 16632 6882 16668
rect 6642 15000 6698 15056
rect 6890 16346 6946 16348
rect 6970 16346 7026 16348
rect 7050 16346 7106 16348
rect 7130 16346 7186 16348
rect 6890 16294 6936 16346
rect 6936 16294 6946 16346
rect 6970 16294 7000 16346
rect 7000 16294 7012 16346
rect 7012 16294 7026 16346
rect 7050 16294 7064 16346
rect 7064 16294 7076 16346
rect 7076 16294 7106 16346
rect 7130 16294 7140 16346
rect 7140 16294 7186 16346
rect 6890 16292 6946 16294
rect 6970 16292 7026 16294
rect 7050 16292 7106 16294
rect 7130 16292 7186 16294
rect 6890 15258 6946 15260
rect 6970 15258 7026 15260
rect 7050 15258 7106 15260
rect 7130 15258 7186 15260
rect 6890 15206 6936 15258
rect 6936 15206 6946 15258
rect 6970 15206 7000 15258
rect 7000 15206 7012 15258
rect 7012 15206 7026 15258
rect 7050 15206 7064 15258
rect 7064 15206 7076 15258
rect 7076 15206 7106 15258
rect 7130 15206 7140 15258
rect 7140 15206 7186 15258
rect 6890 15204 6946 15206
rect 6970 15204 7026 15206
rect 7050 15204 7106 15206
rect 7130 15204 7186 15206
rect 6918 14320 6974 14376
rect 6890 14170 6946 14172
rect 6970 14170 7026 14172
rect 7050 14170 7106 14172
rect 7130 14170 7186 14172
rect 6890 14118 6936 14170
rect 6936 14118 6946 14170
rect 6970 14118 7000 14170
rect 7000 14118 7012 14170
rect 7012 14118 7026 14170
rect 7050 14118 7064 14170
rect 7064 14118 7076 14170
rect 7076 14118 7106 14170
rect 7130 14118 7140 14170
rect 7140 14118 7186 14170
rect 6890 14116 6946 14118
rect 6970 14116 7026 14118
rect 7050 14116 7106 14118
rect 7130 14116 7186 14118
rect 7378 13912 7434 13968
rect 6890 13082 6946 13084
rect 6970 13082 7026 13084
rect 7050 13082 7106 13084
rect 7130 13082 7186 13084
rect 6890 13030 6936 13082
rect 6936 13030 6946 13082
rect 6970 13030 7000 13082
rect 7000 13030 7012 13082
rect 7012 13030 7026 13082
rect 7050 13030 7064 13082
rect 7064 13030 7076 13082
rect 7076 13030 7106 13082
rect 7130 13030 7140 13082
rect 7140 13030 7186 13082
rect 6890 13028 6946 13030
rect 6970 13028 7026 13030
rect 7050 13028 7106 13030
rect 7130 13028 7186 13030
rect 6826 12416 6882 12472
rect 7102 12416 7158 12472
rect 6890 11994 6946 11996
rect 6970 11994 7026 11996
rect 7050 11994 7106 11996
rect 7130 11994 7186 11996
rect 6890 11942 6936 11994
rect 6936 11942 6946 11994
rect 6970 11942 7000 11994
rect 7000 11942 7012 11994
rect 7012 11942 7026 11994
rect 7050 11942 7064 11994
rect 7064 11942 7076 11994
rect 7076 11942 7106 11994
rect 7130 11942 7140 11994
rect 7140 11942 7186 11994
rect 6890 11940 6946 11942
rect 6970 11940 7026 11942
rect 7050 11940 7106 11942
rect 7130 11940 7186 11942
rect 7378 12552 7434 12608
rect 7378 12144 7434 12200
rect 6890 10906 6946 10908
rect 6970 10906 7026 10908
rect 7050 10906 7106 10908
rect 7130 10906 7186 10908
rect 6890 10854 6936 10906
rect 6936 10854 6946 10906
rect 6970 10854 7000 10906
rect 7000 10854 7012 10906
rect 7012 10854 7026 10906
rect 7050 10854 7064 10906
rect 7064 10854 7076 10906
rect 7076 10854 7106 10906
rect 7130 10854 7140 10906
rect 7140 10854 7186 10906
rect 6890 10852 6946 10854
rect 6970 10852 7026 10854
rect 7050 10852 7106 10854
rect 7130 10852 7186 10854
rect 6890 9818 6946 9820
rect 6970 9818 7026 9820
rect 7050 9818 7106 9820
rect 7130 9818 7186 9820
rect 6890 9766 6936 9818
rect 6936 9766 6946 9818
rect 6970 9766 7000 9818
rect 7000 9766 7012 9818
rect 7012 9766 7026 9818
rect 7050 9766 7064 9818
rect 7064 9766 7076 9818
rect 7076 9766 7106 9818
rect 7130 9766 7140 9818
rect 7140 9766 7186 9818
rect 6890 9764 6946 9766
rect 6970 9764 7026 9766
rect 7050 9764 7106 9766
rect 7130 9764 7186 9766
rect 6890 8730 6946 8732
rect 6970 8730 7026 8732
rect 7050 8730 7106 8732
rect 7130 8730 7186 8732
rect 6890 8678 6936 8730
rect 6936 8678 6946 8730
rect 6970 8678 7000 8730
rect 7000 8678 7012 8730
rect 7012 8678 7026 8730
rect 7050 8678 7064 8730
rect 7064 8678 7076 8730
rect 7076 8678 7106 8730
rect 7130 8678 7140 8730
rect 7140 8678 7186 8730
rect 6890 8676 6946 8678
rect 6970 8676 7026 8678
rect 7050 8676 7106 8678
rect 7130 8676 7186 8678
rect 7194 7948 7250 7984
rect 7194 7928 7196 7948
rect 7196 7928 7248 7948
rect 7248 7928 7250 7948
rect 6890 7642 6946 7644
rect 6970 7642 7026 7644
rect 7050 7642 7106 7644
rect 7130 7642 7186 7644
rect 6890 7590 6936 7642
rect 6936 7590 6946 7642
rect 6970 7590 7000 7642
rect 7000 7590 7012 7642
rect 7012 7590 7026 7642
rect 7050 7590 7064 7642
rect 7064 7590 7076 7642
rect 7076 7590 7106 7642
rect 7130 7590 7140 7642
rect 7140 7590 7186 7642
rect 6890 7588 6946 7590
rect 6970 7588 7026 7590
rect 7050 7588 7106 7590
rect 7130 7588 7186 7590
rect 6366 3732 6422 3768
rect 6366 3712 6368 3732
rect 6368 3712 6420 3732
rect 6420 3712 6422 3732
rect 6182 3440 6238 3496
rect 3974 2216 4030 2272
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 4894 2624 4950 2680
rect 6274 2760 6330 2816
rect 6182 2488 6238 2544
rect 4986 2100 5042 2136
rect 4986 2080 4988 2100
rect 4988 2080 5040 2100
rect 5040 2080 5042 2100
rect 5078 1708 5080 1728
rect 5080 1708 5132 1728
rect 5132 1708 5134 1728
rect 5078 1672 5134 1708
rect 5078 1164 5080 1184
rect 5080 1164 5132 1184
rect 5132 1164 5134 1184
rect 5078 1128 5134 1164
rect 5814 2216 5870 2272
rect 6550 2896 6606 2952
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 6826 2896 6882 2952
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 5538 1300 5540 1320
rect 5540 1300 5592 1320
rect 5592 1300 5594 1320
rect 5538 1264 5594 1300
rect 7838 14864 7894 14920
rect 8850 35536 8906 35592
rect 8942 35128 8998 35184
rect 8850 34176 8906 34232
rect 8850 33904 8906 33960
rect 8758 29280 8814 29336
rect 8758 29008 8814 29064
rect 8206 21392 8262 21448
rect 8206 19896 8262 19952
rect 8390 18808 8446 18864
rect 8850 28056 8906 28112
rect 9494 42220 9550 42256
rect 9494 42200 9496 42220
rect 9496 42200 9548 42220
rect 9548 42200 9550 42220
rect 9857 43002 9913 43004
rect 9937 43002 9993 43004
rect 10017 43002 10073 43004
rect 10097 43002 10153 43004
rect 9857 42950 9903 43002
rect 9903 42950 9913 43002
rect 9937 42950 9967 43002
rect 9967 42950 9979 43002
rect 9979 42950 9993 43002
rect 10017 42950 10031 43002
rect 10031 42950 10043 43002
rect 10043 42950 10073 43002
rect 10097 42950 10107 43002
rect 10107 42950 10153 43002
rect 9857 42948 9913 42950
rect 9937 42948 9993 42950
rect 10017 42948 10073 42950
rect 10097 42948 10153 42950
rect 9862 42200 9918 42256
rect 9857 41914 9913 41916
rect 9937 41914 9993 41916
rect 10017 41914 10073 41916
rect 10097 41914 10153 41916
rect 9857 41862 9903 41914
rect 9903 41862 9913 41914
rect 9937 41862 9967 41914
rect 9967 41862 9979 41914
rect 9979 41862 9993 41914
rect 10017 41862 10031 41914
rect 10031 41862 10043 41914
rect 10043 41862 10073 41914
rect 10097 41862 10107 41914
rect 10107 41862 10153 41914
rect 9857 41860 9913 41862
rect 9937 41860 9993 41862
rect 10017 41860 10073 41862
rect 10097 41860 10153 41862
rect 9586 41520 9642 41576
rect 9770 41520 9826 41576
rect 9494 40568 9550 40624
rect 9857 40826 9913 40828
rect 9937 40826 9993 40828
rect 10017 40826 10073 40828
rect 10097 40826 10153 40828
rect 9857 40774 9903 40826
rect 9903 40774 9913 40826
rect 9937 40774 9967 40826
rect 9967 40774 9979 40826
rect 9979 40774 9993 40826
rect 10017 40774 10031 40826
rect 10031 40774 10043 40826
rect 10043 40774 10073 40826
rect 10097 40774 10107 40826
rect 10107 40774 10153 40826
rect 9857 40772 9913 40774
rect 9937 40772 9993 40774
rect 10017 40772 10073 40774
rect 10097 40772 10153 40774
rect 9126 36780 9182 36816
rect 9126 36760 9128 36780
rect 9128 36760 9180 36780
rect 9180 36760 9182 36780
rect 9857 39738 9913 39740
rect 9937 39738 9993 39740
rect 10017 39738 10073 39740
rect 10097 39738 10153 39740
rect 9857 39686 9903 39738
rect 9903 39686 9913 39738
rect 9937 39686 9967 39738
rect 9967 39686 9979 39738
rect 9979 39686 9993 39738
rect 10017 39686 10031 39738
rect 10031 39686 10043 39738
rect 10043 39686 10073 39738
rect 10097 39686 10107 39738
rect 10107 39686 10153 39738
rect 9857 39684 9913 39686
rect 9937 39684 9993 39686
rect 10017 39684 10073 39686
rect 10097 39684 10153 39686
rect 9678 38528 9734 38584
rect 9402 36216 9458 36272
rect 9402 35708 9404 35728
rect 9404 35708 9456 35728
rect 9456 35708 9458 35728
rect 9402 35672 9458 35708
rect 9034 34176 9090 34232
rect 9857 38650 9913 38652
rect 9937 38650 9993 38652
rect 10017 38650 10073 38652
rect 10097 38650 10153 38652
rect 9857 38598 9903 38650
rect 9903 38598 9913 38650
rect 9937 38598 9967 38650
rect 9967 38598 9979 38650
rect 9979 38598 9993 38650
rect 10017 38598 10031 38650
rect 10031 38598 10043 38650
rect 10043 38598 10073 38650
rect 10097 38598 10107 38650
rect 10107 38598 10153 38650
rect 9857 38596 9913 38598
rect 9937 38596 9993 38598
rect 10017 38596 10073 38598
rect 10097 38596 10153 38598
rect 9857 37562 9913 37564
rect 9937 37562 9993 37564
rect 10017 37562 10073 37564
rect 10097 37562 10153 37564
rect 9857 37510 9903 37562
rect 9903 37510 9913 37562
rect 9937 37510 9967 37562
rect 9967 37510 9979 37562
rect 9979 37510 9993 37562
rect 10017 37510 10031 37562
rect 10031 37510 10043 37562
rect 10043 37510 10073 37562
rect 10097 37510 10107 37562
rect 10107 37510 10153 37562
rect 9857 37508 9913 37510
rect 9937 37508 9993 37510
rect 10017 37508 10073 37510
rect 10097 37508 10153 37510
rect 9857 36474 9913 36476
rect 9937 36474 9993 36476
rect 10017 36474 10073 36476
rect 10097 36474 10153 36476
rect 9857 36422 9903 36474
rect 9903 36422 9913 36474
rect 9937 36422 9967 36474
rect 9967 36422 9979 36474
rect 9979 36422 9993 36474
rect 10017 36422 10031 36474
rect 10031 36422 10043 36474
rect 10043 36422 10073 36474
rect 10097 36422 10107 36474
rect 10107 36422 10153 36474
rect 9857 36420 9913 36422
rect 9937 36420 9993 36422
rect 10017 36420 10073 36422
rect 10097 36420 10153 36422
rect 9857 35386 9913 35388
rect 9937 35386 9993 35388
rect 10017 35386 10073 35388
rect 10097 35386 10153 35388
rect 9857 35334 9903 35386
rect 9903 35334 9913 35386
rect 9937 35334 9967 35386
rect 9967 35334 9979 35386
rect 9979 35334 9993 35386
rect 10017 35334 10031 35386
rect 10031 35334 10043 35386
rect 10043 35334 10073 35386
rect 10097 35334 10107 35386
rect 10107 35334 10153 35386
rect 9857 35332 9913 35334
rect 9937 35332 9993 35334
rect 10017 35332 10073 35334
rect 10097 35332 10153 35334
rect 9494 34176 9550 34232
rect 9402 33904 9458 33960
rect 9857 34298 9913 34300
rect 9937 34298 9993 34300
rect 10017 34298 10073 34300
rect 10097 34298 10153 34300
rect 9857 34246 9903 34298
rect 9903 34246 9913 34298
rect 9937 34246 9967 34298
rect 9967 34246 9979 34298
rect 9979 34246 9993 34298
rect 10017 34246 10031 34298
rect 10031 34246 10043 34298
rect 10043 34246 10073 34298
rect 10097 34246 10107 34298
rect 10107 34246 10153 34298
rect 9857 34244 9913 34246
rect 9937 34244 9993 34246
rect 10017 34244 10073 34246
rect 10097 34244 10153 34246
rect 9770 33516 9826 33552
rect 9770 33496 9772 33516
rect 9772 33496 9824 33516
rect 9824 33496 9826 33516
rect 9857 33210 9913 33212
rect 9937 33210 9993 33212
rect 10017 33210 10073 33212
rect 10097 33210 10153 33212
rect 9857 33158 9903 33210
rect 9903 33158 9913 33210
rect 9937 33158 9967 33210
rect 9967 33158 9979 33210
rect 9979 33158 9993 33210
rect 10017 33158 10031 33210
rect 10031 33158 10043 33210
rect 10043 33158 10073 33210
rect 10097 33158 10107 33210
rect 10107 33158 10153 33210
rect 9857 33156 9913 33158
rect 9937 33156 9993 33158
rect 10017 33156 10073 33158
rect 10097 33156 10153 33158
rect 9494 32544 9550 32600
rect 9218 30676 9220 30696
rect 9220 30676 9272 30696
rect 9272 30676 9274 30696
rect 9218 30640 9274 30676
rect 9402 30368 9458 30424
rect 9678 31900 9680 31920
rect 9680 31900 9732 31920
rect 9732 31900 9734 31920
rect 9678 31864 9734 31900
rect 9857 32122 9913 32124
rect 9937 32122 9993 32124
rect 10017 32122 10073 32124
rect 10097 32122 10153 32124
rect 9857 32070 9903 32122
rect 9903 32070 9913 32122
rect 9937 32070 9967 32122
rect 9967 32070 9979 32122
rect 9979 32070 9993 32122
rect 10017 32070 10031 32122
rect 10031 32070 10043 32122
rect 10043 32070 10073 32122
rect 10097 32070 10107 32122
rect 10107 32070 10153 32122
rect 9857 32068 9913 32070
rect 9937 32068 9993 32070
rect 10017 32068 10073 32070
rect 10097 32068 10153 32070
rect 9770 31184 9826 31240
rect 9857 31034 9913 31036
rect 9937 31034 9993 31036
rect 10017 31034 10073 31036
rect 10097 31034 10153 31036
rect 9857 30982 9903 31034
rect 9903 30982 9913 31034
rect 9937 30982 9967 31034
rect 9967 30982 9979 31034
rect 9979 30982 9993 31034
rect 10017 30982 10031 31034
rect 10031 30982 10043 31034
rect 10043 30982 10073 31034
rect 10097 30982 10107 31034
rect 10107 30982 10153 31034
rect 9857 30980 9913 30982
rect 9937 30980 9993 30982
rect 10017 30980 10073 30982
rect 10097 30980 10153 30982
rect 10138 30776 10194 30832
rect 9586 30368 9642 30424
rect 9494 29688 9550 29744
rect 8758 23568 8814 23624
rect 7930 12688 7986 12744
rect 8022 12280 8078 12336
rect 8022 11600 8078 11656
rect 7838 9424 7894 9480
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 8482 13640 8538 13696
rect 8390 12824 8446 12880
rect 8482 12416 8538 12472
rect 8666 16652 8722 16688
rect 8666 16632 8668 16652
rect 8668 16632 8720 16652
rect 8720 16632 8722 16652
rect 8114 7928 8170 7984
rect 8022 4548 8078 4584
rect 8022 4528 8024 4548
rect 8024 4528 8076 4548
rect 8076 4528 8078 4548
rect 8114 2624 8170 2680
rect 7562 856 7618 912
rect 7930 2216 7986 2272
rect 8022 1944 8078 2000
rect 9126 21664 9182 21720
rect 8850 20168 8906 20224
rect 8942 18944 8998 19000
rect 9586 29008 9642 29064
rect 9494 28464 9550 28520
rect 9857 29946 9913 29948
rect 9937 29946 9993 29948
rect 10017 29946 10073 29948
rect 10097 29946 10153 29948
rect 9857 29894 9903 29946
rect 9903 29894 9913 29946
rect 9937 29894 9967 29946
rect 9967 29894 9979 29946
rect 9979 29894 9993 29946
rect 10017 29894 10031 29946
rect 10031 29894 10043 29946
rect 10043 29894 10073 29946
rect 10097 29894 10107 29946
rect 10107 29894 10153 29946
rect 9857 29892 9913 29894
rect 9937 29892 9993 29894
rect 10017 29892 10073 29894
rect 10097 29892 10153 29894
rect 10138 29280 10194 29336
rect 10322 42064 10378 42120
rect 10414 40976 10470 41032
rect 10782 38800 10838 38856
rect 10322 35672 10378 35728
rect 10598 36216 10654 36272
rect 10782 34176 10838 34232
rect 10506 31048 10562 31104
rect 10782 30776 10838 30832
rect 10598 30640 10654 30696
rect 9857 28858 9913 28860
rect 9937 28858 9993 28860
rect 10017 28858 10073 28860
rect 10097 28858 10153 28860
rect 9857 28806 9903 28858
rect 9903 28806 9913 28858
rect 9937 28806 9967 28858
rect 9967 28806 9979 28858
rect 9979 28806 9993 28858
rect 10017 28806 10031 28858
rect 10031 28806 10043 28858
rect 10043 28806 10073 28858
rect 10097 28806 10107 28858
rect 10107 28806 10153 28858
rect 9857 28804 9913 28806
rect 9937 28804 9993 28806
rect 10017 28804 10073 28806
rect 10097 28804 10153 28806
rect 9586 26560 9642 26616
rect 10046 28192 10102 28248
rect 9857 27770 9913 27772
rect 9937 27770 9993 27772
rect 10017 27770 10073 27772
rect 10097 27770 10153 27772
rect 9857 27718 9903 27770
rect 9903 27718 9913 27770
rect 9937 27718 9967 27770
rect 9967 27718 9979 27770
rect 9979 27718 9993 27770
rect 10017 27718 10031 27770
rect 10031 27718 10043 27770
rect 10043 27718 10073 27770
rect 10097 27718 10107 27770
rect 10107 27718 10153 27770
rect 9857 27716 9913 27718
rect 9937 27716 9993 27718
rect 10017 27716 10073 27718
rect 10097 27716 10153 27718
rect 9954 26968 10010 27024
rect 9857 26682 9913 26684
rect 9937 26682 9993 26684
rect 10017 26682 10073 26684
rect 10097 26682 10153 26684
rect 9857 26630 9903 26682
rect 9903 26630 9913 26682
rect 9937 26630 9967 26682
rect 9967 26630 9979 26682
rect 9979 26630 9993 26682
rect 10017 26630 10031 26682
rect 10031 26630 10043 26682
rect 10043 26630 10073 26682
rect 10097 26630 10107 26682
rect 10107 26630 10153 26682
rect 9857 26628 9913 26630
rect 9937 26628 9993 26630
rect 10017 26628 10073 26630
rect 10097 26628 10153 26630
rect 10138 26424 10194 26480
rect 9586 23976 9642 24032
rect 9586 22616 9642 22672
rect 9857 25594 9913 25596
rect 9937 25594 9993 25596
rect 10017 25594 10073 25596
rect 10097 25594 10153 25596
rect 9857 25542 9903 25594
rect 9903 25542 9913 25594
rect 9937 25542 9967 25594
rect 9967 25542 9979 25594
rect 9979 25542 9993 25594
rect 10017 25542 10031 25594
rect 10031 25542 10043 25594
rect 10043 25542 10073 25594
rect 10097 25542 10107 25594
rect 10107 25542 10153 25594
rect 9857 25540 9913 25542
rect 9937 25540 9993 25542
rect 10017 25540 10073 25542
rect 10097 25540 10153 25542
rect 9857 24506 9913 24508
rect 9937 24506 9993 24508
rect 10017 24506 10073 24508
rect 10097 24506 10153 24508
rect 9857 24454 9903 24506
rect 9903 24454 9913 24506
rect 9937 24454 9967 24506
rect 9967 24454 9979 24506
rect 9979 24454 9993 24506
rect 10017 24454 10031 24506
rect 10031 24454 10043 24506
rect 10043 24454 10073 24506
rect 10097 24454 10107 24506
rect 10107 24454 10153 24506
rect 9857 24452 9913 24454
rect 9937 24452 9993 24454
rect 10017 24452 10073 24454
rect 10097 24452 10153 24454
rect 10138 24112 10194 24168
rect 9857 23418 9913 23420
rect 9937 23418 9993 23420
rect 10017 23418 10073 23420
rect 10097 23418 10153 23420
rect 9857 23366 9903 23418
rect 9903 23366 9913 23418
rect 9937 23366 9967 23418
rect 9967 23366 9979 23418
rect 9979 23366 9993 23418
rect 10017 23366 10031 23418
rect 10031 23366 10043 23418
rect 10043 23366 10073 23418
rect 10097 23366 10107 23418
rect 10107 23366 10153 23418
rect 9857 23364 9913 23366
rect 9937 23364 9993 23366
rect 10017 23364 10073 23366
rect 10097 23364 10153 23366
rect 10046 22752 10102 22808
rect 9857 22330 9913 22332
rect 9937 22330 9993 22332
rect 10017 22330 10073 22332
rect 10097 22330 10153 22332
rect 9857 22278 9903 22330
rect 9903 22278 9913 22330
rect 9937 22278 9967 22330
rect 9967 22278 9979 22330
rect 9979 22278 9993 22330
rect 10017 22278 10031 22330
rect 10031 22278 10043 22330
rect 10043 22278 10073 22330
rect 10097 22278 10107 22330
rect 10107 22278 10153 22330
rect 9857 22276 9913 22278
rect 9937 22276 9993 22278
rect 10017 22276 10073 22278
rect 10097 22276 10153 22278
rect 9770 21936 9826 21992
rect 9586 21664 9642 21720
rect 9402 21256 9458 21312
rect 9857 21242 9913 21244
rect 9937 21242 9993 21244
rect 10017 21242 10073 21244
rect 10097 21242 10153 21244
rect 9857 21190 9903 21242
rect 9903 21190 9913 21242
rect 9937 21190 9967 21242
rect 9967 21190 9979 21242
rect 9979 21190 9993 21242
rect 10017 21190 10031 21242
rect 10031 21190 10043 21242
rect 10043 21190 10073 21242
rect 10097 21190 10107 21242
rect 10107 21190 10153 21242
rect 9857 21188 9913 21190
rect 9937 21188 9993 21190
rect 10017 21188 10073 21190
rect 10097 21188 10153 21190
rect 9862 20984 9918 21040
rect 10138 21004 10194 21040
rect 10138 20984 10140 21004
rect 10140 20984 10192 21004
rect 10192 20984 10194 21004
rect 9954 20476 9956 20496
rect 9956 20476 10008 20496
rect 10008 20476 10010 20496
rect 9954 20440 10010 20476
rect 10322 25880 10378 25936
rect 9857 20154 9913 20156
rect 9937 20154 9993 20156
rect 10017 20154 10073 20156
rect 10097 20154 10153 20156
rect 9857 20102 9903 20154
rect 9903 20102 9913 20154
rect 9937 20102 9967 20154
rect 9967 20102 9979 20154
rect 9979 20102 9993 20154
rect 10017 20102 10031 20154
rect 10031 20102 10043 20154
rect 10043 20102 10073 20154
rect 10097 20102 10107 20154
rect 10107 20102 10153 20154
rect 9857 20100 9913 20102
rect 9937 20100 9993 20102
rect 10017 20100 10073 20102
rect 10097 20100 10153 20102
rect 9494 19352 9550 19408
rect 9126 17040 9182 17096
rect 8850 16496 8906 16552
rect 8758 8336 8814 8392
rect 9402 15544 9458 15600
rect 9862 19896 9918 19952
rect 10230 19352 10286 19408
rect 9857 19066 9913 19068
rect 9937 19066 9993 19068
rect 10017 19066 10073 19068
rect 10097 19066 10153 19068
rect 9857 19014 9903 19066
rect 9903 19014 9913 19066
rect 9937 19014 9967 19066
rect 9967 19014 9979 19066
rect 9979 19014 9993 19066
rect 10017 19014 10031 19066
rect 10031 19014 10043 19066
rect 10043 19014 10073 19066
rect 10097 19014 10107 19066
rect 10107 19014 10153 19066
rect 9857 19012 9913 19014
rect 9937 19012 9993 19014
rect 10017 19012 10073 19014
rect 10097 19012 10153 19014
rect 9586 17312 9642 17368
rect 9857 17978 9913 17980
rect 9937 17978 9993 17980
rect 10017 17978 10073 17980
rect 10097 17978 10153 17980
rect 9857 17926 9903 17978
rect 9903 17926 9913 17978
rect 9937 17926 9967 17978
rect 9967 17926 9979 17978
rect 9979 17926 9993 17978
rect 10017 17926 10031 17978
rect 10031 17926 10043 17978
rect 10043 17926 10073 17978
rect 10097 17926 10107 17978
rect 10107 17926 10153 17978
rect 9857 17924 9913 17926
rect 9937 17924 9993 17926
rect 10017 17924 10073 17926
rect 10097 17924 10153 17926
rect 12824 43546 12880 43548
rect 12904 43546 12960 43548
rect 12984 43546 13040 43548
rect 13064 43546 13120 43548
rect 12824 43494 12870 43546
rect 12870 43494 12880 43546
rect 12904 43494 12934 43546
rect 12934 43494 12946 43546
rect 12946 43494 12960 43546
rect 12984 43494 12998 43546
rect 12998 43494 13010 43546
rect 13010 43494 13040 43546
rect 13064 43494 13074 43546
rect 13074 43494 13120 43546
rect 12824 43492 12880 43494
rect 12904 43492 12960 43494
rect 12984 43492 13040 43494
rect 13064 43492 13120 43494
rect 12898 43288 12954 43344
rect 11242 36236 11298 36272
rect 11242 36216 11244 36236
rect 11244 36216 11296 36236
rect 11296 36216 11298 36236
rect 10966 30640 11022 30696
rect 11242 32680 11298 32736
rect 11150 31356 11152 31376
rect 11152 31356 11204 31376
rect 11204 31356 11206 31376
rect 11150 31320 11206 31356
rect 11058 30232 11114 30288
rect 11242 30096 11298 30152
rect 11794 41928 11850 41984
rect 11518 35808 11574 35864
rect 12530 42880 12586 42936
rect 12070 42064 12126 42120
rect 12824 42458 12880 42460
rect 12904 42458 12960 42460
rect 12984 42458 13040 42460
rect 13064 42458 13120 42460
rect 12824 42406 12870 42458
rect 12870 42406 12880 42458
rect 12904 42406 12934 42458
rect 12934 42406 12946 42458
rect 12946 42406 12960 42458
rect 12984 42406 12998 42458
rect 12998 42406 13010 42458
rect 13010 42406 13040 42458
rect 13064 42406 13074 42458
rect 13074 42406 13120 42458
rect 12824 42404 12880 42406
rect 12904 42404 12960 42406
rect 12984 42404 13040 42406
rect 13064 42404 13120 42406
rect 11978 38936 12034 38992
rect 12824 41370 12880 41372
rect 12904 41370 12960 41372
rect 12984 41370 13040 41372
rect 13064 41370 13120 41372
rect 12824 41318 12870 41370
rect 12870 41318 12880 41370
rect 12904 41318 12934 41370
rect 12934 41318 12946 41370
rect 12946 41318 12960 41370
rect 12984 41318 12998 41370
rect 12998 41318 13010 41370
rect 13010 41318 13040 41370
rect 13064 41318 13074 41370
rect 13074 41318 13120 41370
rect 12824 41316 12880 41318
rect 12904 41316 12960 41318
rect 12984 41316 13040 41318
rect 13064 41316 13120 41318
rect 12824 40282 12880 40284
rect 12904 40282 12960 40284
rect 12984 40282 13040 40284
rect 13064 40282 13120 40284
rect 12824 40230 12870 40282
rect 12870 40230 12880 40282
rect 12904 40230 12934 40282
rect 12934 40230 12946 40282
rect 12946 40230 12960 40282
rect 12984 40230 12998 40282
rect 12998 40230 13010 40282
rect 13010 40230 13040 40282
rect 13064 40230 13074 40282
rect 13074 40230 13120 40282
rect 12824 40228 12880 40230
rect 12904 40228 12960 40230
rect 12984 40228 13040 40230
rect 13064 40228 13120 40230
rect 12824 39194 12880 39196
rect 12904 39194 12960 39196
rect 12984 39194 13040 39196
rect 13064 39194 13120 39196
rect 12824 39142 12870 39194
rect 12870 39142 12880 39194
rect 12904 39142 12934 39194
rect 12934 39142 12946 39194
rect 12946 39142 12960 39194
rect 12984 39142 12998 39194
rect 12998 39142 13010 39194
rect 13010 39142 13040 39194
rect 13064 39142 13074 39194
rect 13074 39142 13120 39194
rect 12824 39140 12880 39142
rect 12904 39140 12960 39142
rect 12984 39140 13040 39142
rect 13064 39140 13120 39142
rect 12070 36896 12126 36952
rect 12254 37168 12310 37224
rect 12070 35028 12072 35048
rect 12072 35028 12124 35048
rect 12124 35028 12126 35048
rect 12070 34992 12126 35028
rect 11610 30640 11666 30696
rect 11058 29180 11060 29200
rect 11060 29180 11112 29200
rect 11112 29180 11114 29200
rect 11058 29144 11114 29180
rect 10782 27396 10838 27432
rect 10782 27376 10784 27396
rect 10784 27376 10836 27396
rect 10836 27376 10838 27396
rect 10782 26444 10838 26480
rect 10782 26424 10784 26444
rect 10784 26424 10836 26444
rect 10836 26424 10838 26444
rect 10598 24248 10654 24304
rect 11334 26424 11390 26480
rect 10874 23840 10930 23896
rect 10874 23432 10930 23488
rect 11150 22888 11206 22944
rect 10414 19216 10470 19272
rect 10598 19760 10654 19816
rect 10414 17992 10470 18048
rect 9857 16890 9913 16892
rect 9937 16890 9993 16892
rect 10017 16890 10073 16892
rect 10097 16890 10153 16892
rect 9857 16838 9903 16890
rect 9903 16838 9913 16890
rect 9937 16838 9967 16890
rect 9967 16838 9979 16890
rect 9979 16838 9993 16890
rect 10017 16838 10031 16890
rect 10031 16838 10043 16890
rect 10043 16838 10073 16890
rect 10097 16838 10107 16890
rect 10107 16838 10153 16890
rect 9857 16836 9913 16838
rect 9937 16836 9993 16838
rect 10017 16836 10073 16838
rect 10097 16836 10153 16838
rect 9857 15802 9913 15804
rect 9937 15802 9993 15804
rect 10017 15802 10073 15804
rect 10097 15802 10153 15804
rect 9857 15750 9903 15802
rect 9903 15750 9913 15802
rect 9937 15750 9967 15802
rect 9967 15750 9979 15802
rect 9979 15750 9993 15802
rect 10017 15750 10031 15802
rect 10031 15750 10043 15802
rect 10043 15750 10073 15802
rect 10097 15750 10107 15802
rect 10107 15750 10153 15802
rect 9857 15748 9913 15750
rect 9937 15748 9993 15750
rect 10017 15748 10073 15750
rect 10097 15748 10153 15750
rect 9954 15136 10010 15192
rect 9857 14714 9913 14716
rect 9937 14714 9993 14716
rect 10017 14714 10073 14716
rect 10097 14714 10153 14716
rect 9857 14662 9903 14714
rect 9903 14662 9913 14714
rect 9937 14662 9967 14714
rect 9967 14662 9979 14714
rect 9979 14662 9993 14714
rect 10017 14662 10031 14714
rect 10031 14662 10043 14714
rect 10043 14662 10073 14714
rect 10097 14662 10107 14714
rect 10107 14662 10153 14714
rect 9857 14660 9913 14662
rect 9937 14660 9993 14662
rect 10017 14660 10073 14662
rect 10097 14660 10153 14662
rect 10046 14184 10102 14240
rect 8942 8880 8998 8936
rect 9034 7792 9090 7848
rect 9310 9580 9366 9616
rect 9310 9560 9312 9580
rect 9312 9560 9364 9580
rect 9364 9560 9366 9580
rect 9402 8880 9458 8936
rect 9857 13626 9913 13628
rect 9937 13626 9993 13628
rect 10017 13626 10073 13628
rect 10097 13626 10153 13628
rect 9857 13574 9903 13626
rect 9903 13574 9913 13626
rect 9937 13574 9967 13626
rect 9967 13574 9979 13626
rect 9979 13574 9993 13626
rect 10017 13574 10031 13626
rect 10031 13574 10043 13626
rect 10043 13574 10073 13626
rect 10097 13574 10107 13626
rect 10107 13574 10153 13626
rect 9857 13572 9913 13574
rect 9937 13572 9993 13574
rect 10017 13572 10073 13574
rect 10097 13572 10153 13574
rect 10874 21528 10930 21584
rect 11058 21936 11114 21992
rect 11334 24132 11390 24168
rect 11334 24112 11336 24132
rect 11336 24112 11388 24132
rect 11388 24112 11390 24132
rect 11518 23160 11574 23216
rect 11334 22480 11390 22536
rect 11242 20324 11298 20360
rect 11242 20304 11244 20324
rect 11244 20304 11296 20324
rect 11296 20304 11298 20324
rect 11426 19352 11482 19408
rect 10690 14864 10746 14920
rect 10414 14184 10470 14240
rect 10138 13096 10194 13152
rect 9857 12538 9913 12540
rect 9937 12538 9993 12540
rect 10017 12538 10073 12540
rect 10097 12538 10153 12540
rect 9857 12486 9903 12538
rect 9903 12486 9913 12538
rect 9937 12486 9967 12538
rect 9967 12486 9979 12538
rect 9979 12486 9993 12538
rect 10017 12486 10031 12538
rect 10031 12486 10043 12538
rect 10043 12486 10073 12538
rect 10097 12486 10107 12538
rect 10107 12486 10153 12538
rect 9857 12484 9913 12486
rect 9937 12484 9993 12486
rect 10017 12484 10073 12486
rect 10097 12484 10153 12486
rect 9857 11450 9913 11452
rect 9937 11450 9993 11452
rect 10017 11450 10073 11452
rect 10097 11450 10153 11452
rect 9857 11398 9903 11450
rect 9903 11398 9913 11450
rect 9937 11398 9967 11450
rect 9967 11398 9979 11450
rect 9979 11398 9993 11450
rect 10017 11398 10031 11450
rect 10031 11398 10043 11450
rect 10043 11398 10073 11450
rect 10097 11398 10107 11450
rect 10107 11398 10153 11450
rect 9857 11396 9913 11398
rect 9937 11396 9993 11398
rect 10017 11396 10073 11398
rect 10097 11396 10153 11398
rect 9857 10362 9913 10364
rect 9937 10362 9993 10364
rect 10017 10362 10073 10364
rect 10097 10362 10153 10364
rect 9857 10310 9903 10362
rect 9903 10310 9913 10362
rect 9937 10310 9967 10362
rect 9967 10310 9979 10362
rect 9979 10310 9993 10362
rect 10017 10310 10031 10362
rect 10031 10310 10043 10362
rect 10043 10310 10073 10362
rect 10097 10310 10107 10362
rect 10107 10310 10153 10362
rect 9857 10308 9913 10310
rect 9937 10308 9993 10310
rect 10017 10308 10073 10310
rect 10097 10308 10153 10310
rect 9770 10104 9826 10160
rect 9678 9560 9734 9616
rect 9586 9460 9588 9480
rect 9588 9460 9640 9480
rect 9640 9460 9642 9480
rect 9586 9424 9642 9460
rect 9857 9274 9913 9276
rect 9937 9274 9993 9276
rect 10017 9274 10073 9276
rect 10097 9274 10153 9276
rect 9857 9222 9903 9274
rect 9903 9222 9913 9274
rect 9937 9222 9967 9274
rect 9967 9222 9979 9274
rect 9979 9222 9993 9274
rect 10017 9222 10031 9274
rect 10031 9222 10043 9274
rect 10043 9222 10073 9274
rect 10097 9222 10107 9274
rect 10107 9222 10153 9274
rect 9857 9220 9913 9222
rect 9937 9220 9993 9222
rect 10017 9220 10073 9222
rect 10097 9220 10153 9222
rect 9857 8186 9913 8188
rect 9937 8186 9993 8188
rect 10017 8186 10073 8188
rect 10097 8186 10153 8188
rect 9857 8134 9903 8186
rect 9903 8134 9913 8186
rect 9937 8134 9967 8186
rect 9967 8134 9979 8186
rect 9979 8134 9993 8186
rect 10017 8134 10031 8186
rect 10031 8134 10043 8186
rect 10043 8134 10073 8186
rect 10097 8134 10107 8186
rect 10107 8134 10153 8186
rect 9857 8132 9913 8134
rect 9937 8132 9993 8134
rect 10017 8132 10073 8134
rect 10097 8132 10153 8134
rect 9770 7948 9826 7984
rect 9770 7928 9772 7948
rect 9772 7928 9824 7948
rect 9824 7928 9826 7948
rect 8574 6840 8630 6896
rect 9310 6024 9366 6080
rect 10414 13232 10470 13288
rect 10506 12280 10562 12336
rect 10690 13268 10692 13288
rect 10692 13268 10744 13288
rect 10744 13268 10746 13288
rect 10690 13232 10746 13268
rect 11058 17196 11114 17232
rect 11058 17176 11060 17196
rect 11060 17176 11112 17196
rect 11112 17176 11114 17196
rect 11426 19216 11482 19272
rect 11150 13912 11206 13968
rect 10782 10240 10838 10296
rect 9857 7098 9913 7100
rect 9937 7098 9993 7100
rect 10017 7098 10073 7100
rect 10097 7098 10153 7100
rect 9857 7046 9903 7098
rect 9903 7046 9913 7098
rect 9937 7046 9967 7098
rect 9967 7046 9979 7098
rect 9979 7046 9993 7098
rect 10017 7046 10031 7098
rect 10031 7046 10043 7098
rect 10043 7046 10073 7098
rect 10097 7046 10107 7098
rect 10107 7046 10153 7098
rect 9857 7044 9913 7046
rect 9937 7044 9993 7046
rect 10017 7044 10073 7046
rect 10097 7044 10153 7046
rect 9678 5616 9734 5672
rect 9310 5480 9366 5536
rect 9218 4664 9274 4720
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 9034 3596 9090 3632
rect 9034 3576 9036 3596
rect 9036 3576 9088 3596
rect 9088 3576 9090 3596
rect 9034 1300 9036 1320
rect 9036 1300 9088 1320
rect 9088 1300 9090 1320
rect 9034 1264 9090 1300
rect 9678 3712 9734 3768
rect 9678 3304 9734 3360
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 10966 10104 11022 10160
rect 11886 30504 11942 30560
rect 11794 30232 11850 30288
rect 11794 29028 11850 29064
rect 11794 29008 11796 29028
rect 11796 29008 11848 29028
rect 11848 29008 11850 29028
rect 11702 26152 11758 26208
rect 12070 28192 12126 28248
rect 11886 26016 11942 26072
rect 11794 25336 11850 25392
rect 11978 25064 12034 25120
rect 11886 24248 11942 24304
rect 12824 38106 12880 38108
rect 12904 38106 12960 38108
rect 12984 38106 13040 38108
rect 13064 38106 13120 38108
rect 12824 38054 12870 38106
rect 12870 38054 12880 38106
rect 12904 38054 12934 38106
rect 12934 38054 12946 38106
rect 12946 38054 12960 38106
rect 12984 38054 12998 38106
rect 12998 38054 13010 38106
rect 13010 38054 13040 38106
rect 13064 38054 13074 38106
rect 13074 38054 13120 38106
rect 12824 38052 12880 38054
rect 12904 38052 12960 38054
rect 12984 38052 13040 38054
rect 13064 38052 13120 38054
rect 12824 37018 12880 37020
rect 12904 37018 12960 37020
rect 12984 37018 13040 37020
rect 13064 37018 13120 37020
rect 12824 36966 12870 37018
rect 12870 36966 12880 37018
rect 12904 36966 12934 37018
rect 12934 36966 12946 37018
rect 12946 36966 12960 37018
rect 12984 36966 12998 37018
rect 12998 36966 13010 37018
rect 13010 36966 13040 37018
rect 13064 36966 13074 37018
rect 13074 36966 13120 37018
rect 12824 36964 12880 36966
rect 12904 36964 12960 36966
rect 12984 36964 13040 36966
rect 13064 36964 13120 36966
rect 12438 35808 12494 35864
rect 12824 35930 12880 35932
rect 12904 35930 12960 35932
rect 12984 35930 13040 35932
rect 13064 35930 13120 35932
rect 12824 35878 12870 35930
rect 12870 35878 12880 35930
rect 12904 35878 12934 35930
rect 12934 35878 12946 35930
rect 12946 35878 12960 35930
rect 12984 35878 12998 35930
rect 12998 35878 13010 35930
rect 13010 35878 13040 35930
rect 13064 35878 13074 35930
rect 13074 35878 13120 35930
rect 12824 35876 12880 35878
rect 12904 35876 12960 35878
rect 12984 35876 13040 35878
rect 13064 35876 13120 35878
rect 12990 35556 13046 35592
rect 12990 35536 12992 35556
rect 12992 35536 13044 35556
rect 13044 35536 13046 35556
rect 13450 35400 13506 35456
rect 13358 35128 13414 35184
rect 12824 34842 12880 34844
rect 12904 34842 12960 34844
rect 12984 34842 13040 34844
rect 13064 34842 13120 34844
rect 12824 34790 12870 34842
rect 12870 34790 12880 34842
rect 12904 34790 12934 34842
rect 12934 34790 12946 34842
rect 12946 34790 12960 34842
rect 12984 34790 12998 34842
rect 12998 34790 13010 34842
rect 13010 34790 13040 34842
rect 13064 34790 13074 34842
rect 13074 34790 13120 34842
rect 12824 34788 12880 34790
rect 12904 34788 12960 34790
rect 12984 34788 13040 34790
rect 13064 34788 13120 34790
rect 13266 34720 13322 34776
rect 13082 34448 13138 34504
rect 12530 34060 12586 34096
rect 12530 34040 12532 34060
rect 12532 34040 12584 34060
rect 12584 34040 12586 34060
rect 12346 33924 12402 33960
rect 12346 33904 12348 33924
rect 12348 33904 12400 33924
rect 12400 33904 12402 33924
rect 12530 33904 12586 33960
rect 12824 33754 12880 33756
rect 12904 33754 12960 33756
rect 12984 33754 13040 33756
rect 13064 33754 13120 33756
rect 12824 33702 12870 33754
rect 12870 33702 12880 33754
rect 12904 33702 12934 33754
rect 12934 33702 12946 33754
rect 12946 33702 12960 33754
rect 12984 33702 12998 33754
rect 12998 33702 13010 33754
rect 13010 33702 13040 33754
rect 13064 33702 13074 33754
rect 13074 33702 13120 33754
rect 12824 33700 12880 33702
rect 12904 33700 12960 33702
rect 12984 33700 13040 33702
rect 13064 33700 13120 33702
rect 12622 31456 12678 31512
rect 12824 32666 12880 32668
rect 12904 32666 12960 32668
rect 12984 32666 13040 32668
rect 13064 32666 13120 32668
rect 12824 32614 12870 32666
rect 12870 32614 12880 32666
rect 12904 32614 12934 32666
rect 12934 32614 12946 32666
rect 12946 32614 12960 32666
rect 12984 32614 12998 32666
rect 12998 32614 13010 32666
rect 13010 32614 13040 32666
rect 13064 32614 13074 32666
rect 13074 32614 13120 32666
rect 12824 32612 12880 32614
rect 12904 32612 12960 32614
rect 12984 32612 13040 32614
rect 13064 32612 13120 32614
rect 12824 31578 12880 31580
rect 12904 31578 12960 31580
rect 12984 31578 13040 31580
rect 13064 31578 13120 31580
rect 12824 31526 12870 31578
rect 12870 31526 12880 31578
rect 12904 31526 12934 31578
rect 12934 31526 12946 31578
rect 12946 31526 12960 31578
rect 12984 31526 12998 31578
rect 12998 31526 13010 31578
rect 13010 31526 13040 31578
rect 13064 31526 13074 31578
rect 13074 31526 13120 31578
rect 12824 31524 12880 31526
rect 12904 31524 12960 31526
rect 12984 31524 13040 31526
rect 13064 31524 13120 31526
rect 12622 31184 12678 31240
rect 13266 31048 13322 31104
rect 12824 30490 12880 30492
rect 12904 30490 12960 30492
rect 12984 30490 13040 30492
rect 13064 30490 13120 30492
rect 12824 30438 12870 30490
rect 12870 30438 12880 30490
rect 12904 30438 12934 30490
rect 12934 30438 12946 30490
rect 12946 30438 12960 30490
rect 12984 30438 12998 30490
rect 12998 30438 13010 30490
rect 13010 30438 13040 30490
rect 13064 30438 13074 30490
rect 13074 30438 13120 30490
rect 12824 30436 12880 30438
rect 12904 30436 12960 30438
rect 12984 30436 13040 30438
rect 13064 30436 13120 30438
rect 12622 30368 12678 30424
rect 12824 29402 12880 29404
rect 12904 29402 12960 29404
rect 12984 29402 13040 29404
rect 13064 29402 13120 29404
rect 12824 29350 12870 29402
rect 12870 29350 12880 29402
rect 12904 29350 12934 29402
rect 12934 29350 12946 29402
rect 12946 29350 12960 29402
rect 12984 29350 12998 29402
rect 12998 29350 13010 29402
rect 13010 29350 13040 29402
rect 13064 29350 13074 29402
rect 13074 29350 13120 29402
rect 12824 29348 12880 29350
rect 12904 29348 12960 29350
rect 12984 29348 13040 29350
rect 13064 29348 13120 29350
rect 12530 28872 12586 28928
rect 12438 28056 12494 28112
rect 12824 28314 12880 28316
rect 12904 28314 12960 28316
rect 12984 28314 13040 28316
rect 13064 28314 13120 28316
rect 12824 28262 12870 28314
rect 12870 28262 12880 28314
rect 12904 28262 12934 28314
rect 12934 28262 12946 28314
rect 12946 28262 12960 28314
rect 12984 28262 12998 28314
rect 12998 28262 13010 28314
rect 13010 28262 13040 28314
rect 13064 28262 13074 28314
rect 13074 28262 13120 28314
rect 12824 28260 12880 28262
rect 12904 28260 12960 28262
rect 12984 28260 13040 28262
rect 13064 28260 13120 28262
rect 13174 27376 13230 27432
rect 12824 27226 12880 27228
rect 12904 27226 12960 27228
rect 12984 27226 13040 27228
rect 13064 27226 13120 27228
rect 12824 27174 12870 27226
rect 12870 27174 12880 27226
rect 12904 27174 12934 27226
rect 12934 27174 12946 27226
rect 12946 27174 12960 27226
rect 12984 27174 12998 27226
rect 12998 27174 13010 27226
rect 13010 27174 13040 27226
rect 13064 27174 13074 27226
rect 13074 27174 13120 27226
rect 12824 27172 12880 27174
rect 12904 27172 12960 27174
rect 12984 27172 13040 27174
rect 13064 27172 13120 27174
rect 12824 26138 12880 26140
rect 12904 26138 12960 26140
rect 12984 26138 13040 26140
rect 13064 26138 13120 26140
rect 12824 26086 12870 26138
rect 12870 26086 12880 26138
rect 12904 26086 12934 26138
rect 12934 26086 12946 26138
rect 12946 26086 12960 26138
rect 12984 26086 12998 26138
rect 12998 26086 13010 26138
rect 13010 26086 13040 26138
rect 13064 26086 13074 26138
rect 13074 26086 13120 26138
rect 12824 26084 12880 26086
rect 12904 26084 12960 26086
rect 12984 26084 13040 26086
rect 13064 26084 13120 26086
rect 12824 25050 12880 25052
rect 12904 25050 12960 25052
rect 12984 25050 13040 25052
rect 13064 25050 13120 25052
rect 12824 24998 12870 25050
rect 12870 24998 12880 25050
rect 12904 24998 12934 25050
rect 12934 24998 12946 25050
rect 12946 24998 12960 25050
rect 12984 24998 12998 25050
rect 12998 24998 13010 25050
rect 13010 24998 13040 25050
rect 13064 24998 13074 25050
rect 13074 24998 13120 25050
rect 12824 24996 12880 24998
rect 12904 24996 12960 24998
rect 12984 24996 13040 24998
rect 13064 24996 13120 24998
rect 12070 23568 12126 23624
rect 11794 22752 11850 22808
rect 11702 21392 11758 21448
rect 11794 21004 11850 21040
rect 11794 20984 11796 21004
rect 11796 20984 11848 21004
rect 11848 20984 11850 21004
rect 11518 17720 11574 17776
rect 11242 12280 11298 12336
rect 10506 5752 10562 5808
rect 9954 3440 10010 3496
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 10322 2216 10378 2272
rect 11058 9424 11114 9480
rect 10966 8472 11022 8528
rect 11242 6976 11298 7032
rect 10966 5888 11022 5944
rect 11058 3732 11114 3768
rect 11058 3712 11060 3732
rect 11060 3712 11112 3732
rect 11112 3712 11114 3732
rect 10690 3304 10746 3360
rect 11058 3068 11060 3088
rect 11060 3068 11112 3088
rect 11112 3068 11114 3088
rect 11058 3032 11114 3068
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 12622 24112 12678 24168
rect 12622 23024 12678 23080
rect 12824 23962 12880 23964
rect 12904 23962 12960 23964
rect 12984 23962 13040 23964
rect 13064 23962 13120 23964
rect 12824 23910 12870 23962
rect 12870 23910 12880 23962
rect 12904 23910 12934 23962
rect 12934 23910 12946 23962
rect 12946 23910 12960 23962
rect 12984 23910 12998 23962
rect 12998 23910 13010 23962
rect 13010 23910 13040 23962
rect 13064 23910 13074 23962
rect 13074 23910 13120 23962
rect 12824 23908 12880 23910
rect 12904 23908 12960 23910
rect 12984 23908 13040 23910
rect 13064 23908 13120 23910
rect 13266 23568 13322 23624
rect 12824 22874 12880 22876
rect 12904 22874 12960 22876
rect 12984 22874 13040 22876
rect 13064 22874 13120 22876
rect 12824 22822 12870 22874
rect 12870 22822 12880 22874
rect 12904 22822 12934 22874
rect 12934 22822 12946 22874
rect 12946 22822 12960 22874
rect 12984 22822 12998 22874
rect 12998 22822 13010 22874
rect 13010 22822 13040 22874
rect 13064 22822 13074 22874
rect 13074 22822 13120 22874
rect 12824 22820 12880 22822
rect 12904 22820 12960 22822
rect 12984 22820 13040 22822
rect 13064 22820 13120 22822
rect 12824 21786 12880 21788
rect 12904 21786 12960 21788
rect 12984 21786 13040 21788
rect 13064 21786 13120 21788
rect 12824 21734 12870 21786
rect 12870 21734 12880 21786
rect 12904 21734 12934 21786
rect 12934 21734 12946 21786
rect 12946 21734 12960 21786
rect 12984 21734 12998 21786
rect 12998 21734 13010 21786
rect 13010 21734 13040 21786
rect 13064 21734 13074 21786
rect 13074 21734 13120 21786
rect 12824 21732 12880 21734
rect 12904 21732 12960 21734
rect 12984 21732 13040 21734
rect 13064 21732 13120 21734
rect 12622 20712 12678 20768
rect 13174 20848 13230 20904
rect 12824 20698 12880 20700
rect 12904 20698 12960 20700
rect 12984 20698 13040 20700
rect 13064 20698 13120 20700
rect 12824 20646 12870 20698
rect 12870 20646 12880 20698
rect 12904 20646 12934 20698
rect 12934 20646 12946 20698
rect 12946 20646 12960 20698
rect 12984 20646 12998 20698
rect 12998 20646 13010 20698
rect 13010 20646 13040 20698
rect 13064 20646 13074 20698
rect 13074 20646 13120 20698
rect 12824 20644 12880 20646
rect 12904 20644 12960 20646
rect 12984 20644 13040 20646
rect 13064 20644 13120 20646
rect 12346 19352 12402 19408
rect 11610 13096 11666 13152
rect 12070 15136 12126 15192
rect 11426 4528 11482 4584
rect 12254 17584 12310 17640
rect 12530 19896 12586 19952
rect 12824 19610 12880 19612
rect 12904 19610 12960 19612
rect 12984 19610 13040 19612
rect 13064 19610 13120 19612
rect 12824 19558 12870 19610
rect 12870 19558 12880 19610
rect 12904 19558 12934 19610
rect 12934 19558 12946 19610
rect 12946 19558 12960 19610
rect 12984 19558 12998 19610
rect 12998 19558 13010 19610
rect 13010 19558 13040 19610
rect 13064 19558 13074 19610
rect 13074 19558 13120 19610
rect 12824 19556 12880 19558
rect 12904 19556 12960 19558
rect 12984 19556 13040 19558
rect 13064 19556 13120 19558
rect 12622 18400 12678 18456
rect 12824 18522 12880 18524
rect 12904 18522 12960 18524
rect 12984 18522 13040 18524
rect 13064 18522 13120 18524
rect 12824 18470 12870 18522
rect 12870 18470 12880 18522
rect 12904 18470 12934 18522
rect 12934 18470 12946 18522
rect 12946 18470 12960 18522
rect 12984 18470 12998 18522
rect 12998 18470 13010 18522
rect 13010 18470 13040 18522
rect 13064 18470 13074 18522
rect 13074 18470 13120 18522
rect 12824 18468 12880 18470
rect 12904 18468 12960 18470
rect 12984 18468 13040 18470
rect 13064 18468 13120 18470
rect 12530 17992 12586 18048
rect 12530 16632 12586 16688
rect 12346 15408 12402 15464
rect 13542 32836 13598 32872
rect 13542 32816 13544 32836
rect 13544 32816 13596 32836
rect 13596 32816 13598 32836
rect 14278 42880 14334 42936
rect 14922 42880 14978 42936
rect 15290 43052 15292 43072
rect 15292 43052 15344 43072
rect 15344 43052 15346 43072
rect 15290 43016 15346 43052
rect 15474 42608 15530 42664
rect 13910 33940 13912 33960
rect 13912 33940 13964 33960
rect 13964 33940 13966 33960
rect 13910 33904 13966 33940
rect 13910 31592 13966 31648
rect 13818 29008 13874 29064
rect 13634 26968 13690 27024
rect 14462 37712 14518 37768
rect 14278 36080 14334 36136
rect 14094 27784 14150 27840
rect 14094 25880 14150 25936
rect 13726 24656 13782 24712
rect 13818 23568 13874 23624
rect 13266 20440 13322 20496
rect 13542 19760 13598 19816
rect 13174 17992 13230 18048
rect 12824 17434 12880 17436
rect 12904 17434 12960 17436
rect 12984 17434 13040 17436
rect 13064 17434 13120 17436
rect 12824 17382 12870 17434
rect 12870 17382 12880 17434
rect 12904 17382 12934 17434
rect 12934 17382 12946 17434
rect 12946 17382 12960 17434
rect 12984 17382 12998 17434
rect 12998 17382 13010 17434
rect 13010 17382 13040 17434
rect 13064 17382 13074 17434
rect 13074 17382 13120 17434
rect 12824 17380 12880 17382
rect 12904 17380 12960 17382
rect 12984 17380 13040 17382
rect 13064 17380 13120 17382
rect 12824 16346 12880 16348
rect 12904 16346 12960 16348
rect 12984 16346 13040 16348
rect 13064 16346 13120 16348
rect 12824 16294 12870 16346
rect 12870 16294 12880 16346
rect 12904 16294 12934 16346
rect 12934 16294 12946 16346
rect 12946 16294 12960 16346
rect 12984 16294 12998 16346
rect 12998 16294 13010 16346
rect 13010 16294 13040 16346
rect 13064 16294 13074 16346
rect 13074 16294 13120 16346
rect 12824 16292 12880 16294
rect 12904 16292 12960 16294
rect 12984 16292 13040 16294
rect 13064 16292 13120 16294
rect 12824 15258 12880 15260
rect 12904 15258 12960 15260
rect 12984 15258 13040 15260
rect 13064 15258 13120 15260
rect 12824 15206 12870 15258
rect 12870 15206 12880 15258
rect 12904 15206 12934 15258
rect 12934 15206 12946 15258
rect 12946 15206 12960 15258
rect 12984 15206 12998 15258
rect 12998 15206 13010 15258
rect 13010 15206 13040 15258
rect 13064 15206 13074 15258
rect 13074 15206 13120 15258
rect 12824 15204 12880 15206
rect 12904 15204 12960 15206
rect 12984 15204 13040 15206
rect 13064 15204 13120 15206
rect 12824 14170 12880 14172
rect 12904 14170 12960 14172
rect 12984 14170 13040 14172
rect 13064 14170 13120 14172
rect 12824 14118 12870 14170
rect 12870 14118 12880 14170
rect 12904 14118 12934 14170
rect 12934 14118 12946 14170
rect 12946 14118 12960 14170
rect 12984 14118 12998 14170
rect 12998 14118 13010 14170
rect 13010 14118 13040 14170
rect 13064 14118 13074 14170
rect 13074 14118 13120 14170
rect 12824 14116 12880 14118
rect 12904 14116 12960 14118
rect 12984 14116 13040 14118
rect 13064 14116 13120 14118
rect 13174 13812 13176 13832
rect 13176 13812 13228 13832
rect 13228 13812 13230 13832
rect 13174 13776 13230 13812
rect 12824 13082 12880 13084
rect 12904 13082 12960 13084
rect 12984 13082 13040 13084
rect 13064 13082 13120 13084
rect 12824 13030 12870 13082
rect 12870 13030 12880 13082
rect 12904 13030 12934 13082
rect 12934 13030 12946 13082
rect 12946 13030 12960 13082
rect 12984 13030 12998 13082
rect 12998 13030 13010 13082
rect 13010 13030 13040 13082
rect 13064 13030 13074 13082
rect 13074 13030 13120 13082
rect 12824 13028 12880 13030
rect 12904 13028 12960 13030
rect 12984 13028 13040 13030
rect 13064 13028 13120 13030
rect 12824 11994 12880 11996
rect 12904 11994 12960 11996
rect 12984 11994 13040 11996
rect 13064 11994 13120 11996
rect 12824 11942 12870 11994
rect 12870 11942 12880 11994
rect 12904 11942 12934 11994
rect 12934 11942 12946 11994
rect 12946 11942 12960 11994
rect 12984 11942 12998 11994
rect 12998 11942 13010 11994
rect 13010 11942 13040 11994
rect 13064 11942 13074 11994
rect 13074 11942 13120 11994
rect 12824 11940 12880 11942
rect 12904 11940 12960 11942
rect 12984 11940 13040 11942
rect 13064 11940 13120 11942
rect 12346 9696 12402 9752
rect 11978 8336 12034 8392
rect 11518 3984 11574 4040
rect 11426 3168 11482 3224
rect 11794 3984 11850 4040
rect 11886 2896 11942 2952
rect 12070 2624 12126 2680
rect 11518 1400 11574 1456
rect 12824 10906 12880 10908
rect 12904 10906 12960 10908
rect 12984 10906 13040 10908
rect 13064 10906 13120 10908
rect 12824 10854 12870 10906
rect 12870 10854 12880 10906
rect 12904 10854 12934 10906
rect 12934 10854 12946 10906
rect 12946 10854 12960 10906
rect 12984 10854 12998 10906
rect 12998 10854 13010 10906
rect 13010 10854 13040 10906
rect 13064 10854 13074 10906
rect 13074 10854 13120 10906
rect 12824 10852 12880 10854
rect 12904 10852 12960 10854
rect 12984 10852 13040 10854
rect 13064 10852 13120 10854
rect 12824 9818 12880 9820
rect 12904 9818 12960 9820
rect 12984 9818 13040 9820
rect 13064 9818 13120 9820
rect 12824 9766 12870 9818
rect 12870 9766 12880 9818
rect 12904 9766 12934 9818
rect 12934 9766 12946 9818
rect 12946 9766 12960 9818
rect 12984 9766 12998 9818
rect 12998 9766 13010 9818
rect 13010 9766 13040 9818
rect 13064 9766 13074 9818
rect 13074 9766 13120 9818
rect 12824 9764 12880 9766
rect 12904 9764 12960 9766
rect 12984 9764 13040 9766
rect 13064 9764 13120 9766
rect 12824 8730 12880 8732
rect 12904 8730 12960 8732
rect 12984 8730 13040 8732
rect 13064 8730 13120 8732
rect 12824 8678 12870 8730
rect 12870 8678 12880 8730
rect 12904 8678 12934 8730
rect 12934 8678 12946 8730
rect 12946 8678 12960 8730
rect 12984 8678 12998 8730
rect 12998 8678 13010 8730
rect 13010 8678 13040 8730
rect 13064 8678 13074 8730
rect 13074 8678 13120 8730
rect 12824 8676 12880 8678
rect 12904 8676 12960 8678
rect 12984 8676 13040 8678
rect 13064 8676 13120 8678
rect 12824 7642 12880 7644
rect 12904 7642 12960 7644
rect 12984 7642 13040 7644
rect 13064 7642 13120 7644
rect 12824 7590 12870 7642
rect 12870 7590 12880 7642
rect 12904 7590 12934 7642
rect 12934 7590 12946 7642
rect 12946 7590 12960 7642
rect 12984 7590 12998 7642
rect 12998 7590 13010 7642
rect 13010 7590 13040 7642
rect 13064 7590 13074 7642
rect 13074 7590 13120 7642
rect 12824 7588 12880 7590
rect 12904 7588 12960 7590
rect 12984 7588 13040 7590
rect 13064 7588 13120 7590
rect 13266 9968 13322 10024
rect 13450 13776 13506 13832
rect 13542 13504 13598 13560
rect 13726 11872 13782 11928
rect 13910 19388 13912 19408
rect 13912 19388 13964 19408
rect 13964 19388 13966 19408
rect 13910 19352 13966 19388
rect 14554 34584 14610 34640
rect 14462 27784 14518 27840
rect 14278 22616 14334 22672
rect 14094 17176 14150 17232
rect 14094 16632 14150 16688
rect 14462 23432 14518 23488
rect 15106 40568 15162 40624
rect 15014 34448 15070 34504
rect 15382 32816 15438 32872
rect 15290 31592 15346 31648
rect 14922 30232 14978 30288
rect 14554 22344 14610 22400
rect 15106 28600 15162 28656
rect 14922 27648 14978 27704
rect 15106 26832 15162 26888
rect 15106 24520 15162 24576
rect 15382 31184 15438 31240
rect 15474 29164 15530 29200
rect 15474 29144 15476 29164
rect 15476 29144 15528 29164
rect 15528 29144 15530 29164
rect 15290 24928 15346 24984
rect 15198 24112 15254 24168
rect 15382 24656 15438 24712
rect 15791 43002 15847 43004
rect 15871 43002 15927 43004
rect 15951 43002 16007 43004
rect 16031 43002 16087 43004
rect 15791 42950 15837 43002
rect 15837 42950 15847 43002
rect 15871 42950 15901 43002
rect 15901 42950 15913 43002
rect 15913 42950 15927 43002
rect 15951 42950 15965 43002
rect 15965 42950 15977 43002
rect 15977 42950 16007 43002
rect 16031 42950 16041 43002
rect 16041 42950 16087 43002
rect 15791 42948 15847 42950
rect 15871 42948 15927 42950
rect 15951 42948 16007 42950
rect 16031 42948 16087 42950
rect 15791 41914 15847 41916
rect 15871 41914 15927 41916
rect 15951 41914 16007 41916
rect 16031 41914 16087 41916
rect 15791 41862 15837 41914
rect 15837 41862 15847 41914
rect 15871 41862 15901 41914
rect 15901 41862 15913 41914
rect 15913 41862 15927 41914
rect 15951 41862 15965 41914
rect 15965 41862 15977 41914
rect 15977 41862 16007 41914
rect 16031 41862 16041 41914
rect 16041 41862 16087 41914
rect 15791 41860 15847 41862
rect 15871 41860 15927 41862
rect 15951 41860 16007 41862
rect 16031 41860 16087 41862
rect 15791 40826 15847 40828
rect 15871 40826 15927 40828
rect 15951 40826 16007 40828
rect 16031 40826 16087 40828
rect 15791 40774 15837 40826
rect 15837 40774 15847 40826
rect 15871 40774 15901 40826
rect 15901 40774 15913 40826
rect 15913 40774 15927 40826
rect 15951 40774 15965 40826
rect 15965 40774 15977 40826
rect 15977 40774 16007 40826
rect 16031 40774 16041 40826
rect 16041 40774 16087 40826
rect 15791 40772 15847 40774
rect 15871 40772 15927 40774
rect 15951 40772 16007 40774
rect 16031 40772 16087 40774
rect 15791 39738 15847 39740
rect 15871 39738 15927 39740
rect 15951 39738 16007 39740
rect 16031 39738 16087 39740
rect 15791 39686 15837 39738
rect 15837 39686 15847 39738
rect 15871 39686 15901 39738
rect 15901 39686 15913 39738
rect 15913 39686 15927 39738
rect 15951 39686 15965 39738
rect 15965 39686 15977 39738
rect 15977 39686 16007 39738
rect 16031 39686 16041 39738
rect 16041 39686 16087 39738
rect 15791 39684 15847 39686
rect 15871 39684 15927 39686
rect 15951 39684 16007 39686
rect 16031 39684 16087 39686
rect 15791 38650 15847 38652
rect 15871 38650 15927 38652
rect 15951 38650 16007 38652
rect 16031 38650 16087 38652
rect 15791 38598 15837 38650
rect 15837 38598 15847 38650
rect 15871 38598 15901 38650
rect 15901 38598 15913 38650
rect 15913 38598 15927 38650
rect 15951 38598 15965 38650
rect 15965 38598 15977 38650
rect 15977 38598 16007 38650
rect 16031 38598 16041 38650
rect 16041 38598 16087 38650
rect 15791 38596 15847 38598
rect 15871 38596 15927 38598
rect 15951 38596 16007 38598
rect 16031 38596 16087 38598
rect 15791 37562 15847 37564
rect 15871 37562 15927 37564
rect 15951 37562 16007 37564
rect 16031 37562 16087 37564
rect 15791 37510 15837 37562
rect 15837 37510 15847 37562
rect 15871 37510 15901 37562
rect 15901 37510 15913 37562
rect 15913 37510 15927 37562
rect 15951 37510 15965 37562
rect 15965 37510 15977 37562
rect 15977 37510 16007 37562
rect 16031 37510 16041 37562
rect 16041 37510 16087 37562
rect 15791 37508 15847 37510
rect 15871 37508 15927 37510
rect 15951 37508 16007 37510
rect 16031 37508 16087 37510
rect 15791 36474 15847 36476
rect 15871 36474 15927 36476
rect 15951 36474 16007 36476
rect 16031 36474 16087 36476
rect 15791 36422 15837 36474
rect 15837 36422 15847 36474
rect 15871 36422 15901 36474
rect 15901 36422 15913 36474
rect 15913 36422 15927 36474
rect 15951 36422 15965 36474
rect 15965 36422 15977 36474
rect 15977 36422 16007 36474
rect 16031 36422 16041 36474
rect 16041 36422 16087 36474
rect 15791 36420 15847 36422
rect 15871 36420 15927 36422
rect 15951 36420 16007 36422
rect 16031 36420 16087 36422
rect 15791 35386 15847 35388
rect 15871 35386 15927 35388
rect 15951 35386 16007 35388
rect 16031 35386 16087 35388
rect 15791 35334 15837 35386
rect 15837 35334 15847 35386
rect 15871 35334 15901 35386
rect 15901 35334 15913 35386
rect 15913 35334 15927 35386
rect 15951 35334 15965 35386
rect 15965 35334 15977 35386
rect 15977 35334 16007 35386
rect 16031 35334 16041 35386
rect 16041 35334 16087 35386
rect 15791 35332 15847 35334
rect 15871 35332 15927 35334
rect 15951 35332 16007 35334
rect 16031 35332 16087 35334
rect 15791 34298 15847 34300
rect 15871 34298 15927 34300
rect 15951 34298 16007 34300
rect 16031 34298 16087 34300
rect 15791 34246 15837 34298
rect 15837 34246 15847 34298
rect 15871 34246 15901 34298
rect 15901 34246 15913 34298
rect 15913 34246 15927 34298
rect 15951 34246 15965 34298
rect 15965 34246 15977 34298
rect 15977 34246 16007 34298
rect 16031 34246 16041 34298
rect 16041 34246 16087 34298
rect 15791 34244 15847 34246
rect 15871 34244 15927 34246
rect 15951 34244 16007 34246
rect 16031 34244 16087 34246
rect 15791 33210 15847 33212
rect 15871 33210 15927 33212
rect 15951 33210 16007 33212
rect 16031 33210 16087 33212
rect 15791 33158 15837 33210
rect 15837 33158 15847 33210
rect 15871 33158 15901 33210
rect 15901 33158 15913 33210
rect 15913 33158 15927 33210
rect 15951 33158 15965 33210
rect 15965 33158 15977 33210
rect 15977 33158 16007 33210
rect 16031 33158 16041 33210
rect 16041 33158 16087 33210
rect 15791 33156 15847 33158
rect 15871 33156 15927 33158
rect 15951 33156 16007 33158
rect 16031 33156 16087 33158
rect 15791 32122 15847 32124
rect 15871 32122 15927 32124
rect 15951 32122 16007 32124
rect 16031 32122 16087 32124
rect 15791 32070 15837 32122
rect 15837 32070 15847 32122
rect 15871 32070 15901 32122
rect 15901 32070 15913 32122
rect 15913 32070 15927 32122
rect 15951 32070 15965 32122
rect 15965 32070 15977 32122
rect 15977 32070 16007 32122
rect 16031 32070 16041 32122
rect 16041 32070 16087 32122
rect 15791 32068 15847 32070
rect 15871 32068 15927 32070
rect 15951 32068 16007 32070
rect 16031 32068 16087 32070
rect 15750 31184 15806 31240
rect 16026 31728 16082 31784
rect 15791 31034 15847 31036
rect 15871 31034 15927 31036
rect 15951 31034 16007 31036
rect 16031 31034 16087 31036
rect 15791 30982 15837 31034
rect 15837 30982 15847 31034
rect 15871 30982 15901 31034
rect 15901 30982 15913 31034
rect 15913 30982 15927 31034
rect 15951 30982 15965 31034
rect 15965 30982 15977 31034
rect 15977 30982 16007 31034
rect 16031 30982 16041 31034
rect 16041 30982 16087 31034
rect 15791 30980 15847 30982
rect 15871 30980 15927 30982
rect 15951 30980 16007 30982
rect 16031 30980 16087 30982
rect 15791 29946 15847 29948
rect 15871 29946 15927 29948
rect 15951 29946 16007 29948
rect 16031 29946 16087 29948
rect 15791 29894 15837 29946
rect 15837 29894 15847 29946
rect 15871 29894 15901 29946
rect 15901 29894 15913 29946
rect 15913 29894 15927 29946
rect 15951 29894 15965 29946
rect 15965 29894 15977 29946
rect 15977 29894 16007 29946
rect 16031 29894 16041 29946
rect 16041 29894 16087 29946
rect 15791 29892 15847 29894
rect 15871 29892 15927 29894
rect 15951 29892 16007 29894
rect 16031 29892 16087 29894
rect 15842 29280 15898 29336
rect 15791 28858 15847 28860
rect 15871 28858 15927 28860
rect 15951 28858 16007 28860
rect 16031 28858 16087 28860
rect 15791 28806 15837 28858
rect 15837 28806 15847 28858
rect 15871 28806 15901 28858
rect 15901 28806 15913 28858
rect 15913 28806 15927 28858
rect 15951 28806 15965 28858
rect 15965 28806 15977 28858
rect 15977 28806 16007 28858
rect 16031 28806 16041 28858
rect 16041 28806 16087 28858
rect 15791 28804 15847 28806
rect 15871 28804 15927 28806
rect 15951 28804 16007 28806
rect 16031 28804 16087 28806
rect 15791 27770 15847 27772
rect 15871 27770 15927 27772
rect 15951 27770 16007 27772
rect 16031 27770 16087 27772
rect 15791 27718 15837 27770
rect 15837 27718 15847 27770
rect 15871 27718 15901 27770
rect 15901 27718 15913 27770
rect 15913 27718 15927 27770
rect 15951 27718 15965 27770
rect 15965 27718 15977 27770
rect 15977 27718 16007 27770
rect 16031 27718 16041 27770
rect 16041 27718 16087 27770
rect 15791 27716 15847 27718
rect 15871 27716 15927 27718
rect 15951 27716 16007 27718
rect 16031 27716 16087 27718
rect 15791 26682 15847 26684
rect 15871 26682 15927 26684
rect 15951 26682 16007 26684
rect 16031 26682 16087 26684
rect 15791 26630 15837 26682
rect 15837 26630 15847 26682
rect 15871 26630 15901 26682
rect 15901 26630 15913 26682
rect 15913 26630 15927 26682
rect 15951 26630 15965 26682
rect 15965 26630 15977 26682
rect 15977 26630 16007 26682
rect 16031 26630 16041 26682
rect 16041 26630 16087 26682
rect 15791 26628 15847 26630
rect 15871 26628 15927 26630
rect 15951 26628 16007 26630
rect 16031 26628 16087 26630
rect 14554 17176 14610 17232
rect 14094 16088 14150 16144
rect 13634 9832 13690 9888
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 13082 4936 13138 4992
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 13358 6180 13414 6216
rect 13358 6160 13360 6180
rect 13360 6160 13412 6180
rect 13412 6160 13414 6180
rect 13174 4120 13230 4176
rect 12346 3848 12402 3904
rect 12898 3712 12954 3768
rect 13450 6024 13506 6080
rect 13818 9696 13874 9752
rect 13726 6316 13782 6352
rect 13726 6296 13728 6316
rect 13728 6296 13780 6316
rect 13780 6296 13782 6316
rect 13726 5480 13782 5536
rect 13450 5208 13506 5264
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 13818 5208 13874 5264
rect 13542 2388 13544 2408
rect 13544 2388 13596 2408
rect 13596 2388 13598 2408
rect 13542 2352 13598 2388
rect 13818 2624 13874 2680
rect 13818 1808 13874 1864
rect 14278 13932 14334 13968
rect 14278 13912 14280 13932
rect 14280 13912 14332 13932
rect 14332 13912 14334 13932
rect 15014 17992 15070 18048
rect 15014 16632 15070 16688
rect 14370 8916 14372 8936
rect 14372 8916 14424 8936
rect 14424 8916 14426 8936
rect 14370 8880 14426 8916
rect 14922 12008 14978 12064
rect 14922 9016 14978 9072
rect 14738 5908 14794 5944
rect 14738 5888 14740 5908
rect 14740 5888 14792 5908
rect 14792 5888 14794 5908
rect 14370 4684 14426 4720
rect 14370 4664 14372 4684
rect 14372 4664 14424 4684
rect 14424 4664 14426 4684
rect 14922 4936 14978 4992
rect 14922 4564 14924 4584
rect 14924 4564 14976 4584
rect 14976 4564 14978 4584
rect 14922 4528 14978 4564
rect 14278 2352 14334 2408
rect 14186 1944 14242 2000
rect 15934 25880 15990 25936
rect 15791 25594 15847 25596
rect 15871 25594 15927 25596
rect 15951 25594 16007 25596
rect 16031 25594 16087 25596
rect 15791 25542 15837 25594
rect 15837 25542 15847 25594
rect 15871 25542 15901 25594
rect 15901 25542 15913 25594
rect 15913 25542 15927 25594
rect 15951 25542 15965 25594
rect 15965 25542 15977 25594
rect 15977 25542 16007 25594
rect 16031 25542 16041 25594
rect 16041 25542 16087 25594
rect 15791 25540 15847 25542
rect 15871 25540 15927 25542
rect 15951 25540 16007 25542
rect 16031 25540 16087 25542
rect 15934 25200 15990 25256
rect 16210 27532 16266 27568
rect 16210 27512 16212 27532
rect 16212 27512 16264 27532
rect 16264 27512 16266 27532
rect 16118 25064 16174 25120
rect 15791 24506 15847 24508
rect 15871 24506 15927 24508
rect 15951 24506 16007 24508
rect 16031 24506 16087 24508
rect 15791 24454 15837 24506
rect 15837 24454 15847 24506
rect 15871 24454 15901 24506
rect 15901 24454 15913 24506
rect 15913 24454 15927 24506
rect 15951 24454 15965 24506
rect 15965 24454 15977 24506
rect 15977 24454 16007 24506
rect 16031 24454 16041 24506
rect 16041 24454 16087 24506
rect 15791 24452 15847 24454
rect 15871 24452 15927 24454
rect 15951 24452 16007 24454
rect 16031 24452 16087 24454
rect 15791 23418 15847 23420
rect 15871 23418 15927 23420
rect 15951 23418 16007 23420
rect 16031 23418 16087 23420
rect 15791 23366 15837 23418
rect 15837 23366 15847 23418
rect 15871 23366 15901 23418
rect 15901 23366 15913 23418
rect 15913 23366 15927 23418
rect 15951 23366 15965 23418
rect 15965 23366 15977 23418
rect 15977 23366 16007 23418
rect 16031 23366 16041 23418
rect 16041 23366 16087 23418
rect 15791 23364 15847 23366
rect 15871 23364 15927 23366
rect 15951 23364 16007 23366
rect 16031 23364 16087 23366
rect 15791 22330 15847 22332
rect 15871 22330 15927 22332
rect 15951 22330 16007 22332
rect 16031 22330 16087 22332
rect 15791 22278 15837 22330
rect 15837 22278 15847 22330
rect 15871 22278 15901 22330
rect 15901 22278 15913 22330
rect 15913 22278 15927 22330
rect 15951 22278 15965 22330
rect 15965 22278 15977 22330
rect 15977 22278 16007 22330
rect 16031 22278 16041 22330
rect 16041 22278 16087 22330
rect 15791 22276 15847 22278
rect 15871 22276 15927 22278
rect 15951 22276 16007 22278
rect 16031 22276 16087 22278
rect 15750 22072 15806 22128
rect 15791 21242 15847 21244
rect 15871 21242 15927 21244
rect 15951 21242 16007 21244
rect 16031 21242 16087 21244
rect 15791 21190 15837 21242
rect 15837 21190 15847 21242
rect 15871 21190 15901 21242
rect 15901 21190 15913 21242
rect 15913 21190 15927 21242
rect 15951 21190 15965 21242
rect 15965 21190 15977 21242
rect 15977 21190 16007 21242
rect 16031 21190 16041 21242
rect 16041 21190 16087 21242
rect 15791 21188 15847 21190
rect 15871 21188 15927 21190
rect 15951 21188 16007 21190
rect 16031 21188 16087 21190
rect 15791 20154 15847 20156
rect 15871 20154 15927 20156
rect 15951 20154 16007 20156
rect 16031 20154 16087 20156
rect 15791 20102 15837 20154
rect 15837 20102 15847 20154
rect 15871 20102 15901 20154
rect 15901 20102 15913 20154
rect 15913 20102 15927 20154
rect 15951 20102 15965 20154
rect 15965 20102 15977 20154
rect 15977 20102 16007 20154
rect 16031 20102 16041 20154
rect 16041 20102 16087 20154
rect 15791 20100 15847 20102
rect 15871 20100 15927 20102
rect 15951 20100 16007 20102
rect 16031 20100 16087 20102
rect 16946 41656 17002 41712
rect 17314 41792 17370 41848
rect 17038 41520 17094 41576
rect 18758 43546 18814 43548
rect 18838 43546 18894 43548
rect 18918 43546 18974 43548
rect 18998 43546 19054 43548
rect 18758 43494 18804 43546
rect 18804 43494 18814 43546
rect 18838 43494 18868 43546
rect 18868 43494 18880 43546
rect 18880 43494 18894 43546
rect 18918 43494 18932 43546
rect 18932 43494 18944 43546
rect 18944 43494 18974 43546
rect 18998 43494 19008 43546
rect 19008 43494 19054 43546
rect 18758 43492 18814 43494
rect 18838 43492 18894 43494
rect 18918 43492 18974 43494
rect 18998 43492 19054 43494
rect 18418 42608 18474 42664
rect 17682 41656 17738 41712
rect 17038 33924 17094 33960
rect 17038 33904 17040 33924
rect 17040 33904 17092 33924
rect 17092 33904 17094 33924
rect 16762 29552 16818 29608
rect 16578 27648 16634 27704
rect 16486 27276 16488 27296
rect 16488 27276 16540 27296
rect 16540 27276 16542 27296
rect 16486 27240 16542 27276
rect 16486 25880 16542 25936
rect 16854 29416 16910 29472
rect 16486 21528 16542 21584
rect 17130 27920 17186 27976
rect 17774 34040 17830 34096
rect 17958 33224 18014 33280
rect 17590 29280 17646 29336
rect 17498 28056 17554 28112
rect 17314 27532 17370 27568
rect 17314 27512 17316 27532
rect 17316 27512 17368 27532
rect 17368 27512 17370 27532
rect 17222 27412 17224 27432
rect 17224 27412 17276 27432
rect 17276 27412 17278 27432
rect 17222 27376 17278 27412
rect 17314 26696 17370 26752
rect 16854 21800 16910 21856
rect 16486 21392 16542 21448
rect 16210 19352 16266 19408
rect 15791 19066 15847 19068
rect 15871 19066 15927 19068
rect 15951 19066 16007 19068
rect 16031 19066 16087 19068
rect 15791 19014 15837 19066
rect 15837 19014 15847 19066
rect 15871 19014 15901 19066
rect 15901 19014 15913 19066
rect 15913 19014 15927 19066
rect 15951 19014 15965 19066
rect 15965 19014 15977 19066
rect 15977 19014 16007 19066
rect 16031 19014 16041 19066
rect 16041 19014 16087 19066
rect 15791 19012 15847 19014
rect 15871 19012 15927 19014
rect 15951 19012 16007 19014
rect 16031 19012 16087 19014
rect 16210 18708 16212 18728
rect 16212 18708 16264 18728
rect 16264 18708 16266 18728
rect 15566 17992 15622 18048
rect 16210 18672 16266 18708
rect 15791 17978 15847 17980
rect 15871 17978 15927 17980
rect 15951 17978 16007 17980
rect 16031 17978 16087 17980
rect 15791 17926 15837 17978
rect 15837 17926 15847 17978
rect 15871 17926 15901 17978
rect 15901 17926 15913 17978
rect 15913 17926 15927 17978
rect 15951 17926 15965 17978
rect 15965 17926 15977 17978
rect 15977 17926 16007 17978
rect 16031 17926 16041 17978
rect 16041 17926 16087 17978
rect 15791 17924 15847 17926
rect 15871 17924 15927 17926
rect 15951 17924 16007 17926
rect 16031 17924 16087 17926
rect 15791 16890 15847 16892
rect 15871 16890 15927 16892
rect 15951 16890 16007 16892
rect 16031 16890 16087 16892
rect 15791 16838 15837 16890
rect 15837 16838 15847 16890
rect 15871 16838 15901 16890
rect 15901 16838 15913 16890
rect 15913 16838 15927 16890
rect 15951 16838 15965 16890
rect 15965 16838 15977 16890
rect 15977 16838 16007 16890
rect 16031 16838 16041 16890
rect 16041 16838 16087 16890
rect 15791 16836 15847 16838
rect 15871 16836 15927 16838
rect 15951 16836 16007 16838
rect 16031 16836 16087 16838
rect 16302 17856 16358 17912
rect 15290 14456 15346 14512
rect 15198 13368 15254 13424
rect 15198 10240 15254 10296
rect 15290 6976 15346 7032
rect 16026 16496 16082 16552
rect 15791 15802 15847 15804
rect 15871 15802 15927 15804
rect 15951 15802 16007 15804
rect 16031 15802 16087 15804
rect 15791 15750 15837 15802
rect 15837 15750 15847 15802
rect 15871 15750 15901 15802
rect 15901 15750 15913 15802
rect 15913 15750 15927 15802
rect 15951 15750 15965 15802
rect 15965 15750 15977 15802
rect 15977 15750 16007 15802
rect 16031 15750 16041 15802
rect 16041 15750 16087 15802
rect 15791 15748 15847 15750
rect 15871 15748 15927 15750
rect 15951 15748 16007 15750
rect 16031 15748 16087 15750
rect 15791 14714 15847 14716
rect 15871 14714 15927 14716
rect 15951 14714 16007 14716
rect 16031 14714 16087 14716
rect 15791 14662 15837 14714
rect 15837 14662 15847 14714
rect 15871 14662 15901 14714
rect 15901 14662 15913 14714
rect 15913 14662 15927 14714
rect 15951 14662 15965 14714
rect 15965 14662 15977 14714
rect 15977 14662 16007 14714
rect 16031 14662 16041 14714
rect 16041 14662 16087 14714
rect 15791 14660 15847 14662
rect 15871 14660 15927 14662
rect 15951 14660 16007 14662
rect 16031 14660 16087 14662
rect 16210 14592 16266 14648
rect 16026 14476 16082 14512
rect 16026 14456 16028 14476
rect 16028 14456 16080 14476
rect 16080 14456 16082 14476
rect 15791 13626 15847 13628
rect 15871 13626 15927 13628
rect 15951 13626 16007 13628
rect 16031 13626 16087 13628
rect 15791 13574 15837 13626
rect 15837 13574 15847 13626
rect 15871 13574 15901 13626
rect 15901 13574 15913 13626
rect 15913 13574 15927 13626
rect 15951 13574 15965 13626
rect 15965 13574 15977 13626
rect 15977 13574 16007 13626
rect 16031 13574 16041 13626
rect 16041 13574 16087 13626
rect 15791 13572 15847 13574
rect 15871 13572 15927 13574
rect 15951 13572 16007 13574
rect 16031 13572 16087 13574
rect 15791 12538 15847 12540
rect 15871 12538 15927 12540
rect 15951 12538 16007 12540
rect 16031 12538 16087 12540
rect 15791 12486 15837 12538
rect 15837 12486 15847 12538
rect 15871 12486 15901 12538
rect 15901 12486 15913 12538
rect 15913 12486 15927 12538
rect 15951 12486 15965 12538
rect 15965 12486 15977 12538
rect 15977 12486 16007 12538
rect 16031 12486 16041 12538
rect 16041 12486 16087 12538
rect 15791 12484 15847 12486
rect 15871 12484 15927 12486
rect 15951 12484 16007 12486
rect 16031 12484 16087 12486
rect 15842 12008 15898 12064
rect 15791 11450 15847 11452
rect 15871 11450 15927 11452
rect 15951 11450 16007 11452
rect 16031 11450 16087 11452
rect 15791 11398 15837 11450
rect 15837 11398 15847 11450
rect 15871 11398 15901 11450
rect 15901 11398 15913 11450
rect 15913 11398 15927 11450
rect 15951 11398 15965 11450
rect 15965 11398 15977 11450
rect 15977 11398 16007 11450
rect 16031 11398 16041 11450
rect 16041 11398 16087 11450
rect 15791 11396 15847 11398
rect 15871 11396 15927 11398
rect 15951 11396 16007 11398
rect 16031 11396 16087 11398
rect 16302 14456 16358 14512
rect 16578 15544 16634 15600
rect 15791 10362 15847 10364
rect 15871 10362 15927 10364
rect 15951 10362 16007 10364
rect 16031 10362 16087 10364
rect 15791 10310 15837 10362
rect 15837 10310 15847 10362
rect 15871 10310 15901 10362
rect 15901 10310 15913 10362
rect 15913 10310 15927 10362
rect 15951 10310 15965 10362
rect 15965 10310 15977 10362
rect 15977 10310 16007 10362
rect 16031 10310 16041 10362
rect 16041 10310 16087 10362
rect 15791 10308 15847 10310
rect 15871 10308 15927 10310
rect 15951 10308 16007 10310
rect 16031 10308 16087 10310
rect 15658 9560 15714 9616
rect 15791 9274 15847 9276
rect 15871 9274 15927 9276
rect 15951 9274 16007 9276
rect 16031 9274 16087 9276
rect 15791 9222 15837 9274
rect 15837 9222 15847 9274
rect 15871 9222 15901 9274
rect 15901 9222 15913 9274
rect 15913 9222 15927 9274
rect 15951 9222 15965 9274
rect 15965 9222 15977 9274
rect 15977 9222 16007 9274
rect 16031 9222 16041 9274
rect 16041 9222 16087 9274
rect 15791 9220 15847 9222
rect 15871 9220 15927 9222
rect 15951 9220 16007 9222
rect 16031 9220 16087 9222
rect 15750 9016 15806 9072
rect 17314 24148 17316 24168
rect 17316 24148 17368 24168
rect 17368 24148 17370 24168
rect 17314 24112 17370 24148
rect 17590 25608 17646 25664
rect 17590 25236 17592 25256
rect 17592 25236 17644 25256
rect 17644 25236 17646 25256
rect 17590 25200 17646 25236
rect 16762 14456 16818 14512
rect 16762 14184 16818 14240
rect 15791 8186 15847 8188
rect 15871 8186 15927 8188
rect 15951 8186 16007 8188
rect 16031 8186 16087 8188
rect 15791 8134 15837 8186
rect 15837 8134 15847 8186
rect 15871 8134 15901 8186
rect 15901 8134 15913 8186
rect 15913 8134 15927 8186
rect 15951 8134 15965 8186
rect 15965 8134 15977 8186
rect 15977 8134 16007 8186
rect 16031 8134 16041 8186
rect 16041 8134 16087 8186
rect 15791 8132 15847 8134
rect 15871 8132 15927 8134
rect 15951 8132 16007 8134
rect 16031 8132 16087 8134
rect 15658 7656 15714 7712
rect 15566 6296 15622 6352
rect 15198 5072 15254 5128
rect 15791 7098 15847 7100
rect 15871 7098 15927 7100
rect 15951 7098 16007 7100
rect 16031 7098 16087 7100
rect 15791 7046 15837 7098
rect 15837 7046 15847 7098
rect 15871 7046 15901 7098
rect 15901 7046 15913 7098
rect 15913 7046 15927 7098
rect 15951 7046 15965 7098
rect 15965 7046 15977 7098
rect 15977 7046 16007 7098
rect 16031 7046 16041 7098
rect 16041 7046 16087 7098
rect 15791 7044 15847 7046
rect 15871 7044 15927 7046
rect 15951 7044 16007 7046
rect 16031 7044 16087 7046
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 16210 7928 16266 7984
rect 16394 5616 16450 5672
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 16302 2624 16358 2680
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 17314 21120 17370 21176
rect 17130 14864 17186 14920
rect 17222 14476 17278 14512
rect 17222 14456 17224 14476
rect 17224 14456 17276 14476
rect 17276 14456 17278 14476
rect 17038 11228 17040 11248
rect 17040 11228 17092 11248
rect 17092 11228 17094 11248
rect 17038 11192 17094 11228
rect 17774 21548 17830 21584
rect 17774 21528 17776 21548
rect 17776 21528 17828 21548
rect 17828 21528 17830 21548
rect 17958 21664 18014 21720
rect 19246 43016 19302 43072
rect 18878 42608 18934 42664
rect 18758 42458 18814 42460
rect 18838 42458 18894 42460
rect 18918 42458 18974 42460
rect 18998 42458 19054 42460
rect 18758 42406 18804 42458
rect 18804 42406 18814 42458
rect 18838 42406 18868 42458
rect 18868 42406 18880 42458
rect 18880 42406 18894 42458
rect 18918 42406 18932 42458
rect 18932 42406 18944 42458
rect 18944 42406 18974 42458
rect 18998 42406 19008 42458
rect 19008 42406 19054 42458
rect 18758 42404 18814 42406
rect 18838 42404 18894 42406
rect 18918 42404 18974 42406
rect 18998 42404 19054 42406
rect 18970 42200 19026 42256
rect 18326 41656 18382 41712
rect 18234 41556 18236 41576
rect 18236 41556 18288 41576
rect 18288 41556 18290 41576
rect 18234 41520 18290 41556
rect 18418 41420 18420 41440
rect 18420 41420 18472 41440
rect 18472 41420 18474 41440
rect 18418 41384 18474 41420
rect 18418 41112 18474 41168
rect 18326 35808 18382 35864
rect 17314 10104 17370 10160
rect 16670 6840 16726 6896
rect 17222 5208 17278 5264
rect 17038 4800 17094 4856
rect 17222 3848 17278 3904
rect 17590 9968 17646 10024
rect 17498 5752 17554 5808
rect 17406 5480 17462 5536
rect 18142 21392 18198 21448
rect 18418 33224 18474 33280
rect 19246 42200 19302 42256
rect 18758 41370 18814 41372
rect 18838 41370 18894 41372
rect 18918 41370 18974 41372
rect 18998 41370 19054 41372
rect 18758 41318 18804 41370
rect 18804 41318 18814 41370
rect 18838 41318 18868 41370
rect 18868 41318 18880 41370
rect 18880 41318 18894 41370
rect 18918 41318 18932 41370
rect 18932 41318 18944 41370
rect 18944 41318 18974 41370
rect 18998 41318 19008 41370
rect 19008 41318 19054 41370
rect 18758 41316 18814 41318
rect 18838 41316 18894 41318
rect 18918 41316 18974 41318
rect 18998 41316 19054 41318
rect 19522 41656 19578 41712
rect 19706 41520 19762 41576
rect 19798 41268 19854 41304
rect 19798 41248 19800 41268
rect 19800 41248 19852 41268
rect 19852 41248 19854 41268
rect 18758 40282 18814 40284
rect 18838 40282 18894 40284
rect 18918 40282 18974 40284
rect 18998 40282 19054 40284
rect 18758 40230 18804 40282
rect 18804 40230 18814 40282
rect 18838 40230 18868 40282
rect 18868 40230 18880 40282
rect 18880 40230 18894 40282
rect 18918 40230 18932 40282
rect 18932 40230 18944 40282
rect 18944 40230 18974 40282
rect 18998 40230 19008 40282
rect 19008 40230 19054 40282
rect 18758 40228 18814 40230
rect 18838 40228 18894 40230
rect 18918 40228 18974 40230
rect 18998 40228 19054 40230
rect 18758 39194 18814 39196
rect 18838 39194 18894 39196
rect 18918 39194 18974 39196
rect 18998 39194 19054 39196
rect 18758 39142 18804 39194
rect 18804 39142 18814 39194
rect 18838 39142 18868 39194
rect 18868 39142 18880 39194
rect 18880 39142 18894 39194
rect 18918 39142 18932 39194
rect 18932 39142 18944 39194
rect 18944 39142 18974 39194
rect 18998 39142 19008 39194
rect 19008 39142 19054 39194
rect 18758 39140 18814 39142
rect 18838 39140 18894 39142
rect 18918 39140 18974 39142
rect 18998 39140 19054 39142
rect 19430 38664 19486 38720
rect 18758 38106 18814 38108
rect 18838 38106 18894 38108
rect 18918 38106 18974 38108
rect 18998 38106 19054 38108
rect 18758 38054 18804 38106
rect 18804 38054 18814 38106
rect 18838 38054 18868 38106
rect 18868 38054 18880 38106
rect 18880 38054 18894 38106
rect 18918 38054 18932 38106
rect 18932 38054 18944 38106
rect 18944 38054 18974 38106
rect 18998 38054 19008 38106
rect 19008 38054 19054 38106
rect 18758 38052 18814 38054
rect 18838 38052 18894 38054
rect 18918 38052 18974 38054
rect 18998 38052 19054 38054
rect 18758 37018 18814 37020
rect 18838 37018 18894 37020
rect 18918 37018 18974 37020
rect 18998 37018 19054 37020
rect 18758 36966 18804 37018
rect 18804 36966 18814 37018
rect 18838 36966 18868 37018
rect 18868 36966 18880 37018
rect 18880 36966 18894 37018
rect 18918 36966 18932 37018
rect 18932 36966 18944 37018
rect 18944 36966 18974 37018
rect 18998 36966 19008 37018
rect 19008 36966 19054 37018
rect 18758 36964 18814 36966
rect 18838 36964 18894 36966
rect 18918 36964 18974 36966
rect 18998 36964 19054 36966
rect 18758 35930 18814 35932
rect 18838 35930 18894 35932
rect 18918 35930 18974 35932
rect 18998 35930 19054 35932
rect 18758 35878 18804 35930
rect 18804 35878 18814 35930
rect 18838 35878 18868 35930
rect 18868 35878 18880 35930
rect 18880 35878 18894 35930
rect 18918 35878 18932 35930
rect 18932 35878 18944 35930
rect 18944 35878 18974 35930
rect 18998 35878 19008 35930
rect 19008 35878 19054 35930
rect 18758 35876 18814 35878
rect 18838 35876 18894 35878
rect 18918 35876 18974 35878
rect 18998 35876 19054 35878
rect 18758 34842 18814 34844
rect 18838 34842 18894 34844
rect 18918 34842 18974 34844
rect 18998 34842 19054 34844
rect 18758 34790 18804 34842
rect 18804 34790 18814 34842
rect 18838 34790 18868 34842
rect 18868 34790 18880 34842
rect 18880 34790 18894 34842
rect 18918 34790 18932 34842
rect 18932 34790 18944 34842
rect 18944 34790 18974 34842
rect 18998 34790 19008 34842
rect 19008 34790 19054 34842
rect 18758 34788 18814 34790
rect 18838 34788 18894 34790
rect 18918 34788 18974 34790
rect 18998 34788 19054 34790
rect 18970 34448 19026 34504
rect 18758 33754 18814 33756
rect 18838 33754 18894 33756
rect 18918 33754 18974 33756
rect 18998 33754 19054 33756
rect 18758 33702 18804 33754
rect 18804 33702 18814 33754
rect 18838 33702 18868 33754
rect 18868 33702 18880 33754
rect 18880 33702 18894 33754
rect 18918 33702 18932 33754
rect 18932 33702 18944 33754
rect 18944 33702 18974 33754
rect 18998 33702 19008 33754
rect 19008 33702 19054 33754
rect 18758 33700 18814 33702
rect 18838 33700 18894 33702
rect 18918 33700 18974 33702
rect 18998 33700 19054 33702
rect 18970 33532 18972 33552
rect 18972 33532 19024 33552
rect 19024 33532 19026 33552
rect 18970 33496 19026 33532
rect 18758 32666 18814 32668
rect 18838 32666 18894 32668
rect 18918 32666 18974 32668
rect 18998 32666 19054 32668
rect 18758 32614 18804 32666
rect 18804 32614 18814 32666
rect 18838 32614 18868 32666
rect 18868 32614 18880 32666
rect 18880 32614 18894 32666
rect 18918 32614 18932 32666
rect 18932 32614 18944 32666
rect 18944 32614 18974 32666
rect 18998 32614 19008 32666
rect 19008 32614 19054 32666
rect 18758 32612 18814 32614
rect 18838 32612 18894 32614
rect 18918 32612 18974 32614
rect 18998 32612 19054 32614
rect 19338 33360 19394 33416
rect 18758 31578 18814 31580
rect 18838 31578 18894 31580
rect 18918 31578 18974 31580
rect 18998 31578 19054 31580
rect 18758 31526 18804 31578
rect 18804 31526 18814 31578
rect 18838 31526 18868 31578
rect 18868 31526 18880 31578
rect 18880 31526 18894 31578
rect 18918 31526 18932 31578
rect 18932 31526 18944 31578
rect 18944 31526 18974 31578
rect 18998 31526 19008 31578
rect 19008 31526 19054 31578
rect 18758 31524 18814 31526
rect 18838 31524 18894 31526
rect 18918 31524 18974 31526
rect 18998 31524 19054 31526
rect 18758 30490 18814 30492
rect 18838 30490 18894 30492
rect 18918 30490 18974 30492
rect 18998 30490 19054 30492
rect 18758 30438 18804 30490
rect 18804 30438 18814 30490
rect 18838 30438 18868 30490
rect 18868 30438 18880 30490
rect 18880 30438 18894 30490
rect 18918 30438 18932 30490
rect 18932 30438 18944 30490
rect 18944 30438 18974 30490
rect 18998 30438 19008 30490
rect 19008 30438 19054 30490
rect 18758 30436 18814 30438
rect 18838 30436 18894 30438
rect 18918 30436 18974 30438
rect 18998 30436 19054 30438
rect 19798 39072 19854 39128
rect 20074 42200 20130 42256
rect 20626 42200 20682 42256
rect 20718 41384 20774 41440
rect 20074 39908 20130 39944
rect 20074 39888 20076 39908
rect 20076 39888 20128 39908
rect 20128 39888 20130 39908
rect 20258 40296 20314 40352
rect 19706 33088 19762 33144
rect 18758 29402 18814 29404
rect 18838 29402 18894 29404
rect 18918 29402 18974 29404
rect 18998 29402 19054 29404
rect 18758 29350 18804 29402
rect 18804 29350 18814 29402
rect 18838 29350 18868 29402
rect 18868 29350 18880 29402
rect 18880 29350 18894 29402
rect 18918 29350 18932 29402
rect 18932 29350 18944 29402
rect 18944 29350 18974 29402
rect 18998 29350 19008 29402
rect 19008 29350 19054 29402
rect 18758 29348 18814 29350
rect 18838 29348 18894 29350
rect 18918 29348 18974 29350
rect 18998 29348 19054 29350
rect 18758 28314 18814 28316
rect 18838 28314 18894 28316
rect 18918 28314 18974 28316
rect 18998 28314 19054 28316
rect 18758 28262 18804 28314
rect 18804 28262 18814 28314
rect 18838 28262 18868 28314
rect 18868 28262 18880 28314
rect 18880 28262 18894 28314
rect 18918 28262 18932 28314
rect 18932 28262 18944 28314
rect 18944 28262 18974 28314
rect 18998 28262 19008 28314
rect 19008 28262 19054 28314
rect 18758 28260 18814 28262
rect 18838 28260 18894 28262
rect 18918 28260 18974 28262
rect 18998 28260 19054 28262
rect 18758 27226 18814 27228
rect 18838 27226 18894 27228
rect 18918 27226 18974 27228
rect 18998 27226 19054 27228
rect 18758 27174 18804 27226
rect 18804 27174 18814 27226
rect 18838 27174 18868 27226
rect 18868 27174 18880 27226
rect 18880 27174 18894 27226
rect 18918 27174 18932 27226
rect 18932 27174 18944 27226
rect 18944 27174 18974 27226
rect 18998 27174 19008 27226
rect 19008 27174 19054 27226
rect 18758 27172 18814 27174
rect 18838 27172 18894 27174
rect 18918 27172 18974 27174
rect 18998 27172 19054 27174
rect 18694 26444 18750 26480
rect 18694 26424 18696 26444
rect 18696 26424 18748 26444
rect 18748 26424 18750 26444
rect 18758 26138 18814 26140
rect 18838 26138 18894 26140
rect 18918 26138 18974 26140
rect 18998 26138 19054 26140
rect 18758 26086 18804 26138
rect 18804 26086 18814 26138
rect 18838 26086 18868 26138
rect 18868 26086 18880 26138
rect 18880 26086 18894 26138
rect 18918 26086 18932 26138
rect 18932 26086 18944 26138
rect 18944 26086 18974 26138
rect 18998 26086 19008 26138
rect 19008 26086 19054 26138
rect 18758 26084 18814 26086
rect 18838 26084 18894 26086
rect 18918 26084 18974 26086
rect 18998 26084 19054 26086
rect 18758 25050 18814 25052
rect 18838 25050 18894 25052
rect 18918 25050 18974 25052
rect 18998 25050 19054 25052
rect 18758 24998 18804 25050
rect 18804 24998 18814 25050
rect 18838 24998 18868 25050
rect 18868 24998 18880 25050
rect 18880 24998 18894 25050
rect 18918 24998 18932 25050
rect 18932 24998 18944 25050
rect 18944 24998 18974 25050
rect 18998 24998 19008 25050
rect 19008 24998 19054 25050
rect 18758 24996 18814 24998
rect 18838 24996 18894 24998
rect 18918 24996 18974 24998
rect 18998 24996 19054 24998
rect 18758 23962 18814 23964
rect 18838 23962 18894 23964
rect 18918 23962 18974 23964
rect 18998 23962 19054 23964
rect 18758 23910 18804 23962
rect 18804 23910 18814 23962
rect 18838 23910 18868 23962
rect 18868 23910 18880 23962
rect 18880 23910 18894 23962
rect 18918 23910 18932 23962
rect 18932 23910 18944 23962
rect 18944 23910 18974 23962
rect 18998 23910 19008 23962
rect 19008 23910 19054 23962
rect 18758 23908 18814 23910
rect 18838 23908 18894 23910
rect 18918 23908 18974 23910
rect 18998 23908 19054 23910
rect 18758 22874 18814 22876
rect 18838 22874 18894 22876
rect 18918 22874 18974 22876
rect 18998 22874 19054 22876
rect 18758 22822 18804 22874
rect 18804 22822 18814 22874
rect 18838 22822 18868 22874
rect 18868 22822 18880 22874
rect 18880 22822 18894 22874
rect 18918 22822 18932 22874
rect 18932 22822 18944 22874
rect 18944 22822 18974 22874
rect 18998 22822 19008 22874
rect 19008 22822 19054 22874
rect 18758 22820 18814 22822
rect 18838 22820 18894 22822
rect 18918 22820 18974 22822
rect 18998 22820 19054 22822
rect 18418 22072 18474 22128
rect 18418 21800 18474 21856
rect 18326 21664 18382 21720
rect 18234 17176 18290 17232
rect 18326 12144 18382 12200
rect 18234 11736 18290 11792
rect 18326 8492 18382 8528
rect 18326 8472 18328 8492
rect 18328 8472 18380 8492
rect 18380 8472 18382 8492
rect 18758 21786 18814 21788
rect 18838 21786 18894 21788
rect 18918 21786 18974 21788
rect 18998 21786 19054 21788
rect 18758 21734 18804 21786
rect 18804 21734 18814 21786
rect 18838 21734 18868 21786
rect 18868 21734 18880 21786
rect 18880 21734 18894 21786
rect 18918 21734 18932 21786
rect 18932 21734 18944 21786
rect 18944 21734 18974 21786
rect 18998 21734 19008 21786
rect 19008 21734 19054 21786
rect 18758 21732 18814 21734
rect 18838 21732 18894 21734
rect 18918 21732 18974 21734
rect 18998 21732 19054 21734
rect 19154 21120 19210 21176
rect 18758 20698 18814 20700
rect 18838 20698 18894 20700
rect 18918 20698 18974 20700
rect 18998 20698 19054 20700
rect 18758 20646 18804 20698
rect 18804 20646 18814 20698
rect 18838 20646 18868 20698
rect 18868 20646 18880 20698
rect 18880 20646 18894 20698
rect 18918 20646 18932 20698
rect 18932 20646 18944 20698
rect 18944 20646 18974 20698
rect 18998 20646 19008 20698
rect 19008 20646 19054 20698
rect 18758 20644 18814 20646
rect 18838 20644 18894 20646
rect 18918 20644 18974 20646
rect 18998 20644 19054 20646
rect 19614 24520 19670 24576
rect 19522 23568 19578 23624
rect 19338 20712 19394 20768
rect 18758 19610 18814 19612
rect 18838 19610 18894 19612
rect 18918 19610 18974 19612
rect 18998 19610 19054 19612
rect 18758 19558 18804 19610
rect 18804 19558 18814 19610
rect 18838 19558 18868 19610
rect 18868 19558 18880 19610
rect 18880 19558 18894 19610
rect 18918 19558 18932 19610
rect 18932 19558 18944 19610
rect 18944 19558 18974 19610
rect 18998 19558 19008 19610
rect 19008 19558 19054 19610
rect 18758 19556 18814 19558
rect 18838 19556 18894 19558
rect 18918 19556 18974 19558
rect 18998 19556 19054 19558
rect 18758 18522 18814 18524
rect 18838 18522 18894 18524
rect 18918 18522 18974 18524
rect 18998 18522 19054 18524
rect 18758 18470 18804 18522
rect 18804 18470 18814 18522
rect 18838 18470 18868 18522
rect 18868 18470 18880 18522
rect 18880 18470 18894 18522
rect 18918 18470 18932 18522
rect 18932 18470 18944 18522
rect 18944 18470 18974 18522
rect 18998 18470 19008 18522
rect 19008 18470 19054 18522
rect 18758 18468 18814 18470
rect 18838 18468 18894 18470
rect 18918 18468 18974 18470
rect 18998 18468 19054 18470
rect 18758 17434 18814 17436
rect 18838 17434 18894 17436
rect 18918 17434 18974 17436
rect 18998 17434 19054 17436
rect 18758 17382 18804 17434
rect 18804 17382 18814 17434
rect 18838 17382 18868 17434
rect 18868 17382 18880 17434
rect 18880 17382 18894 17434
rect 18918 17382 18932 17434
rect 18932 17382 18944 17434
rect 18944 17382 18974 17434
rect 18998 17382 19008 17434
rect 19008 17382 19054 17434
rect 18758 17380 18814 17382
rect 18838 17380 18894 17382
rect 18918 17380 18974 17382
rect 18998 17380 19054 17382
rect 19154 17176 19210 17232
rect 18758 16346 18814 16348
rect 18838 16346 18894 16348
rect 18918 16346 18974 16348
rect 18998 16346 19054 16348
rect 18758 16294 18804 16346
rect 18804 16294 18814 16346
rect 18838 16294 18868 16346
rect 18868 16294 18880 16346
rect 18880 16294 18894 16346
rect 18918 16294 18932 16346
rect 18932 16294 18944 16346
rect 18944 16294 18974 16346
rect 18998 16294 19008 16346
rect 19008 16294 19054 16346
rect 18758 16292 18814 16294
rect 18838 16292 18894 16294
rect 18918 16292 18974 16294
rect 18998 16292 19054 16294
rect 18758 15258 18814 15260
rect 18838 15258 18894 15260
rect 18918 15258 18974 15260
rect 18998 15258 19054 15260
rect 18758 15206 18804 15258
rect 18804 15206 18814 15258
rect 18838 15206 18868 15258
rect 18868 15206 18880 15258
rect 18880 15206 18894 15258
rect 18918 15206 18932 15258
rect 18932 15206 18944 15258
rect 18944 15206 18974 15258
rect 18998 15206 19008 15258
rect 19008 15206 19054 15258
rect 18758 15204 18814 15206
rect 18838 15204 18894 15206
rect 18918 15204 18974 15206
rect 18998 15204 19054 15206
rect 18758 14170 18814 14172
rect 18838 14170 18894 14172
rect 18918 14170 18974 14172
rect 18998 14170 19054 14172
rect 18758 14118 18804 14170
rect 18804 14118 18814 14170
rect 18838 14118 18868 14170
rect 18868 14118 18880 14170
rect 18880 14118 18894 14170
rect 18918 14118 18932 14170
rect 18932 14118 18944 14170
rect 18944 14118 18974 14170
rect 18998 14118 19008 14170
rect 19008 14118 19054 14170
rect 18758 14116 18814 14118
rect 18838 14116 18894 14118
rect 18918 14116 18974 14118
rect 18998 14116 19054 14118
rect 18758 13082 18814 13084
rect 18838 13082 18894 13084
rect 18918 13082 18974 13084
rect 18998 13082 19054 13084
rect 18758 13030 18804 13082
rect 18804 13030 18814 13082
rect 18838 13030 18868 13082
rect 18868 13030 18880 13082
rect 18880 13030 18894 13082
rect 18918 13030 18932 13082
rect 18932 13030 18944 13082
rect 18944 13030 18974 13082
rect 18998 13030 19008 13082
rect 19008 13030 19054 13082
rect 18758 13028 18814 13030
rect 18838 13028 18894 13030
rect 18918 13028 18974 13030
rect 18998 13028 19054 13030
rect 19430 19372 19486 19408
rect 19430 19352 19432 19372
rect 19432 19352 19484 19372
rect 19484 19352 19486 19372
rect 20994 41520 21050 41576
rect 20902 40976 20958 41032
rect 21086 39380 21088 39400
rect 21088 39380 21140 39400
rect 21140 39380 21142 39400
rect 21086 39344 21142 39380
rect 21725 43002 21781 43004
rect 21805 43002 21861 43004
rect 21885 43002 21941 43004
rect 21965 43002 22021 43004
rect 21725 42950 21771 43002
rect 21771 42950 21781 43002
rect 21805 42950 21835 43002
rect 21835 42950 21847 43002
rect 21847 42950 21861 43002
rect 21885 42950 21899 43002
rect 21899 42950 21911 43002
rect 21911 42950 21941 43002
rect 21965 42950 21975 43002
rect 21975 42950 22021 43002
rect 21725 42948 21781 42950
rect 21805 42948 21861 42950
rect 21885 42948 21941 42950
rect 21965 42948 22021 42950
rect 21725 41914 21781 41916
rect 21805 41914 21861 41916
rect 21885 41914 21941 41916
rect 21965 41914 22021 41916
rect 21725 41862 21771 41914
rect 21771 41862 21781 41914
rect 21805 41862 21835 41914
rect 21835 41862 21847 41914
rect 21847 41862 21861 41914
rect 21885 41862 21899 41914
rect 21899 41862 21911 41914
rect 21911 41862 21941 41914
rect 21965 41862 21975 41914
rect 21975 41862 22021 41914
rect 21725 41860 21781 41862
rect 21805 41860 21861 41862
rect 21885 41860 21941 41862
rect 21965 41860 22021 41862
rect 21454 40976 21510 41032
rect 21362 39208 21418 39264
rect 20994 35672 21050 35728
rect 20718 34584 20774 34640
rect 20074 29008 20130 29064
rect 20074 26968 20130 27024
rect 19338 16496 19394 16552
rect 17682 3848 17738 3904
rect 17958 3848 18014 3904
rect 17590 3052 17646 3088
rect 17590 3032 17592 3052
rect 17592 3032 17644 3052
rect 17644 3032 17646 3052
rect 17682 2388 17684 2408
rect 17684 2388 17736 2408
rect 17736 2388 17738 2408
rect 17682 2352 17738 2388
rect 19154 12280 19210 12336
rect 18758 11994 18814 11996
rect 18838 11994 18894 11996
rect 18918 11994 18974 11996
rect 18998 11994 19054 11996
rect 18758 11942 18804 11994
rect 18804 11942 18814 11994
rect 18838 11942 18868 11994
rect 18868 11942 18880 11994
rect 18880 11942 18894 11994
rect 18918 11942 18932 11994
rect 18932 11942 18944 11994
rect 18944 11942 18974 11994
rect 18998 11942 19008 11994
rect 19008 11942 19054 11994
rect 18758 11940 18814 11942
rect 18838 11940 18894 11942
rect 18918 11940 18974 11942
rect 18998 11940 19054 11942
rect 18758 10906 18814 10908
rect 18838 10906 18894 10908
rect 18918 10906 18974 10908
rect 18998 10906 19054 10908
rect 18758 10854 18804 10906
rect 18804 10854 18814 10906
rect 18838 10854 18868 10906
rect 18868 10854 18880 10906
rect 18880 10854 18894 10906
rect 18918 10854 18932 10906
rect 18932 10854 18944 10906
rect 18944 10854 18974 10906
rect 18998 10854 19008 10906
rect 19008 10854 19054 10906
rect 18758 10852 18814 10854
rect 18838 10852 18894 10854
rect 18918 10852 18974 10854
rect 18998 10852 19054 10854
rect 18758 9818 18814 9820
rect 18838 9818 18894 9820
rect 18918 9818 18974 9820
rect 18998 9818 19054 9820
rect 18758 9766 18804 9818
rect 18804 9766 18814 9818
rect 18838 9766 18868 9818
rect 18868 9766 18880 9818
rect 18880 9766 18894 9818
rect 18918 9766 18932 9818
rect 18932 9766 18944 9818
rect 18944 9766 18974 9818
rect 18998 9766 19008 9818
rect 19008 9766 19054 9818
rect 18758 9764 18814 9766
rect 18838 9764 18894 9766
rect 18918 9764 18974 9766
rect 18998 9764 19054 9766
rect 18758 8730 18814 8732
rect 18838 8730 18894 8732
rect 18918 8730 18974 8732
rect 18998 8730 19054 8732
rect 18758 8678 18804 8730
rect 18804 8678 18814 8730
rect 18838 8678 18868 8730
rect 18868 8678 18880 8730
rect 18880 8678 18894 8730
rect 18918 8678 18932 8730
rect 18932 8678 18944 8730
rect 18944 8678 18974 8730
rect 18998 8678 19008 8730
rect 19008 8678 19054 8730
rect 18758 8676 18814 8678
rect 18838 8676 18894 8678
rect 18918 8676 18974 8678
rect 18998 8676 19054 8678
rect 18758 7642 18814 7644
rect 18838 7642 18894 7644
rect 18918 7642 18974 7644
rect 18998 7642 19054 7644
rect 18758 7590 18804 7642
rect 18804 7590 18814 7642
rect 18838 7590 18868 7642
rect 18868 7590 18880 7642
rect 18880 7590 18894 7642
rect 18918 7590 18932 7642
rect 18932 7590 18944 7642
rect 18944 7590 18974 7642
rect 18998 7590 19008 7642
rect 19008 7590 19054 7642
rect 18758 7588 18814 7590
rect 18838 7588 18894 7590
rect 18918 7588 18974 7590
rect 18998 7588 19054 7590
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 19982 21120 20038 21176
rect 20718 28464 20774 28520
rect 20626 25236 20628 25256
rect 20628 25236 20680 25256
rect 20680 25236 20682 25256
rect 20626 25200 20682 25236
rect 20258 21256 20314 21312
rect 20074 15952 20130 16008
rect 19798 13504 19854 13560
rect 19706 11600 19762 11656
rect 19982 13232 20038 13288
rect 20994 22072 21050 22128
rect 20810 20984 20866 21040
rect 21270 34992 21326 35048
rect 21270 26968 21326 27024
rect 21822 41384 21878 41440
rect 22558 41520 22614 41576
rect 22926 43152 22982 43208
rect 21822 41132 21878 41168
rect 21822 41112 21824 41132
rect 21824 41112 21876 41132
rect 21876 41112 21878 41132
rect 22190 40976 22246 41032
rect 21725 40826 21781 40828
rect 21805 40826 21861 40828
rect 21885 40826 21941 40828
rect 21965 40826 22021 40828
rect 21725 40774 21771 40826
rect 21771 40774 21781 40826
rect 21805 40774 21835 40826
rect 21835 40774 21847 40826
rect 21847 40774 21861 40826
rect 21885 40774 21899 40826
rect 21899 40774 21911 40826
rect 21911 40774 21941 40826
rect 21965 40774 21975 40826
rect 21975 40774 22021 40826
rect 21725 40772 21781 40774
rect 21805 40772 21861 40774
rect 21885 40772 21941 40774
rect 21965 40772 22021 40774
rect 22098 40704 22154 40760
rect 21638 40432 21694 40488
rect 22098 40468 22100 40488
rect 22100 40468 22152 40488
rect 22152 40468 22154 40488
rect 22098 40432 22154 40468
rect 21822 40180 21878 40216
rect 21822 40160 21824 40180
rect 21824 40160 21876 40180
rect 21876 40160 21878 40180
rect 21914 40024 21970 40080
rect 21725 39738 21781 39740
rect 21805 39738 21861 39740
rect 21885 39738 21941 39740
rect 21965 39738 22021 39740
rect 21725 39686 21771 39738
rect 21771 39686 21781 39738
rect 21805 39686 21835 39738
rect 21835 39686 21847 39738
rect 21847 39686 21861 39738
rect 21885 39686 21899 39738
rect 21899 39686 21911 39738
rect 21911 39686 21941 39738
rect 21965 39686 21975 39738
rect 21975 39686 22021 39738
rect 21725 39684 21781 39686
rect 21805 39684 21861 39686
rect 21885 39684 21941 39686
rect 21965 39684 22021 39686
rect 22466 40976 22522 41032
rect 22466 40724 22522 40760
rect 22466 40704 22468 40724
rect 22468 40704 22520 40724
rect 22520 40704 22522 40724
rect 22650 40568 22706 40624
rect 22650 40060 22652 40080
rect 22652 40060 22704 40080
rect 22704 40060 22706 40080
rect 22650 40024 22706 40060
rect 21725 38650 21781 38652
rect 21805 38650 21861 38652
rect 21885 38650 21941 38652
rect 21965 38650 22021 38652
rect 21725 38598 21771 38650
rect 21771 38598 21781 38650
rect 21805 38598 21835 38650
rect 21835 38598 21847 38650
rect 21847 38598 21861 38650
rect 21885 38598 21899 38650
rect 21899 38598 21911 38650
rect 21911 38598 21941 38650
rect 21965 38598 21975 38650
rect 21975 38598 22021 38650
rect 21725 38596 21781 38598
rect 21805 38596 21861 38598
rect 21885 38596 21941 38598
rect 21965 38596 22021 38598
rect 21725 37562 21781 37564
rect 21805 37562 21861 37564
rect 21885 37562 21941 37564
rect 21965 37562 22021 37564
rect 21725 37510 21771 37562
rect 21771 37510 21781 37562
rect 21805 37510 21835 37562
rect 21835 37510 21847 37562
rect 21847 37510 21861 37562
rect 21885 37510 21899 37562
rect 21899 37510 21911 37562
rect 21911 37510 21941 37562
rect 21965 37510 21975 37562
rect 21975 37510 22021 37562
rect 21725 37508 21781 37510
rect 21805 37508 21861 37510
rect 21885 37508 21941 37510
rect 21965 37508 22021 37510
rect 21725 36474 21781 36476
rect 21805 36474 21861 36476
rect 21885 36474 21941 36476
rect 21965 36474 22021 36476
rect 21725 36422 21771 36474
rect 21771 36422 21781 36474
rect 21805 36422 21835 36474
rect 21835 36422 21847 36474
rect 21847 36422 21861 36474
rect 21885 36422 21899 36474
rect 21899 36422 21911 36474
rect 21911 36422 21941 36474
rect 21965 36422 21975 36474
rect 21975 36422 22021 36474
rect 21725 36420 21781 36422
rect 21805 36420 21861 36422
rect 21885 36420 21941 36422
rect 21965 36420 22021 36422
rect 21725 35386 21781 35388
rect 21805 35386 21861 35388
rect 21885 35386 21941 35388
rect 21965 35386 22021 35388
rect 21725 35334 21771 35386
rect 21771 35334 21781 35386
rect 21805 35334 21835 35386
rect 21835 35334 21847 35386
rect 21847 35334 21861 35386
rect 21885 35334 21899 35386
rect 21899 35334 21911 35386
rect 21911 35334 21941 35386
rect 21965 35334 21975 35386
rect 21975 35334 22021 35386
rect 21725 35332 21781 35334
rect 21805 35332 21861 35334
rect 21885 35332 21941 35334
rect 21965 35332 22021 35334
rect 21725 34298 21781 34300
rect 21805 34298 21861 34300
rect 21885 34298 21941 34300
rect 21965 34298 22021 34300
rect 21725 34246 21771 34298
rect 21771 34246 21781 34298
rect 21805 34246 21835 34298
rect 21835 34246 21847 34298
rect 21847 34246 21861 34298
rect 21885 34246 21899 34298
rect 21899 34246 21911 34298
rect 21911 34246 21941 34298
rect 21965 34246 21975 34298
rect 21975 34246 22021 34298
rect 21725 34244 21781 34246
rect 21805 34244 21861 34246
rect 21885 34244 21941 34246
rect 21965 34244 22021 34246
rect 21725 33210 21781 33212
rect 21805 33210 21861 33212
rect 21885 33210 21941 33212
rect 21965 33210 22021 33212
rect 21725 33158 21771 33210
rect 21771 33158 21781 33210
rect 21805 33158 21835 33210
rect 21835 33158 21847 33210
rect 21847 33158 21861 33210
rect 21885 33158 21899 33210
rect 21899 33158 21911 33210
rect 21911 33158 21941 33210
rect 21965 33158 21975 33210
rect 21975 33158 22021 33210
rect 21725 33156 21781 33158
rect 21805 33156 21861 33158
rect 21885 33156 21941 33158
rect 21965 33156 22021 33158
rect 21725 32122 21781 32124
rect 21805 32122 21861 32124
rect 21885 32122 21941 32124
rect 21965 32122 22021 32124
rect 21725 32070 21771 32122
rect 21771 32070 21781 32122
rect 21805 32070 21835 32122
rect 21835 32070 21847 32122
rect 21847 32070 21861 32122
rect 21885 32070 21899 32122
rect 21899 32070 21911 32122
rect 21911 32070 21941 32122
rect 21965 32070 21975 32122
rect 21975 32070 22021 32122
rect 21725 32068 21781 32070
rect 21805 32068 21861 32070
rect 21885 32068 21941 32070
rect 21965 32068 22021 32070
rect 21725 31034 21781 31036
rect 21805 31034 21861 31036
rect 21885 31034 21941 31036
rect 21965 31034 22021 31036
rect 21725 30982 21771 31034
rect 21771 30982 21781 31034
rect 21805 30982 21835 31034
rect 21835 30982 21847 31034
rect 21847 30982 21861 31034
rect 21885 30982 21899 31034
rect 21899 30982 21911 31034
rect 21911 30982 21941 31034
rect 21965 30982 21975 31034
rect 21975 30982 22021 31034
rect 21725 30980 21781 30982
rect 21805 30980 21861 30982
rect 21885 30980 21941 30982
rect 21965 30980 22021 30982
rect 21725 29946 21781 29948
rect 21805 29946 21861 29948
rect 21885 29946 21941 29948
rect 21965 29946 22021 29948
rect 21725 29894 21771 29946
rect 21771 29894 21781 29946
rect 21805 29894 21835 29946
rect 21835 29894 21847 29946
rect 21847 29894 21861 29946
rect 21885 29894 21899 29946
rect 21899 29894 21911 29946
rect 21911 29894 21941 29946
rect 21965 29894 21975 29946
rect 21975 29894 22021 29946
rect 21725 29892 21781 29894
rect 21805 29892 21861 29894
rect 21885 29892 21941 29894
rect 21965 29892 22021 29894
rect 22098 29688 22154 29744
rect 21725 28858 21781 28860
rect 21805 28858 21861 28860
rect 21885 28858 21941 28860
rect 21965 28858 22021 28860
rect 21725 28806 21771 28858
rect 21771 28806 21781 28858
rect 21805 28806 21835 28858
rect 21835 28806 21847 28858
rect 21847 28806 21861 28858
rect 21885 28806 21899 28858
rect 21899 28806 21911 28858
rect 21911 28806 21941 28858
rect 21965 28806 21975 28858
rect 21975 28806 22021 28858
rect 21725 28804 21781 28806
rect 21805 28804 21861 28806
rect 21885 28804 21941 28806
rect 21965 28804 22021 28806
rect 21725 27770 21781 27772
rect 21805 27770 21861 27772
rect 21885 27770 21941 27772
rect 21965 27770 22021 27772
rect 21725 27718 21771 27770
rect 21771 27718 21781 27770
rect 21805 27718 21835 27770
rect 21835 27718 21847 27770
rect 21847 27718 21861 27770
rect 21885 27718 21899 27770
rect 21899 27718 21911 27770
rect 21911 27718 21941 27770
rect 21965 27718 21975 27770
rect 21975 27718 22021 27770
rect 21725 27716 21781 27718
rect 21805 27716 21861 27718
rect 21885 27716 21941 27718
rect 21965 27716 22021 27718
rect 22926 41248 22982 41304
rect 23202 43288 23258 43344
rect 23202 41384 23258 41440
rect 23110 40024 23166 40080
rect 23110 39244 23112 39264
rect 23112 39244 23164 39264
rect 23164 39244 23166 39264
rect 23110 39208 23166 39244
rect 23018 39072 23074 39128
rect 23478 40432 23534 40488
rect 23386 39480 23442 39536
rect 23662 40876 23664 40896
rect 23664 40876 23716 40896
rect 23716 40876 23718 40896
rect 23662 40840 23718 40876
rect 23662 40296 23718 40352
rect 24692 43546 24748 43548
rect 24772 43546 24828 43548
rect 24852 43546 24908 43548
rect 24932 43546 24988 43548
rect 24692 43494 24738 43546
rect 24738 43494 24748 43546
rect 24772 43494 24802 43546
rect 24802 43494 24814 43546
rect 24814 43494 24828 43546
rect 24852 43494 24866 43546
rect 24866 43494 24878 43546
rect 24878 43494 24908 43546
rect 24932 43494 24942 43546
rect 24942 43494 24988 43546
rect 24692 43492 24748 43494
rect 24772 43492 24828 43494
rect 24852 43492 24908 43494
rect 24932 43492 24988 43494
rect 24692 42458 24748 42460
rect 24772 42458 24828 42460
rect 24852 42458 24908 42460
rect 24932 42458 24988 42460
rect 24692 42406 24738 42458
rect 24738 42406 24748 42458
rect 24772 42406 24802 42458
rect 24802 42406 24814 42458
rect 24814 42406 24828 42458
rect 24852 42406 24866 42458
rect 24866 42406 24878 42458
rect 24878 42406 24908 42458
rect 24932 42406 24942 42458
rect 24942 42406 24988 42458
rect 24692 42404 24748 42406
rect 24772 42404 24828 42406
rect 24852 42404 24908 42406
rect 24932 42404 24988 42406
rect 24122 41928 24178 41984
rect 23938 40160 23994 40216
rect 22742 35944 22798 36000
rect 24122 39344 24178 39400
rect 24398 39788 24400 39808
rect 24400 39788 24452 39808
rect 24452 39788 24454 39808
rect 24398 39752 24454 39788
rect 24398 38700 24400 38720
rect 24400 38700 24452 38720
rect 24452 38700 24454 38720
rect 24398 38664 24454 38700
rect 24398 37612 24400 37632
rect 24400 37612 24452 37632
rect 24452 37612 24454 37632
rect 24398 37576 24454 37612
rect 24122 37168 24178 37224
rect 22742 33496 22798 33552
rect 22558 33224 22614 33280
rect 21725 26682 21781 26684
rect 21805 26682 21861 26684
rect 21885 26682 21941 26684
rect 21965 26682 22021 26684
rect 21725 26630 21771 26682
rect 21771 26630 21781 26682
rect 21805 26630 21835 26682
rect 21835 26630 21847 26682
rect 21847 26630 21861 26682
rect 21885 26630 21899 26682
rect 21899 26630 21911 26682
rect 21911 26630 21941 26682
rect 21965 26630 21975 26682
rect 21975 26630 22021 26682
rect 21725 26628 21781 26630
rect 21805 26628 21861 26630
rect 21885 26628 21941 26630
rect 21965 26628 22021 26630
rect 21638 26152 21694 26208
rect 21725 25594 21781 25596
rect 21805 25594 21861 25596
rect 21885 25594 21941 25596
rect 21965 25594 22021 25596
rect 21725 25542 21771 25594
rect 21771 25542 21781 25594
rect 21805 25542 21835 25594
rect 21835 25542 21847 25594
rect 21847 25542 21861 25594
rect 21885 25542 21899 25594
rect 21899 25542 21911 25594
rect 21911 25542 21941 25594
rect 21965 25542 21975 25594
rect 21975 25542 22021 25594
rect 21725 25540 21781 25542
rect 21805 25540 21861 25542
rect 21885 25540 21941 25542
rect 21965 25540 22021 25542
rect 22098 24792 22154 24848
rect 21362 22072 21418 22128
rect 21086 19352 21142 19408
rect 19890 8336 19946 8392
rect 20534 13268 20536 13288
rect 20536 13268 20588 13288
rect 20588 13268 20590 13288
rect 20534 13232 20590 13268
rect 20902 16632 20958 16688
rect 20902 13640 20958 13696
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 18694 5208 18750 5264
rect 19430 6432 19486 6488
rect 19430 6160 19486 6216
rect 19338 4800 19394 4856
rect 18510 3848 18566 3904
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 19062 1300 19064 1320
rect 19064 1300 19116 1320
rect 19116 1300 19118 1320
rect 19062 1264 19118 1300
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 19890 4664 19946 4720
rect 20442 7520 20498 7576
rect 20626 7384 20682 7440
rect 20258 6160 20314 6216
rect 20350 5480 20406 5536
rect 19982 3032 20038 3088
rect 20718 6568 20774 6624
rect 20626 6024 20682 6080
rect 21725 24506 21781 24508
rect 21805 24506 21861 24508
rect 21885 24506 21941 24508
rect 21965 24506 22021 24508
rect 21725 24454 21771 24506
rect 21771 24454 21781 24506
rect 21805 24454 21835 24506
rect 21835 24454 21847 24506
rect 21847 24454 21861 24506
rect 21885 24454 21899 24506
rect 21899 24454 21911 24506
rect 21911 24454 21941 24506
rect 21965 24454 21975 24506
rect 21975 24454 22021 24506
rect 21725 24452 21781 24454
rect 21805 24452 21861 24454
rect 21885 24452 21941 24454
rect 21965 24452 22021 24454
rect 21638 23724 21694 23760
rect 21638 23704 21640 23724
rect 21640 23704 21692 23724
rect 21692 23704 21694 23724
rect 21725 23418 21781 23420
rect 21805 23418 21861 23420
rect 21885 23418 21941 23420
rect 21965 23418 22021 23420
rect 21725 23366 21771 23418
rect 21771 23366 21781 23418
rect 21805 23366 21835 23418
rect 21835 23366 21847 23418
rect 21847 23366 21861 23418
rect 21885 23366 21899 23418
rect 21899 23366 21911 23418
rect 21911 23366 21941 23418
rect 21965 23366 21975 23418
rect 21975 23366 22021 23418
rect 21725 23364 21781 23366
rect 21805 23364 21861 23366
rect 21885 23364 21941 23366
rect 21965 23364 22021 23366
rect 22190 23432 22246 23488
rect 21638 22480 21694 22536
rect 21725 22330 21781 22332
rect 21805 22330 21861 22332
rect 21885 22330 21941 22332
rect 21965 22330 22021 22332
rect 21725 22278 21771 22330
rect 21771 22278 21781 22330
rect 21805 22278 21835 22330
rect 21835 22278 21847 22330
rect 21847 22278 21861 22330
rect 21885 22278 21899 22330
rect 21899 22278 21911 22330
rect 21911 22278 21941 22330
rect 21965 22278 21975 22330
rect 21975 22278 22021 22330
rect 21725 22276 21781 22278
rect 21805 22276 21861 22278
rect 21885 22276 21941 22278
rect 21965 22276 22021 22278
rect 21725 21242 21781 21244
rect 21805 21242 21861 21244
rect 21885 21242 21941 21244
rect 21965 21242 22021 21244
rect 21725 21190 21771 21242
rect 21771 21190 21781 21242
rect 21805 21190 21835 21242
rect 21835 21190 21847 21242
rect 21847 21190 21861 21242
rect 21885 21190 21899 21242
rect 21899 21190 21911 21242
rect 21911 21190 21941 21242
rect 21965 21190 21975 21242
rect 21975 21190 22021 21242
rect 21725 21188 21781 21190
rect 21805 21188 21861 21190
rect 21885 21188 21941 21190
rect 21965 21188 22021 21190
rect 22466 22480 22522 22536
rect 21725 20154 21781 20156
rect 21805 20154 21861 20156
rect 21885 20154 21941 20156
rect 21965 20154 22021 20156
rect 21725 20102 21771 20154
rect 21771 20102 21781 20154
rect 21805 20102 21835 20154
rect 21835 20102 21847 20154
rect 21847 20102 21861 20154
rect 21885 20102 21899 20154
rect 21899 20102 21911 20154
rect 21911 20102 21941 20154
rect 21965 20102 21975 20154
rect 21975 20102 22021 20154
rect 21725 20100 21781 20102
rect 21805 20100 21861 20102
rect 21885 20100 21941 20102
rect 21965 20100 22021 20102
rect 21725 19066 21781 19068
rect 21805 19066 21861 19068
rect 21885 19066 21941 19068
rect 21965 19066 22021 19068
rect 21725 19014 21771 19066
rect 21771 19014 21781 19066
rect 21805 19014 21835 19066
rect 21835 19014 21847 19066
rect 21847 19014 21861 19066
rect 21885 19014 21899 19066
rect 21899 19014 21911 19066
rect 21911 19014 21941 19066
rect 21965 19014 21975 19066
rect 21975 19014 22021 19066
rect 21725 19012 21781 19014
rect 21805 19012 21861 19014
rect 21885 19012 21941 19014
rect 21965 19012 22021 19014
rect 21725 17978 21781 17980
rect 21805 17978 21861 17980
rect 21885 17978 21941 17980
rect 21965 17978 22021 17980
rect 21725 17926 21771 17978
rect 21771 17926 21781 17978
rect 21805 17926 21835 17978
rect 21835 17926 21847 17978
rect 21847 17926 21861 17978
rect 21885 17926 21899 17978
rect 21899 17926 21911 17978
rect 21911 17926 21941 17978
rect 21965 17926 21975 17978
rect 21975 17926 22021 17978
rect 21725 17924 21781 17926
rect 21805 17924 21861 17926
rect 21885 17924 21941 17926
rect 21965 17924 22021 17926
rect 21638 17720 21694 17776
rect 21725 16890 21781 16892
rect 21805 16890 21861 16892
rect 21885 16890 21941 16892
rect 21965 16890 22021 16892
rect 21725 16838 21771 16890
rect 21771 16838 21781 16890
rect 21805 16838 21835 16890
rect 21835 16838 21847 16890
rect 21847 16838 21861 16890
rect 21885 16838 21899 16890
rect 21899 16838 21911 16890
rect 21911 16838 21941 16890
rect 21965 16838 21975 16890
rect 21975 16838 22021 16890
rect 21725 16836 21781 16838
rect 21805 16836 21861 16838
rect 21885 16836 21941 16838
rect 21965 16836 22021 16838
rect 22190 16088 22246 16144
rect 21725 15802 21781 15804
rect 21805 15802 21861 15804
rect 21885 15802 21941 15804
rect 21965 15802 22021 15804
rect 21725 15750 21771 15802
rect 21771 15750 21781 15802
rect 21805 15750 21835 15802
rect 21835 15750 21847 15802
rect 21847 15750 21861 15802
rect 21885 15750 21899 15802
rect 21899 15750 21911 15802
rect 21911 15750 21941 15802
rect 21965 15750 21975 15802
rect 21975 15750 22021 15802
rect 21725 15748 21781 15750
rect 21805 15748 21861 15750
rect 21885 15748 21941 15750
rect 21965 15748 22021 15750
rect 21725 14714 21781 14716
rect 21805 14714 21861 14716
rect 21885 14714 21941 14716
rect 21965 14714 22021 14716
rect 21725 14662 21771 14714
rect 21771 14662 21781 14714
rect 21805 14662 21835 14714
rect 21835 14662 21847 14714
rect 21847 14662 21861 14714
rect 21885 14662 21899 14714
rect 21899 14662 21911 14714
rect 21911 14662 21941 14714
rect 21965 14662 21975 14714
rect 21975 14662 22021 14714
rect 21725 14660 21781 14662
rect 21805 14660 21861 14662
rect 21885 14660 21941 14662
rect 21965 14660 22021 14662
rect 21270 6840 21326 6896
rect 20534 5344 20590 5400
rect 20718 5072 20774 5128
rect 21178 5788 21180 5808
rect 21180 5788 21232 5808
rect 21232 5788 21234 5808
rect 21178 5752 21234 5788
rect 20718 3304 20774 3360
rect 21270 4528 21326 4584
rect 21086 4004 21142 4040
rect 21086 3984 21088 4004
rect 21088 3984 21140 4004
rect 21140 3984 21142 4004
rect 20718 2896 20774 2952
rect 20534 2624 20590 2680
rect 21178 3440 21234 3496
rect 20718 1808 20774 1864
rect 20718 584 20774 640
rect 21546 7792 21602 7848
rect 21546 6060 21548 6080
rect 21548 6060 21600 6080
rect 21600 6060 21602 6080
rect 21546 6024 21602 6060
rect 22098 13912 22154 13968
rect 22098 13676 22100 13696
rect 22100 13676 22152 13696
rect 22152 13676 22154 13696
rect 22098 13640 22154 13676
rect 21725 13626 21781 13628
rect 21805 13626 21861 13628
rect 21885 13626 21941 13628
rect 21965 13626 22021 13628
rect 21725 13574 21771 13626
rect 21771 13574 21781 13626
rect 21805 13574 21835 13626
rect 21835 13574 21847 13626
rect 21847 13574 21861 13626
rect 21885 13574 21899 13626
rect 21899 13574 21911 13626
rect 21911 13574 21941 13626
rect 21965 13574 21975 13626
rect 21975 13574 22021 13626
rect 21725 13572 21781 13574
rect 21805 13572 21861 13574
rect 21885 13572 21941 13574
rect 21965 13572 22021 13574
rect 21725 12538 21781 12540
rect 21805 12538 21861 12540
rect 21885 12538 21941 12540
rect 21965 12538 22021 12540
rect 21725 12486 21771 12538
rect 21771 12486 21781 12538
rect 21805 12486 21835 12538
rect 21835 12486 21847 12538
rect 21847 12486 21861 12538
rect 21885 12486 21899 12538
rect 21899 12486 21911 12538
rect 21911 12486 21941 12538
rect 21965 12486 21975 12538
rect 21975 12486 22021 12538
rect 21725 12484 21781 12486
rect 21805 12484 21861 12486
rect 21885 12484 21941 12486
rect 21965 12484 22021 12486
rect 21725 11450 21781 11452
rect 21805 11450 21861 11452
rect 21885 11450 21941 11452
rect 21965 11450 22021 11452
rect 21725 11398 21771 11450
rect 21771 11398 21781 11450
rect 21805 11398 21835 11450
rect 21835 11398 21847 11450
rect 21847 11398 21861 11450
rect 21885 11398 21899 11450
rect 21899 11398 21911 11450
rect 21911 11398 21941 11450
rect 21965 11398 21975 11450
rect 21975 11398 22021 11450
rect 21725 11396 21781 11398
rect 21805 11396 21861 11398
rect 21885 11396 21941 11398
rect 21965 11396 22021 11398
rect 21725 10362 21781 10364
rect 21805 10362 21861 10364
rect 21885 10362 21941 10364
rect 21965 10362 22021 10364
rect 21725 10310 21771 10362
rect 21771 10310 21781 10362
rect 21805 10310 21835 10362
rect 21835 10310 21847 10362
rect 21847 10310 21861 10362
rect 21885 10310 21899 10362
rect 21899 10310 21911 10362
rect 21911 10310 21941 10362
rect 21965 10310 21975 10362
rect 21975 10310 22021 10362
rect 21725 10308 21781 10310
rect 21805 10308 21861 10310
rect 21885 10308 21941 10310
rect 21965 10308 22021 10310
rect 23202 31764 23204 31784
rect 23204 31764 23256 31784
rect 23256 31764 23258 31784
rect 23202 31728 23258 31764
rect 24398 36524 24400 36544
rect 24400 36524 24452 36544
rect 24452 36524 24454 36544
rect 24398 36488 24454 36524
rect 24398 35436 24400 35456
rect 24400 35436 24452 35456
rect 24452 35436 24454 35456
rect 24398 35400 24454 35436
rect 24398 34484 24400 34504
rect 24400 34484 24452 34504
rect 24452 34484 24454 34504
rect 24398 34448 24454 34484
rect 24398 33260 24400 33280
rect 24400 33260 24452 33280
rect 24452 33260 24454 33280
rect 24398 33224 24454 33260
rect 24398 32172 24400 32192
rect 24400 32172 24452 32192
rect 24452 32172 24454 32192
rect 24398 32136 24454 32172
rect 23202 28600 23258 28656
rect 22926 24792 22982 24848
rect 24398 31084 24400 31104
rect 24400 31084 24452 31104
rect 24452 31084 24454 31104
rect 24398 31048 24454 31084
rect 24398 29996 24400 30016
rect 24400 29996 24452 30016
rect 24452 29996 24454 30016
rect 24398 29960 24454 29996
rect 24214 26152 24270 26208
rect 23846 24248 23902 24304
rect 22558 13524 22614 13560
rect 22558 13504 22560 13524
rect 22560 13504 22612 13524
rect 22612 13504 22614 13524
rect 21725 9274 21781 9276
rect 21805 9274 21861 9276
rect 21885 9274 21941 9276
rect 21965 9274 22021 9276
rect 21725 9222 21771 9274
rect 21771 9222 21781 9274
rect 21805 9222 21835 9274
rect 21835 9222 21847 9274
rect 21847 9222 21861 9274
rect 21885 9222 21899 9274
rect 21899 9222 21911 9274
rect 21911 9222 21941 9274
rect 21965 9222 21975 9274
rect 21975 9222 22021 9274
rect 21725 9220 21781 9222
rect 21805 9220 21861 9222
rect 21885 9220 21941 9222
rect 21965 9220 22021 9222
rect 21725 8186 21781 8188
rect 21805 8186 21861 8188
rect 21885 8186 21941 8188
rect 21965 8186 22021 8188
rect 21725 8134 21771 8186
rect 21771 8134 21781 8186
rect 21805 8134 21835 8186
rect 21835 8134 21847 8186
rect 21847 8134 21861 8186
rect 21885 8134 21899 8186
rect 21899 8134 21911 8186
rect 21911 8134 21941 8186
rect 21965 8134 21975 8186
rect 21975 8134 22021 8186
rect 21725 8132 21781 8134
rect 21805 8132 21861 8134
rect 21885 8132 21941 8134
rect 21965 8132 22021 8134
rect 21725 7098 21781 7100
rect 21805 7098 21861 7100
rect 21885 7098 21941 7100
rect 21965 7098 22021 7100
rect 21725 7046 21771 7098
rect 21771 7046 21781 7098
rect 21805 7046 21835 7098
rect 21835 7046 21847 7098
rect 21847 7046 21861 7098
rect 21885 7046 21899 7098
rect 21899 7046 21911 7098
rect 21911 7046 21941 7098
rect 21965 7046 21975 7098
rect 21975 7046 22021 7098
rect 21725 7044 21781 7046
rect 21805 7044 21861 7046
rect 21885 7044 21941 7046
rect 21965 7044 22021 7046
rect 21730 6840 21786 6896
rect 21730 6296 21786 6352
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 21454 4800 21510 4856
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 22006 4664 22062 4720
rect 21638 3984 21694 4040
rect 21822 3984 21878 4040
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 21914 2488 21970 2544
rect 22098 2216 22154 2272
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 21638 1300 21640 1320
rect 21640 1300 21692 1320
rect 21692 1300 21694 1320
rect 21638 1264 21694 1300
rect 21362 1128 21418 1184
rect 23846 21292 23848 21312
rect 23848 21292 23900 21312
rect 23900 21292 23902 21312
rect 23846 21256 23902 21292
rect 23846 19116 23848 19136
rect 23848 19116 23900 19136
rect 23900 19116 23902 19136
rect 23846 19080 23902 19116
rect 22926 13912 22982 13968
rect 23294 13676 23296 13696
rect 23296 13676 23348 13696
rect 23348 13676 23350 13696
rect 23294 13640 23350 13676
rect 23202 13504 23258 13560
rect 24030 20168 24086 20224
rect 24398 28872 24454 28928
rect 24398 27820 24400 27840
rect 24400 27820 24452 27840
rect 24452 27820 24454 27840
rect 24398 27784 24454 27820
rect 24398 26732 24400 26752
rect 24400 26732 24452 26752
rect 24452 26732 24454 26752
rect 24398 26696 24454 26732
rect 24398 25644 24400 25664
rect 24400 25644 24452 25664
rect 24452 25644 24454 25664
rect 24398 25608 24454 25644
rect 24398 24556 24400 24576
rect 24400 24556 24452 24576
rect 24452 24556 24454 24576
rect 24398 24520 24454 24556
rect 24398 23468 24400 23488
rect 24400 23468 24452 23488
rect 24452 23468 24454 23488
rect 24398 23432 24454 23468
rect 24692 41370 24748 41372
rect 24772 41370 24828 41372
rect 24852 41370 24908 41372
rect 24932 41370 24988 41372
rect 24692 41318 24738 41370
rect 24738 41318 24748 41370
rect 24772 41318 24802 41370
rect 24802 41318 24814 41370
rect 24814 41318 24828 41370
rect 24852 41318 24866 41370
rect 24866 41318 24878 41370
rect 24878 41318 24908 41370
rect 24932 41318 24942 41370
rect 24942 41318 24988 41370
rect 24692 41316 24748 41318
rect 24772 41316 24828 41318
rect 24852 41316 24908 41318
rect 24932 41316 24988 41318
rect 25134 42472 25190 42528
rect 25318 43016 25374 43072
rect 25134 41384 25190 41440
rect 25134 40296 25190 40352
rect 24692 40282 24748 40284
rect 24772 40282 24828 40284
rect 24852 40282 24908 40284
rect 24932 40282 24988 40284
rect 24692 40230 24738 40282
rect 24738 40230 24748 40282
rect 24772 40230 24802 40282
rect 24802 40230 24814 40282
rect 24814 40230 24828 40282
rect 24852 40230 24866 40282
rect 24866 40230 24878 40282
rect 24878 40230 24908 40282
rect 24932 40230 24942 40282
rect 24942 40230 24988 40282
rect 24692 40228 24748 40230
rect 24772 40228 24828 40230
rect 24852 40228 24908 40230
rect 24932 40228 24988 40230
rect 25226 39244 25228 39264
rect 25228 39244 25280 39264
rect 25280 39244 25282 39264
rect 25226 39208 25282 39244
rect 24692 39194 24748 39196
rect 24772 39194 24828 39196
rect 24852 39194 24908 39196
rect 24932 39194 24988 39196
rect 24692 39142 24738 39194
rect 24738 39142 24748 39194
rect 24772 39142 24802 39194
rect 24802 39142 24814 39194
rect 24814 39142 24828 39194
rect 24852 39142 24866 39194
rect 24866 39142 24878 39194
rect 24878 39142 24908 39194
rect 24932 39142 24942 39194
rect 24942 39142 24988 39194
rect 24692 39140 24748 39142
rect 24772 39140 24828 39142
rect 24852 39140 24908 39142
rect 24932 39140 24988 39142
rect 25226 38156 25228 38176
rect 25228 38156 25280 38176
rect 25280 38156 25282 38176
rect 25226 38120 25282 38156
rect 24692 38106 24748 38108
rect 24772 38106 24828 38108
rect 24852 38106 24908 38108
rect 24932 38106 24988 38108
rect 24692 38054 24738 38106
rect 24738 38054 24748 38106
rect 24772 38054 24802 38106
rect 24802 38054 24814 38106
rect 24814 38054 24828 38106
rect 24852 38054 24866 38106
rect 24866 38054 24878 38106
rect 24878 38054 24908 38106
rect 24932 38054 24942 38106
rect 24942 38054 24988 38106
rect 24692 38052 24748 38054
rect 24772 38052 24828 38054
rect 24852 38052 24908 38054
rect 24932 38052 24988 38054
rect 24692 37018 24748 37020
rect 24772 37018 24828 37020
rect 24852 37018 24908 37020
rect 24932 37018 24988 37020
rect 24692 36966 24738 37018
rect 24738 36966 24748 37018
rect 24772 36966 24802 37018
rect 24802 36966 24814 37018
rect 24814 36966 24828 37018
rect 24852 36966 24866 37018
rect 24866 36966 24878 37018
rect 24878 36966 24908 37018
rect 24932 36966 24942 37018
rect 24942 36966 24988 37018
rect 24692 36964 24748 36966
rect 24772 36964 24828 36966
rect 24852 36964 24908 36966
rect 24932 36964 24988 36966
rect 24692 35930 24748 35932
rect 24772 35930 24828 35932
rect 24852 35930 24908 35932
rect 24932 35930 24988 35932
rect 24692 35878 24738 35930
rect 24738 35878 24748 35930
rect 24772 35878 24802 35930
rect 24802 35878 24814 35930
rect 24814 35878 24828 35930
rect 24852 35878 24866 35930
rect 24866 35878 24878 35930
rect 24878 35878 24908 35930
rect 24932 35878 24942 35930
rect 24942 35878 24988 35930
rect 24692 35876 24748 35878
rect 24772 35876 24828 35878
rect 24852 35876 24908 35878
rect 24932 35876 24988 35878
rect 24692 34842 24748 34844
rect 24772 34842 24828 34844
rect 24852 34842 24908 34844
rect 24932 34842 24988 34844
rect 24692 34790 24738 34842
rect 24738 34790 24748 34842
rect 24772 34790 24802 34842
rect 24802 34790 24814 34842
rect 24814 34790 24828 34842
rect 24852 34790 24866 34842
rect 24866 34790 24878 34842
rect 24878 34790 24908 34842
rect 24932 34790 24942 34842
rect 24942 34790 24988 34842
rect 24692 34788 24748 34790
rect 24772 34788 24828 34790
rect 24852 34788 24908 34790
rect 24932 34788 24988 34790
rect 24692 33754 24748 33756
rect 24772 33754 24828 33756
rect 24852 33754 24908 33756
rect 24932 33754 24988 33756
rect 24692 33702 24738 33754
rect 24738 33702 24748 33754
rect 24772 33702 24802 33754
rect 24802 33702 24814 33754
rect 24814 33702 24828 33754
rect 24852 33702 24866 33754
rect 24866 33702 24878 33754
rect 24878 33702 24908 33754
rect 24932 33702 24942 33754
rect 24942 33702 24988 33754
rect 24692 33700 24748 33702
rect 24772 33700 24828 33702
rect 24852 33700 24908 33702
rect 24932 33700 24988 33702
rect 24692 32666 24748 32668
rect 24772 32666 24828 32668
rect 24852 32666 24908 32668
rect 24932 32666 24988 32668
rect 24692 32614 24738 32666
rect 24738 32614 24748 32666
rect 24772 32614 24802 32666
rect 24802 32614 24814 32666
rect 24814 32614 24828 32666
rect 24852 32614 24866 32666
rect 24866 32614 24878 32666
rect 24878 32614 24908 32666
rect 24932 32614 24942 32666
rect 24942 32614 24988 32666
rect 24692 32612 24748 32614
rect 24772 32612 24828 32614
rect 24852 32612 24908 32614
rect 24932 32612 24988 32614
rect 24692 31578 24748 31580
rect 24772 31578 24828 31580
rect 24852 31578 24908 31580
rect 24932 31578 24988 31580
rect 24692 31526 24738 31578
rect 24738 31526 24748 31578
rect 24772 31526 24802 31578
rect 24802 31526 24814 31578
rect 24814 31526 24828 31578
rect 24852 31526 24866 31578
rect 24866 31526 24878 31578
rect 24878 31526 24908 31578
rect 24932 31526 24942 31578
rect 24942 31526 24988 31578
rect 24692 31524 24748 31526
rect 24772 31524 24828 31526
rect 24852 31524 24908 31526
rect 24932 31524 24988 31526
rect 24582 30776 24638 30832
rect 24122 16940 24124 16960
rect 24124 16940 24176 16960
rect 24176 16940 24178 16960
rect 24122 16904 24178 16940
rect 24122 15816 24178 15872
rect 24030 14764 24032 14784
rect 24032 14764 24084 14784
rect 24084 14764 24086 14784
rect 24030 14728 24086 14764
rect 24490 22344 24546 22400
rect 24398 18028 24400 18048
rect 24400 18028 24452 18048
rect 24452 18028 24454 18048
rect 24398 17992 24454 18028
rect 24398 13676 24400 13696
rect 24400 13676 24452 13696
rect 24452 13676 24454 13696
rect 24398 13640 24454 13676
rect 24214 12588 24216 12608
rect 24216 12588 24268 12608
rect 24268 12588 24270 12608
rect 24214 12552 24270 12588
rect 22558 5480 22614 5536
rect 22374 3712 22430 3768
rect 22374 2352 22430 2408
rect 23018 5616 23074 5672
rect 23846 11500 23848 11520
rect 23848 11500 23900 11520
rect 23900 11500 23902 11520
rect 23846 11464 23902 11500
rect 23294 10376 23350 10432
rect 23202 10104 23258 10160
rect 23570 8916 23572 8936
rect 23572 8916 23624 8936
rect 23624 8916 23626 8936
rect 23570 8880 23626 8916
rect 24030 9288 24086 9344
rect 23754 7112 23810 7168
rect 23202 6704 23258 6760
rect 23754 3440 23810 3496
rect 24692 30490 24748 30492
rect 24772 30490 24828 30492
rect 24852 30490 24908 30492
rect 24932 30490 24988 30492
rect 24692 30438 24738 30490
rect 24738 30438 24748 30490
rect 24772 30438 24802 30490
rect 24802 30438 24814 30490
rect 24814 30438 24828 30490
rect 24852 30438 24866 30490
rect 24866 30438 24878 30490
rect 24878 30438 24908 30490
rect 24932 30438 24942 30490
rect 24942 30438 24988 30490
rect 24692 30436 24748 30438
rect 24772 30436 24828 30438
rect 24852 30436 24908 30438
rect 24932 30436 24988 30438
rect 24692 29402 24748 29404
rect 24772 29402 24828 29404
rect 24852 29402 24908 29404
rect 24932 29402 24988 29404
rect 24692 29350 24738 29402
rect 24738 29350 24748 29402
rect 24772 29350 24802 29402
rect 24802 29350 24814 29402
rect 24814 29350 24828 29402
rect 24852 29350 24866 29402
rect 24866 29350 24878 29402
rect 24878 29350 24908 29402
rect 24932 29350 24942 29402
rect 24942 29350 24988 29402
rect 24692 29348 24748 29350
rect 24772 29348 24828 29350
rect 24852 29348 24908 29350
rect 24932 29348 24988 29350
rect 24692 28314 24748 28316
rect 24772 28314 24828 28316
rect 24852 28314 24908 28316
rect 24932 28314 24988 28316
rect 24692 28262 24738 28314
rect 24738 28262 24748 28314
rect 24772 28262 24802 28314
rect 24802 28262 24814 28314
rect 24814 28262 24828 28314
rect 24852 28262 24866 28314
rect 24866 28262 24878 28314
rect 24878 28262 24908 28314
rect 24932 28262 24942 28314
rect 24942 28262 24988 28314
rect 24692 28260 24748 28262
rect 24772 28260 24828 28262
rect 24852 28260 24908 28262
rect 24932 28260 24988 28262
rect 24692 27226 24748 27228
rect 24772 27226 24828 27228
rect 24852 27226 24908 27228
rect 24932 27226 24988 27228
rect 24692 27174 24738 27226
rect 24738 27174 24748 27226
rect 24772 27174 24802 27226
rect 24802 27174 24814 27226
rect 24814 27174 24828 27226
rect 24852 27174 24866 27226
rect 24866 27174 24878 27226
rect 24878 27174 24908 27226
rect 24932 27174 24942 27226
rect 24942 27174 24988 27226
rect 24692 27172 24748 27174
rect 24772 27172 24828 27174
rect 24852 27172 24908 27174
rect 24932 27172 24988 27174
rect 24692 26138 24748 26140
rect 24772 26138 24828 26140
rect 24852 26138 24908 26140
rect 24932 26138 24988 26140
rect 24692 26086 24738 26138
rect 24738 26086 24748 26138
rect 24772 26086 24802 26138
rect 24802 26086 24814 26138
rect 24814 26086 24828 26138
rect 24852 26086 24866 26138
rect 24866 26086 24878 26138
rect 24878 26086 24908 26138
rect 24932 26086 24942 26138
rect 24942 26086 24988 26138
rect 24692 26084 24748 26086
rect 24772 26084 24828 26086
rect 24852 26084 24908 26086
rect 24932 26084 24988 26086
rect 24692 25050 24748 25052
rect 24772 25050 24828 25052
rect 24852 25050 24908 25052
rect 24932 25050 24988 25052
rect 24692 24998 24738 25050
rect 24738 24998 24748 25050
rect 24772 24998 24802 25050
rect 24802 24998 24814 25050
rect 24814 24998 24828 25050
rect 24852 24998 24866 25050
rect 24866 24998 24878 25050
rect 24878 24998 24908 25050
rect 24932 24998 24942 25050
rect 24942 24998 24988 25050
rect 24692 24996 24748 24998
rect 24772 24996 24828 24998
rect 24852 24996 24908 24998
rect 24932 24996 24988 24998
rect 24692 23962 24748 23964
rect 24772 23962 24828 23964
rect 24852 23962 24908 23964
rect 24932 23962 24988 23964
rect 24692 23910 24738 23962
rect 24738 23910 24748 23962
rect 24772 23910 24802 23962
rect 24802 23910 24814 23962
rect 24814 23910 24828 23962
rect 24852 23910 24866 23962
rect 24866 23910 24878 23962
rect 24878 23910 24908 23962
rect 24932 23910 24942 23962
rect 24942 23910 24988 23962
rect 24692 23908 24748 23910
rect 24772 23908 24828 23910
rect 24852 23908 24908 23910
rect 24932 23908 24988 23910
rect 24692 22874 24748 22876
rect 24772 22874 24828 22876
rect 24852 22874 24908 22876
rect 24932 22874 24988 22876
rect 24692 22822 24738 22874
rect 24738 22822 24748 22874
rect 24772 22822 24802 22874
rect 24802 22822 24814 22874
rect 24814 22822 24828 22874
rect 24852 22822 24866 22874
rect 24866 22822 24878 22874
rect 24878 22822 24908 22874
rect 24932 22822 24942 22874
rect 24942 22822 24988 22874
rect 24692 22820 24748 22822
rect 24772 22820 24828 22822
rect 24852 22820 24908 22822
rect 24932 22820 24988 22822
rect 24692 21786 24748 21788
rect 24772 21786 24828 21788
rect 24852 21786 24908 21788
rect 24932 21786 24988 21788
rect 24692 21734 24738 21786
rect 24738 21734 24748 21786
rect 24772 21734 24802 21786
rect 24802 21734 24814 21786
rect 24814 21734 24828 21786
rect 24852 21734 24866 21786
rect 24866 21734 24878 21786
rect 24878 21734 24908 21786
rect 24932 21734 24942 21786
rect 24942 21734 24988 21786
rect 24692 21732 24748 21734
rect 24772 21732 24828 21734
rect 24852 21732 24908 21734
rect 24932 21732 24988 21734
rect 24692 20698 24748 20700
rect 24772 20698 24828 20700
rect 24852 20698 24908 20700
rect 24932 20698 24988 20700
rect 24692 20646 24738 20698
rect 24738 20646 24748 20698
rect 24772 20646 24802 20698
rect 24802 20646 24814 20698
rect 24814 20646 24828 20698
rect 24852 20646 24866 20698
rect 24866 20646 24878 20698
rect 24878 20646 24908 20698
rect 24932 20646 24942 20698
rect 24942 20646 24988 20698
rect 24692 20644 24748 20646
rect 24772 20644 24828 20646
rect 24852 20644 24908 20646
rect 24932 20644 24988 20646
rect 24692 19610 24748 19612
rect 24772 19610 24828 19612
rect 24852 19610 24908 19612
rect 24932 19610 24988 19612
rect 24692 19558 24738 19610
rect 24738 19558 24748 19610
rect 24772 19558 24802 19610
rect 24802 19558 24814 19610
rect 24814 19558 24828 19610
rect 24852 19558 24866 19610
rect 24866 19558 24878 19610
rect 24878 19558 24908 19610
rect 24932 19558 24942 19610
rect 24942 19558 24988 19610
rect 24692 19556 24748 19558
rect 24772 19556 24828 19558
rect 24852 19556 24908 19558
rect 24932 19556 24988 19558
rect 24692 18522 24748 18524
rect 24772 18522 24828 18524
rect 24852 18522 24908 18524
rect 24932 18522 24988 18524
rect 24692 18470 24738 18522
rect 24738 18470 24748 18522
rect 24772 18470 24802 18522
rect 24802 18470 24814 18522
rect 24814 18470 24828 18522
rect 24852 18470 24866 18522
rect 24866 18470 24878 18522
rect 24878 18470 24908 18522
rect 24932 18470 24942 18522
rect 24942 18470 24988 18522
rect 24692 18468 24748 18470
rect 24772 18468 24828 18470
rect 24852 18468 24908 18470
rect 24932 18468 24988 18470
rect 25134 35944 25190 36000
rect 25226 34892 25228 34912
rect 25228 34892 25280 34912
rect 25280 34892 25282 34912
rect 25226 34856 25282 34892
rect 25226 33804 25228 33824
rect 25228 33804 25280 33824
rect 25280 33804 25282 33824
rect 25226 33768 25282 33804
rect 25226 32716 25228 32736
rect 25228 32716 25280 32736
rect 25280 32716 25282 32736
rect 25226 32680 25282 32716
rect 25134 31592 25190 31648
rect 25134 30504 25190 30560
rect 25134 29452 25136 29472
rect 25136 29452 25188 29472
rect 25188 29452 25190 29472
rect 25134 29416 25190 29452
rect 25134 28364 25136 28384
rect 25136 28364 25188 28384
rect 25188 28364 25190 28384
rect 25134 28328 25190 28364
rect 25134 27276 25136 27296
rect 25136 27276 25188 27296
rect 25188 27276 25190 27296
rect 25134 27240 25190 27276
rect 25134 26152 25190 26208
rect 25134 25064 25190 25120
rect 25134 24012 25136 24032
rect 25136 24012 25188 24032
rect 25188 24012 25190 24032
rect 25134 23976 25190 24012
rect 25134 22924 25136 22944
rect 25136 22924 25188 22944
rect 25188 22924 25190 22944
rect 25134 22888 25190 22924
rect 25134 21800 25190 21856
rect 25134 20712 25190 20768
rect 25134 18536 25190 18592
rect 25134 17448 25190 17504
rect 24692 17434 24748 17436
rect 24772 17434 24828 17436
rect 24852 17434 24908 17436
rect 24932 17434 24988 17436
rect 24692 17382 24738 17434
rect 24738 17382 24748 17434
rect 24772 17382 24802 17434
rect 24802 17382 24814 17434
rect 24814 17382 24828 17434
rect 24852 17382 24866 17434
rect 24866 17382 24878 17434
rect 24878 17382 24908 17434
rect 24932 17382 24942 17434
rect 24942 17382 24988 17434
rect 24692 17380 24748 17382
rect 24772 17380 24828 17382
rect 24852 17380 24908 17382
rect 24932 17380 24988 17382
rect 25594 38936 25650 38992
rect 25502 24112 25558 24168
rect 25318 19624 25374 19680
rect 24692 16346 24748 16348
rect 24772 16346 24828 16348
rect 24852 16346 24908 16348
rect 24932 16346 24988 16348
rect 24692 16294 24738 16346
rect 24738 16294 24748 16346
rect 24772 16294 24802 16346
rect 24802 16294 24814 16346
rect 24814 16294 24828 16346
rect 24852 16294 24866 16346
rect 24866 16294 24878 16346
rect 24878 16294 24908 16346
rect 24932 16294 24942 16346
rect 24942 16294 24988 16346
rect 24692 16292 24748 16294
rect 24772 16292 24828 16294
rect 24852 16292 24908 16294
rect 24932 16292 24988 16294
rect 24692 15258 24748 15260
rect 24772 15258 24828 15260
rect 24852 15258 24908 15260
rect 24932 15258 24988 15260
rect 24692 15206 24738 15258
rect 24738 15206 24748 15258
rect 24772 15206 24802 15258
rect 24802 15206 24814 15258
rect 24814 15206 24828 15258
rect 24852 15206 24866 15258
rect 24866 15206 24878 15258
rect 24878 15206 24908 15258
rect 24932 15206 24942 15258
rect 24942 15206 24988 15258
rect 24692 15204 24748 15206
rect 24772 15204 24828 15206
rect 24852 15204 24908 15206
rect 24932 15204 24988 15206
rect 24692 14170 24748 14172
rect 24772 14170 24828 14172
rect 24852 14170 24908 14172
rect 24932 14170 24988 14172
rect 24692 14118 24738 14170
rect 24738 14118 24748 14170
rect 24772 14118 24802 14170
rect 24802 14118 24814 14170
rect 24814 14118 24828 14170
rect 24852 14118 24866 14170
rect 24866 14118 24878 14170
rect 24878 14118 24908 14170
rect 24932 14118 24942 14170
rect 24942 14118 24988 14170
rect 24692 14116 24748 14118
rect 24772 14116 24828 14118
rect 24852 14116 24908 14118
rect 24932 14116 24988 14118
rect 24692 13082 24748 13084
rect 24772 13082 24828 13084
rect 24852 13082 24908 13084
rect 24932 13082 24988 13084
rect 24692 13030 24738 13082
rect 24738 13030 24748 13082
rect 24772 13030 24802 13082
rect 24802 13030 24814 13082
rect 24814 13030 24828 13082
rect 24852 13030 24866 13082
rect 24866 13030 24878 13082
rect 24878 13030 24908 13082
rect 24932 13030 24942 13082
rect 24942 13030 24988 13082
rect 24692 13028 24748 13030
rect 24772 13028 24828 13030
rect 24852 13028 24908 13030
rect 24932 13028 24988 13030
rect 24692 11994 24748 11996
rect 24772 11994 24828 11996
rect 24852 11994 24908 11996
rect 24932 11994 24988 11996
rect 24692 11942 24738 11994
rect 24738 11942 24748 11994
rect 24772 11942 24802 11994
rect 24802 11942 24814 11994
rect 24814 11942 24828 11994
rect 24852 11942 24866 11994
rect 24866 11942 24878 11994
rect 24878 11942 24908 11994
rect 24932 11942 24942 11994
rect 24942 11942 24988 11994
rect 24692 11940 24748 11942
rect 24772 11940 24828 11942
rect 24852 11940 24908 11942
rect 24932 11940 24988 11942
rect 25226 16360 25282 16416
rect 25318 15272 25374 15328
rect 25134 14184 25190 14240
rect 25134 12688 25190 12744
rect 25226 12008 25282 12064
rect 24692 10906 24748 10908
rect 24772 10906 24828 10908
rect 24852 10906 24908 10908
rect 24932 10906 24988 10908
rect 24692 10854 24738 10906
rect 24738 10854 24748 10906
rect 24772 10854 24802 10906
rect 24802 10854 24814 10906
rect 24814 10854 24828 10906
rect 24852 10854 24866 10906
rect 24866 10854 24878 10906
rect 24878 10854 24908 10906
rect 24932 10854 24942 10906
rect 24942 10854 24988 10906
rect 24692 10852 24748 10854
rect 24772 10852 24828 10854
rect 24852 10852 24908 10854
rect 24932 10852 24988 10854
rect 24692 9818 24748 9820
rect 24772 9818 24828 9820
rect 24852 9818 24908 9820
rect 24932 9818 24988 9820
rect 24692 9766 24738 9818
rect 24738 9766 24748 9818
rect 24772 9766 24802 9818
rect 24802 9766 24814 9818
rect 24814 9766 24828 9818
rect 24852 9766 24866 9818
rect 24866 9766 24878 9818
rect 24878 9766 24908 9818
rect 24932 9766 24942 9818
rect 24942 9766 24988 9818
rect 24692 9764 24748 9766
rect 24772 9764 24828 9766
rect 24852 9764 24908 9766
rect 24932 9764 24988 9766
rect 24490 8200 24546 8256
rect 24030 3032 24086 3088
rect 24692 8730 24748 8732
rect 24772 8730 24828 8732
rect 24852 8730 24908 8732
rect 24932 8730 24988 8732
rect 24692 8678 24738 8730
rect 24738 8678 24748 8730
rect 24772 8678 24802 8730
rect 24802 8678 24814 8730
rect 24814 8678 24828 8730
rect 24852 8678 24866 8730
rect 24866 8678 24878 8730
rect 24878 8678 24908 8730
rect 24932 8678 24942 8730
rect 24942 8678 24988 8730
rect 24692 8676 24748 8678
rect 24772 8676 24828 8678
rect 24852 8676 24908 8678
rect 24932 8676 24988 8678
rect 24692 7642 24748 7644
rect 24772 7642 24828 7644
rect 24852 7642 24908 7644
rect 24932 7642 24988 7644
rect 24692 7590 24738 7642
rect 24738 7590 24748 7642
rect 24772 7590 24802 7642
rect 24802 7590 24814 7642
rect 24814 7590 24828 7642
rect 24852 7590 24866 7642
rect 24866 7590 24878 7642
rect 24878 7590 24908 7642
rect 24932 7590 24942 7642
rect 24942 7590 24988 7642
rect 24692 7588 24748 7590
rect 24772 7588 24828 7590
rect 24852 7588 24908 7590
rect 24932 7588 24988 7590
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 25226 10920 25282 10976
rect 25134 9832 25190 9888
rect 25042 5752 25098 5808
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
rect 25226 3712 25282 3768
rect 25502 6840 25558 6896
rect 25594 3576 25650 3632
rect 25502 1128 25558 1184
<< metal3 >>
rect 18454 44508 18460 44572
rect 18524 44570 18530 44572
rect 18597 44570 18663 44573
rect 18524 44568 18663 44570
rect 18524 44512 18602 44568
rect 18658 44512 18663 44568
rect 18524 44510 18663 44512
rect 18524 44508 18530 44510
rect 18597 44507 18663 44510
rect 25840 43618 26000 43648
rect 25086 43558 26000 43618
rect 6880 43552 7196 43553
rect 6880 43488 6886 43552
rect 6950 43488 6966 43552
rect 7030 43488 7046 43552
rect 7110 43488 7126 43552
rect 7190 43488 7196 43552
rect 6880 43487 7196 43488
rect 12814 43552 13130 43553
rect 12814 43488 12820 43552
rect 12884 43488 12900 43552
rect 12964 43488 12980 43552
rect 13044 43488 13060 43552
rect 13124 43488 13130 43552
rect 12814 43487 13130 43488
rect 18748 43552 19064 43553
rect 18748 43488 18754 43552
rect 18818 43488 18834 43552
rect 18898 43488 18914 43552
rect 18978 43488 18994 43552
rect 19058 43488 19064 43552
rect 18748 43487 19064 43488
rect 24682 43552 24998 43553
rect 24682 43488 24688 43552
rect 24752 43488 24768 43552
rect 24832 43488 24848 43552
rect 24912 43488 24928 43552
rect 24992 43488 24998 43552
rect 24682 43487 24998 43488
rect 12893 43346 12959 43349
rect 15510 43346 15516 43348
rect 12893 43344 15516 43346
rect 12893 43288 12898 43344
rect 12954 43288 15516 43344
rect 12893 43286 15516 43288
rect 12893 43283 12959 43286
rect 15510 43284 15516 43286
rect 15580 43284 15586 43348
rect 23197 43346 23263 43349
rect 25086 43346 25146 43558
rect 25840 43528 26000 43558
rect 23197 43344 25146 43346
rect 23197 43288 23202 43344
rect 23258 43288 25146 43344
rect 23197 43286 25146 43288
rect 23197 43283 23263 43286
rect 21582 43148 21588 43212
rect 21652 43210 21658 43212
rect 22921 43210 22987 43213
rect 21652 43208 22987 43210
rect 21652 43152 22926 43208
rect 22982 43152 22987 43208
rect 21652 43150 22987 43152
rect 21652 43148 21658 43150
rect 22921 43147 22987 43150
rect 14590 43012 14596 43076
rect 14660 43074 14666 43076
rect 15285 43074 15351 43077
rect 19241 43074 19307 43077
rect 14660 43072 15351 43074
rect 14660 43016 15290 43072
rect 15346 43016 15351 43072
rect 14660 43014 15351 43016
rect 14660 43012 14666 43014
rect 15285 43011 15351 43014
rect 19198 43072 19307 43074
rect 19198 43016 19246 43072
rect 19302 43016 19307 43072
rect 19198 43011 19307 43016
rect 25313 43074 25379 43077
rect 25840 43074 26000 43104
rect 25313 43072 26000 43074
rect 25313 43016 25318 43072
rect 25374 43016 26000 43072
rect 25313 43014 26000 43016
rect 25313 43011 25379 43014
rect 3913 43008 4229 43009
rect 3913 42944 3919 43008
rect 3983 42944 3999 43008
rect 4063 42944 4079 43008
rect 4143 42944 4159 43008
rect 4223 42944 4229 43008
rect 3913 42943 4229 42944
rect 9847 43008 10163 43009
rect 9847 42944 9853 43008
rect 9917 42944 9933 43008
rect 9997 42944 10013 43008
rect 10077 42944 10093 43008
rect 10157 42944 10163 43008
rect 9847 42943 10163 42944
rect 15781 43008 16097 43009
rect 15781 42944 15787 43008
rect 15851 42944 15867 43008
rect 15931 42944 15947 43008
rect 16011 42944 16027 43008
rect 16091 42944 16097 43008
rect 15781 42943 16097 42944
rect 10358 42876 10364 42940
rect 10428 42938 10434 42940
rect 12525 42938 12591 42941
rect 10428 42936 12591 42938
rect 10428 42880 12530 42936
rect 12586 42880 12591 42936
rect 10428 42878 12591 42880
rect 10428 42876 10434 42878
rect 12525 42875 12591 42878
rect 13302 42876 13308 42940
rect 13372 42938 13378 42940
rect 14273 42938 14339 42941
rect 13372 42936 14339 42938
rect 13372 42880 14278 42936
rect 14334 42880 14339 42936
rect 13372 42878 14339 42880
rect 13372 42876 13378 42878
rect 14273 42875 14339 42878
rect 14917 42940 14983 42941
rect 14917 42936 14964 42940
rect 15028 42938 15034 42940
rect 14917 42880 14922 42936
rect 14917 42876 14964 42880
rect 15028 42878 15074 42938
rect 15028 42876 15034 42878
rect 14917 42875 14983 42876
rect 8845 42666 8911 42669
rect 15469 42666 15535 42669
rect 8845 42664 15535 42666
rect 8845 42608 8850 42664
rect 8906 42608 15474 42664
rect 15530 42608 15535 42664
rect 8845 42606 15535 42608
rect 8845 42603 8911 42606
rect 15469 42603 15535 42606
rect 18413 42666 18479 42669
rect 18873 42666 18939 42669
rect 18413 42664 18939 42666
rect 18413 42608 18418 42664
rect 18474 42608 18878 42664
rect 18934 42608 18939 42664
rect 18413 42606 18939 42608
rect 18413 42603 18479 42606
rect 18873 42603 18939 42606
rect 6880 42464 7196 42465
rect 6880 42400 6886 42464
rect 6950 42400 6966 42464
rect 7030 42400 7046 42464
rect 7110 42400 7126 42464
rect 7190 42400 7196 42464
rect 6880 42399 7196 42400
rect 12814 42464 13130 42465
rect 12814 42400 12820 42464
rect 12884 42400 12900 42464
rect 12964 42400 12980 42464
rect 13044 42400 13060 42464
rect 13124 42400 13130 42464
rect 12814 42399 13130 42400
rect 18748 42464 19064 42465
rect 18748 42400 18754 42464
rect 18818 42400 18834 42464
rect 18898 42400 18914 42464
rect 18978 42400 18994 42464
rect 19058 42400 19064 42464
rect 18748 42399 19064 42400
rect 2037 42394 2103 42397
rect 5809 42394 5875 42397
rect 2037 42392 5875 42394
rect 2037 42336 2042 42392
rect 2098 42336 5814 42392
rect 5870 42336 5875 42392
rect 2037 42334 5875 42336
rect 2037 42331 2103 42334
rect 5809 42331 5875 42334
rect 19198 42261 19258 43011
rect 21715 43008 22031 43009
rect 21715 42944 21721 43008
rect 21785 42944 21801 43008
rect 21865 42944 21881 43008
rect 21945 42944 21961 43008
rect 22025 42944 22031 43008
rect 25840 42984 26000 43014
rect 21715 42943 22031 42944
rect 25129 42530 25195 42533
rect 25840 42530 26000 42560
rect 25129 42528 26000 42530
rect 25129 42472 25134 42528
rect 25190 42472 26000 42528
rect 25129 42470 26000 42472
rect 25129 42467 25195 42470
rect 24682 42464 24998 42465
rect 24682 42400 24688 42464
rect 24752 42400 24768 42464
rect 24832 42400 24848 42464
rect 24912 42400 24928 42464
rect 24992 42400 24998 42464
rect 25840 42440 26000 42470
rect 24682 42399 24998 42400
rect 1158 42196 1164 42260
rect 1228 42258 1234 42260
rect 4705 42258 4771 42261
rect 1228 42256 4771 42258
rect 1228 42200 4710 42256
rect 4766 42200 4771 42256
rect 1228 42198 4771 42200
rect 1228 42196 1234 42198
rect 4705 42195 4771 42198
rect 9489 42258 9555 42261
rect 9857 42258 9923 42261
rect 9489 42256 17970 42258
rect 9489 42200 9494 42256
rect 9550 42200 9862 42256
rect 9918 42200 17970 42256
rect 9489 42198 17970 42200
rect 9489 42195 9555 42198
rect 9857 42195 9923 42198
rect 3417 42122 3483 42125
rect 3969 42122 4035 42125
rect 3417 42120 4035 42122
rect 3417 42064 3422 42120
rect 3478 42064 3974 42120
rect 4030 42064 4035 42120
rect 3417 42062 4035 42064
rect 3417 42059 3483 42062
rect 3969 42059 4035 42062
rect 7097 42122 7163 42125
rect 10317 42122 10383 42125
rect 7097 42120 10383 42122
rect 7097 42064 7102 42120
rect 7158 42064 10322 42120
rect 10378 42064 10383 42120
rect 7097 42062 10383 42064
rect 7097 42059 7163 42062
rect 10317 42059 10383 42062
rect 11646 42060 11652 42124
rect 11716 42122 11722 42124
rect 12065 42122 12131 42125
rect 11716 42120 12131 42122
rect 11716 42064 12070 42120
rect 12126 42064 12131 42120
rect 11716 42062 12131 42064
rect 17910 42122 17970 42198
rect 18454 42196 18460 42260
rect 18524 42258 18530 42260
rect 18965 42258 19031 42261
rect 18524 42256 19031 42258
rect 18524 42200 18970 42256
rect 19026 42200 19031 42256
rect 18524 42198 19031 42200
rect 19198 42256 19307 42261
rect 19198 42200 19246 42256
rect 19302 42200 19307 42256
rect 19198 42198 19307 42200
rect 18524 42196 18530 42198
rect 18965 42195 19031 42198
rect 19241 42195 19307 42198
rect 20069 42258 20135 42261
rect 20621 42258 20687 42261
rect 20069 42256 20687 42258
rect 20069 42200 20074 42256
rect 20130 42200 20626 42256
rect 20682 42200 20687 42256
rect 20069 42198 20687 42200
rect 20069 42195 20135 42198
rect 20621 42195 20687 42198
rect 20662 42122 20668 42124
rect 17910 42062 20668 42122
rect 11716 42060 11722 42062
rect 12065 42059 12131 42062
rect 20662 42060 20668 42062
rect 20732 42060 20738 42124
rect 11789 41988 11855 41989
rect 11789 41984 11836 41988
rect 11900 41986 11906 41988
rect 24117 41986 24183 41989
rect 25840 41986 26000 42016
rect 11789 41928 11794 41984
rect 11789 41924 11836 41928
rect 11900 41926 11946 41986
rect 24117 41984 26000 41986
rect 24117 41928 24122 41984
rect 24178 41928 26000 41984
rect 24117 41926 26000 41928
rect 11900 41924 11906 41926
rect 11789 41923 11855 41924
rect 24117 41923 24183 41926
rect 3913 41920 4229 41921
rect 3913 41856 3919 41920
rect 3983 41856 3999 41920
rect 4063 41856 4079 41920
rect 4143 41856 4159 41920
rect 4223 41856 4229 41920
rect 3913 41855 4229 41856
rect 9847 41920 10163 41921
rect 9847 41856 9853 41920
rect 9917 41856 9933 41920
rect 9997 41856 10013 41920
rect 10077 41856 10093 41920
rect 10157 41856 10163 41920
rect 9847 41855 10163 41856
rect 15781 41920 16097 41921
rect 15781 41856 15787 41920
rect 15851 41856 15867 41920
rect 15931 41856 15947 41920
rect 16011 41856 16027 41920
rect 16091 41856 16097 41920
rect 15781 41855 16097 41856
rect 21715 41920 22031 41921
rect 21715 41856 21721 41920
rect 21785 41856 21801 41920
rect 21865 41856 21881 41920
rect 21945 41856 21961 41920
rect 22025 41856 22031 41920
rect 25840 41896 26000 41926
rect 21715 41855 22031 41856
rect 6269 41852 6335 41853
rect 6269 41850 6316 41852
rect 6224 41848 6316 41850
rect 6224 41792 6274 41848
rect 6224 41790 6316 41792
rect 6269 41788 6316 41790
rect 6380 41788 6386 41852
rect 7465 41850 7531 41853
rect 8201 41852 8267 41853
rect 7598 41850 7604 41852
rect 7465 41848 7604 41850
rect 7465 41792 7470 41848
rect 7526 41792 7604 41848
rect 7465 41790 7604 41792
rect 6269 41787 6335 41788
rect 7465 41787 7531 41790
rect 7598 41788 7604 41790
rect 7668 41788 7674 41852
rect 8150 41850 8156 41852
rect 8110 41790 8156 41850
rect 8220 41848 8267 41852
rect 8262 41792 8267 41848
rect 8150 41788 8156 41790
rect 8220 41788 8267 41792
rect 8201 41787 8267 41788
rect 17309 41850 17375 41853
rect 17309 41848 19810 41850
rect 17309 41792 17314 41848
rect 17370 41792 19810 41848
rect 17309 41790 19810 41792
rect 17309 41787 17375 41790
rect 16941 41716 17007 41717
rect 17677 41716 17743 41717
rect 18321 41716 18387 41717
rect 16941 41712 16988 41716
rect 17052 41714 17058 41716
rect 16941 41656 16946 41712
rect 16941 41652 16988 41656
rect 17052 41654 17098 41714
rect 17677 41712 17724 41716
rect 17788 41714 17794 41716
rect 18270 41714 18276 41716
rect 17677 41656 17682 41712
rect 17052 41652 17058 41654
rect 17677 41652 17724 41656
rect 17788 41654 17834 41714
rect 18230 41654 18276 41714
rect 18340 41712 18387 41716
rect 18382 41656 18387 41712
rect 17788 41652 17794 41654
rect 18270 41652 18276 41654
rect 18340 41652 18387 41656
rect 16941 41651 17007 41652
rect 17677 41651 17743 41652
rect 18321 41651 18387 41652
rect 19517 41716 19583 41717
rect 19517 41712 19564 41716
rect 19628 41714 19634 41716
rect 19750 41714 19810 41790
rect 19517 41656 19522 41712
rect 19517 41652 19564 41656
rect 19628 41654 19674 41714
rect 19750 41654 22754 41714
rect 19628 41652 19634 41654
rect 19517 41651 19583 41652
rect 473 41578 539 41581
rect 9581 41578 9647 41581
rect 473 41576 9647 41578
rect 473 41520 478 41576
rect 534 41520 9586 41576
rect 9642 41520 9647 41576
rect 473 41518 9647 41520
rect 473 41515 539 41518
rect 9581 41515 9647 41518
rect 9765 41578 9831 41581
rect 17033 41578 17099 41581
rect 9765 41576 17099 41578
rect 9765 41520 9770 41576
rect 9826 41520 17038 41576
rect 17094 41520 17099 41576
rect 9765 41518 17099 41520
rect 9765 41515 9831 41518
rect 17033 41515 17099 41518
rect 18229 41578 18295 41581
rect 19701 41578 19767 41581
rect 18229 41576 19767 41578
rect 18229 41520 18234 41576
rect 18290 41520 19706 41576
rect 19762 41520 19767 41576
rect 18229 41518 19767 41520
rect 18229 41515 18295 41518
rect 19701 41515 19767 41518
rect 20989 41578 21055 41581
rect 22553 41578 22619 41581
rect 20989 41576 22619 41578
rect 20989 41520 20994 41576
rect 21050 41520 22558 41576
rect 22614 41520 22619 41576
rect 20989 41518 22619 41520
rect 20989 41515 21055 41518
rect 22553 41515 22619 41518
rect 974 41380 980 41444
rect 1044 41442 1050 41444
rect 2865 41442 2931 41445
rect 1044 41440 2931 41442
rect 1044 41384 2870 41440
rect 2926 41384 2931 41440
rect 1044 41382 2931 41384
rect 1044 41380 1050 41382
rect 2865 41379 2931 41382
rect 18413 41444 18479 41445
rect 18413 41440 18460 41444
rect 18524 41442 18530 41444
rect 20713 41442 20779 41445
rect 21817 41442 21883 41445
rect 18413 41384 18418 41440
rect 18413 41380 18460 41384
rect 18524 41382 18570 41442
rect 20713 41440 21883 41442
rect 20713 41384 20718 41440
rect 20774 41384 21822 41440
rect 21878 41384 21883 41440
rect 20713 41382 21883 41384
rect 22694 41442 22754 41654
rect 23197 41442 23263 41445
rect 22694 41440 23263 41442
rect 22694 41384 23202 41440
rect 23258 41384 23263 41440
rect 22694 41382 23263 41384
rect 18524 41380 18530 41382
rect 18413 41379 18479 41380
rect 20713 41379 20779 41382
rect 21817 41379 21883 41382
rect 23197 41379 23263 41382
rect 25129 41442 25195 41445
rect 25840 41442 26000 41472
rect 25129 41440 26000 41442
rect 25129 41384 25134 41440
rect 25190 41384 26000 41440
rect 25129 41382 26000 41384
rect 25129 41379 25195 41382
rect 6880 41376 7196 41377
rect 6880 41312 6886 41376
rect 6950 41312 6966 41376
rect 7030 41312 7046 41376
rect 7110 41312 7126 41376
rect 7190 41312 7196 41376
rect 6880 41311 7196 41312
rect 12814 41376 13130 41377
rect 12814 41312 12820 41376
rect 12884 41312 12900 41376
rect 12964 41312 12980 41376
rect 13044 41312 13060 41376
rect 13124 41312 13130 41376
rect 12814 41311 13130 41312
rect 18748 41376 19064 41377
rect 18748 41312 18754 41376
rect 18818 41312 18834 41376
rect 18898 41312 18914 41376
rect 18978 41312 18994 41376
rect 19058 41312 19064 41376
rect 18748 41311 19064 41312
rect 24682 41376 24998 41377
rect 24682 41312 24688 41376
rect 24752 41312 24768 41376
rect 24832 41312 24848 41376
rect 24912 41312 24928 41376
rect 24992 41312 24998 41376
rect 25840 41352 26000 41382
rect 24682 41311 24998 41312
rect 19793 41306 19859 41309
rect 22921 41306 22987 41309
rect 19793 41304 22987 41306
rect 19793 41248 19798 41304
rect 19854 41248 22926 41304
rect 22982 41248 22987 41304
rect 19793 41246 22987 41248
rect 19793 41243 19859 41246
rect 22921 41243 22987 41246
rect 2221 41170 2287 41173
rect 18413 41170 18479 41173
rect 21817 41170 21883 41173
rect 2221 41168 21883 41170
rect 2221 41112 2226 41168
rect 2282 41112 18418 41168
rect 18474 41112 21822 41168
rect 21878 41112 21883 41168
rect 2221 41110 21883 41112
rect 2221 41107 2287 41110
rect 18413 41107 18479 41110
rect 21817 41107 21883 41110
rect 10409 41034 10475 41037
rect 20897 41034 20963 41037
rect 10409 41032 20963 41034
rect 10409 40976 10414 41032
rect 10470 40976 20902 41032
rect 20958 40976 20963 41032
rect 10409 40974 20963 40976
rect 10409 40971 10475 40974
rect 20897 40971 20963 40974
rect 21449 41034 21515 41037
rect 21582 41034 21588 41036
rect 21449 41032 21588 41034
rect 21449 40976 21454 41032
rect 21510 40976 21588 41032
rect 21449 40974 21588 40976
rect 21449 40971 21515 40974
rect 21582 40972 21588 40974
rect 21652 40972 21658 41036
rect 22185 41034 22251 41037
rect 22461 41034 22527 41037
rect 22185 41032 22527 41034
rect 22185 40976 22190 41032
rect 22246 40976 22466 41032
rect 22522 40976 22527 41032
rect 22185 40974 22527 40976
rect 22185 40971 22251 40974
rect 22461 40971 22527 40974
rect 23657 40898 23723 40901
rect 25840 40898 26000 40928
rect 23657 40896 26000 40898
rect 23657 40840 23662 40896
rect 23718 40840 26000 40896
rect 23657 40838 26000 40840
rect 23657 40835 23723 40838
rect 3913 40832 4229 40833
rect 3913 40768 3919 40832
rect 3983 40768 3999 40832
rect 4063 40768 4079 40832
rect 4143 40768 4159 40832
rect 4223 40768 4229 40832
rect 3913 40767 4229 40768
rect 9847 40832 10163 40833
rect 9847 40768 9853 40832
rect 9917 40768 9933 40832
rect 9997 40768 10013 40832
rect 10077 40768 10093 40832
rect 10157 40768 10163 40832
rect 9847 40767 10163 40768
rect 15781 40832 16097 40833
rect 15781 40768 15787 40832
rect 15851 40768 15867 40832
rect 15931 40768 15947 40832
rect 16011 40768 16027 40832
rect 16091 40768 16097 40832
rect 15781 40767 16097 40768
rect 21715 40832 22031 40833
rect 21715 40768 21721 40832
rect 21785 40768 21801 40832
rect 21865 40768 21881 40832
rect 21945 40768 21961 40832
rect 22025 40768 22031 40832
rect 25840 40808 26000 40838
rect 21715 40767 22031 40768
rect 22093 40762 22159 40765
rect 22461 40762 22527 40765
rect 22093 40760 22527 40762
rect 22093 40704 22098 40760
rect 22154 40704 22466 40760
rect 22522 40704 22527 40760
rect 22093 40702 22527 40704
rect 22093 40699 22159 40702
rect 22461 40699 22527 40702
rect 606 40564 612 40628
rect 676 40626 682 40628
rect 4889 40626 4955 40629
rect 676 40624 4955 40626
rect 676 40568 4894 40624
rect 4950 40568 4955 40624
rect 676 40566 4955 40568
rect 676 40564 682 40566
rect 4889 40563 4955 40566
rect 5625 40626 5691 40629
rect 9489 40626 9555 40629
rect 5625 40624 9555 40626
rect 5625 40568 5630 40624
rect 5686 40568 9494 40624
rect 9550 40568 9555 40624
rect 5625 40566 9555 40568
rect 5625 40563 5691 40566
rect 9489 40563 9555 40566
rect 15101 40626 15167 40629
rect 22645 40626 22711 40629
rect 15101 40624 22711 40626
rect 15101 40568 15106 40624
rect 15162 40568 22650 40624
rect 22706 40568 22711 40624
rect 15101 40566 22711 40568
rect 15101 40563 15167 40566
rect 22645 40563 22711 40566
rect 7281 40490 7347 40493
rect 21633 40490 21699 40493
rect 7281 40488 21699 40490
rect 7281 40432 7286 40488
rect 7342 40432 21638 40488
rect 21694 40432 21699 40488
rect 7281 40430 21699 40432
rect 7281 40427 7347 40430
rect 21633 40427 21699 40430
rect 22093 40490 22159 40493
rect 23473 40490 23539 40493
rect 22093 40488 23539 40490
rect 22093 40432 22098 40488
rect 22154 40432 23478 40488
rect 23534 40432 23539 40488
rect 22093 40430 23539 40432
rect 22093 40427 22159 40430
rect 23473 40427 23539 40430
rect 790 40292 796 40356
rect 860 40354 866 40356
rect 4245 40354 4311 40357
rect 860 40352 4311 40354
rect 860 40296 4250 40352
rect 4306 40296 4311 40352
rect 860 40294 4311 40296
rect 860 40292 866 40294
rect 4245 40291 4311 40294
rect 20253 40354 20319 40357
rect 23657 40354 23723 40357
rect 20253 40352 23723 40354
rect 20253 40296 20258 40352
rect 20314 40296 23662 40352
rect 23718 40296 23723 40352
rect 20253 40294 23723 40296
rect 20253 40291 20319 40294
rect 23657 40291 23723 40294
rect 25129 40354 25195 40357
rect 25840 40354 26000 40384
rect 25129 40352 26000 40354
rect 25129 40296 25134 40352
rect 25190 40296 26000 40352
rect 25129 40294 26000 40296
rect 25129 40291 25195 40294
rect 6880 40288 7196 40289
rect 6880 40224 6886 40288
rect 6950 40224 6966 40288
rect 7030 40224 7046 40288
rect 7110 40224 7126 40288
rect 7190 40224 7196 40288
rect 6880 40223 7196 40224
rect 12814 40288 13130 40289
rect 12814 40224 12820 40288
rect 12884 40224 12900 40288
rect 12964 40224 12980 40288
rect 13044 40224 13060 40288
rect 13124 40224 13130 40288
rect 12814 40223 13130 40224
rect 18748 40288 19064 40289
rect 18748 40224 18754 40288
rect 18818 40224 18834 40288
rect 18898 40224 18914 40288
rect 18978 40224 18994 40288
rect 19058 40224 19064 40288
rect 18748 40223 19064 40224
rect 24682 40288 24998 40289
rect 24682 40224 24688 40288
rect 24752 40224 24768 40288
rect 24832 40224 24848 40288
rect 24912 40224 24928 40288
rect 24992 40224 24998 40288
rect 25840 40264 26000 40294
rect 24682 40223 24998 40224
rect 2630 40156 2636 40220
rect 2700 40218 2706 40220
rect 5349 40218 5415 40221
rect 2700 40216 5415 40218
rect 2700 40160 5354 40216
rect 5410 40160 5415 40216
rect 2700 40158 5415 40160
rect 2700 40156 2706 40158
rect 5349 40155 5415 40158
rect 21817 40218 21883 40221
rect 23933 40218 23999 40221
rect 21817 40216 23999 40218
rect 21817 40160 21822 40216
rect 21878 40160 23938 40216
rect 23994 40160 23999 40216
rect 21817 40158 23999 40160
rect 21817 40155 21883 40158
rect 23933 40155 23999 40158
rect 3233 40082 3299 40085
rect 3366 40082 3372 40084
rect 3233 40080 3372 40082
rect 3233 40024 3238 40080
rect 3294 40024 3372 40080
rect 3233 40022 3372 40024
rect 3233 40019 3299 40022
rect 3366 40020 3372 40022
rect 3436 40020 3442 40084
rect 7741 40082 7807 40085
rect 9622 40082 9628 40084
rect 7741 40080 9628 40082
rect 7741 40024 7746 40080
rect 7802 40024 9628 40080
rect 7741 40022 9628 40024
rect 7741 40019 7807 40022
rect 9622 40020 9628 40022
rect 9692 40020 9698 40084
rect 21909 40082 21975 40085
rect 22645 40082 22711 40085
rect 23105 40082 23171 40085
rect 21909 40080 22711 40082
rect 21909 40024 21914 40080
rect 21970 40024 22650 40080
rect 22706 40024 22711 40080
rect 21909 40022 22711 40024
rect 21909 40019 21975 40022
rect 22645 40019 22711 40022
rect 22878 40080 23171 40082
rect 22878 40024 23110 40080
rect 23166 40024 23171 40080
rect 22878 40022 23171 40024
rect 1209 39946 1275 39949
rect 798 39944 1275 39946
rect 798 39888 1214 39944
rect 1270 39888 1275 39944
rect 798 39886 1275 39888
rect 0 39538 160 39568
rect 798 39538 858 39886
rect 1209 39883 1275 39886
rect 20069 39946 20135 39949
rect 22878 39946 22938 40022
rect 23105 40019 23171 40022
rect 20069 39944 22938 39946
rect 20069 39888 20074 39944
rect 20130 39888 22938 39944
rect 20069 39886 22938 39888
rect 20069 39883 20135 39886
rect 24393 39810 24459 39813
rect 25840 39810 26000 39840
rect 24393 39808 26000 39810
rect 24393 39752 24398 39808
rect 24454 39752 26000 39808
rect 24393 39750 26000 39752
rect 24393 39747 24459 39750
rect 3913 39744 4229 39745
rect 3913 39680 3919 39744
rect 3983 39680 3999 39744
rect 4063 39680 4079 39744
rect 4143 39680 4159 39744
rect 4223 39680 4229 39744
rect 3913 39679 4229 39680
rect 9847 39744 10163 39745
rect 9847 39680 9853 39744
rect 9917 39680 9933 39744
rect 9997 39680 10013 39744
rect 10077 39680 10093 39744
rect 10157 39680 10163 39744
rect 9847 39679 10163 39680
rect 15781 39744 16097 39745
rect 15781 39680 15787 39744
rect 15851 39680 15867 39744
rect 15931 39680 15947 39744
rect 16011 39680 16027 39744
rect 16091 39680 16097 39744
rect 15781 39679 16097 39680
rect 21715 39744 22031 39745
rect 21715 39680 21721 39744
rect 21785 39680 21801 39744
rect 21865 39680 21881 39744
rect 21945 39680 21961 39744
rect 22025 39680 22031 39744
rect 25840 39720 26000 39750
rect 21715 39679 22031 39680
rect 2221 39676 2287 39677
rect 2221 39674 2268 39676
rect 2140 39672 2268 39674
rect 2332 39674 2338 39676
rect 3785 39674 3851 39677
rect 2332 39672 3851 39674
rect 2140 39616 2226 39672
rect 2332 39616 3790 39672
rect 3846 39616 3851 39672
rect 2140 39614 2268 39616
rect 2221 39612 2268 39614
rect 2332 39614 3851 39616
rect 2332 39612 2338 39614
rect 2221 39611 2287 39612
rect 3785 39611 3851 39614
rect 0 39478 858 39538
rect 7557 39538 7623 39541
rect 16430 39538 16436 39540
rect 7557 39536 16436 39538
rect 7557 39480 7562 39536
rect 7618 39480 16436 39536
rect 7557 39478 16436 39480
rect 0 39448 160 39478
rect 7557 39475 7623 39478
rect 16430 39476 16436 39478
rect 16500 39538 16506 39540
rect 23381 39538 23447 39541
rect 16500 39536 23447 39538
rect 16500 39480 23386 39536
rect 23442 39480 23447 39536
rect 16500 39478 23447 39480
rect 16500 39476 16506 39478
rect 23381 39475 23447 39478
rect 1393 39400 1459 39405
rect 1393 39344 1398 39400
rect 1454 39344 1459 39400
rect 1393 39339 1459 39344
rect 1669 39402 1735 39405
rect 12566 39402 12572 39404
rect 1669 39400 12572 39402
rect 1669 39344 1674 39400
rect 1730 39344 12572 39400
rect 1669 39342 12572 39344
rect 1669 39339 1735 39342
rect 12566 39340 12572 39342
rect 12636 39340 12642 39404
rect 21081 39402 21147 39405
rect 24117 39402 24183 39405
rect 21081 39400 24183 39402
rect 21081 39344 21086 39400
rect 21142 39344 24122 39400
rect 24178 39344 24183 39400
rect 21081 39342 24183 39344
rect 21081 39339 21147 39342
rect 24117 39339 24183 39342
rect 0 39266 160 39296
rect 1396 39266 1456 39339
rect 0 39206 1456 39266
rect 21357 39266 21423 39269
rect 23105 39266 23171 39269
rect 21357 39264 23171 39266
rect 21357 39208 21362 39264
rect 21418 39208 23110 39264
rect 23166 39208 23171 39264
rect 21357 39206 23171 39208
rect 0 39176 160 39206
rect 21357 39203 21423 39206
rect 23105 39203 23171 39206
rect 25221 39266 25287 39269
rect 25840 39266 26000 39296
rect 25221 39264 26000 39266
rect 25221 39208 25226 39264
rect 25282 39208 26000 39264
rect 25221 39206 26000 39208
rect 25221 39203 25287 39206
rect 6880 39200 7196 39201
rect 6880 39136 6886 39200
rect 6950 39136 6966 39200
rect 7030 39136 7046 39200
rect 7110 39136 7126 39200
rect 7190 39136 7196 39200
rect 6880 39135 7196 39136
rect 12814 39200 13130 39201
rect 12814 39136 12820 39200
rect 12884 39136 12900 39200
rect 12964 39136 12980 39200
rect 13044 39136 13060 39200
rect 13124 39136 13130 39200
rect 12814 39135 13130 39136
rect 18748 39200 19064 39201
rect 18748 39136 18754 39200
rect 18818 39136 18834 39200
rect 18898 39136 18914 39200
rect 18978 39136 18994 39200
rect 19058 39136 19064 39200
rect 18748 39135 19064 39136
rect 24682 39200 24998 39201
rect 24682 39136 24688 39200
rect 24752 39136 24768 39200
rect 24832 39136 24848 39200
rect 24912 39136 24928 39200
rect 24992 39136 24998 39200
rect 25840 39176 26000 39206
rect 24682 39135 24998 39136
rect 19793 39130 19859 39133
rect 23013 39130 23079 39133
rect 19793 39128 23079 39130
rect 19793 39072 19798 39128
rect 19854 39072 23018 39128
rect 23074 39072 23079 39128
rect 19793 39070 23079 39072
rect 19793 39067 19859 39070
rect 23013 39067 23079 39070
rect 0 38994 160 39024
rect 2773 38994 2839 38997
rect 0 38992 2839 38994
rect 0 38936 2778 38992
rect 2834 38936 2839 38992
rect 0 38934 2839 38936
rect 0 38904 160 38934
rect 2773 38931 2839 38934
rect 11973 38994 12039 38997
rect 25589 38994 25655 38997
rect 11973 38992 25655 38994
rect 11973 38936 11978 38992
rect 12034 38936 25594 38992
rect 25650 38936 25655 38992
rect 11973 38934 25655 38936
rect 11973 38931 12039 38934
rect 25589 38931 25655 38934
rect 3877 38858 3943 38861
rect 4337 38860 4403 38861
rect 4286 38858 4292 38860
rect 2730 38856 3943 38858
rect 2730 38800 3882 38856
rect 3938 38800 3943 38856
rect 2730 38798 3943 38800
rect 4246 38798 4292 38858
rect 4356 38856 4403 38860
rect 4398 38800 4403 38856
rect 0 38722 160 38752
rect 2730 38722 2790 38798
rect 3877 38795 3943 38798
rect 4286 38796 4292 38798
rect 4356 38796 4403 38800
rect 4337 38795 4403 38796
rect 10777 38858 10843 38861
rect 19742 38858 19748 38860
rect 10777 38856 19748 38858
rect 10777 38800 10782 38856
rect 10838 38800 19748 38856
rect 10777 38798 19748 38800
rect 10777 38795 10843 38798
rect 19742 38796 19748 38798
rect 19812 38796 19818 38860
rect 0 38662 2790 38722
rect 19425 38722 19491 38725
rect 20110 38722 20116 38724
rect 19425 38720 20116 38722
rect 19425 38664 19430 38720
rect 19486 38664 20116 38720
rect 19425 38662 20116 38664
rect 0 38632 160 38662
rect 19425 38659 19491 38662
rect 20110 38660 20116 38662
rect 20180 38660 20186 38724
rect 24393 38722 24459 38725
rect 25840 38722 26000 38752
rect 24393 38720 26000 38722
rect 24393 38664 24398 38720
rect 24454 38664 26000 38720
rect 24393 38662 26000 38664
rect 24393 38659 24459 38662
rect 3913 38656 4229 38657
rect 3913 38592 3919 38656
rect 3983 38592 3999 38656
rect 4063 38592 4079 38656
rect 4143 38592 4159 38656
rect 4223 38592 4229 38656
rect 3913 38591 4229 38592
rect 9847 38656 10163 38657
rect 9847 38592 9853 38656
rect 9917 38592 9933 38656
rect 9997 38592 10013 38656
rect 10077 38592 10093 38656
rect 10157 38592 10163 38656
rect 9847 38591 10163 38592
rect 15781 38656 16097 38657
rect 15781 38592 15787 38656
rect 15851 38592 15867 38656
rect 15931 38592 15947 38656
rect 16011 38592 16027 38656
rect 16091 38592 16097 38656
rect 15781 38591 16097 38592
rect 21715 38656 22031 38657
rect 21715 38592 21721 38656
rect 21785 38592 21801 38656
rect 21865 38592 21881 38656
rect 21945 38592 21961 38656
rect 22025 38592 22031 38656
rect 25840 38632 26000 38662
rect 21715 38591 22031 38592
rect 2078 38524 2084 38588
rect 2148 38586 2154 38588
rect 8201 38586 8267 38589
rect 9673 38586 9739 38589
rect 2148 38526 3848 38586
rect 2148 38524 2154 38526
rect 0 38450 160 38480
rect 3049 38450 3115 38453
rect 0 38448 3115 38450
rect 0 38392 3054 38448
rect 3110 38392 3115 38448
rect 0 38390 3115 38392
rect 3788 38450 3848 38526
rect 8201 38584 9739 38586
rect 8201 38528 8206 38584
rect 8262 38528 9678 38584
rect 9734 38528 9739 38584
rect 8201 38526 9739 38528
rect 8201 38523 8267 38526
rect 9673 38523 9739 38526
rect 4613 38450 4679 38453
rect 3788 38448 4679 38450
rect 3788 38392 4618 38448
rect 4674 38392 4679 38448
rect 3788 38390 4679 38392
rect 0 38360 160 38390
rect 3049 38387 3115 38390
rect 4613 38387 4679 38390
rect 4429 38314 4495 38317
rect 13854 38314 13860 38316
rect 4429 38312 13860 38314
rect 4429 38256 4434 38312
rect 4490 38256 13860 38312
rect 4429 38254 13860 38256
rect 4429 38251 4495 38254
rect 13854 38252 13860 38254
rect 13924 38252 13930 38316
rect 0 38178 160 38208
rect 1209 38178 1275 38181
rect 0 38176 1275 38178
rect 0 38120 1214 38176
rect 1270 38120 1275 38176
rect 0 38118 1275 38120
rect 0 38088 160 38118
rect 1209 38115 1275 38118
rect 25221 38178 25287 38181
rect 25840 38178 26000 38208
rect 25221 38176 26000 38178
rect 25221 38120 25226 38176
rect 25282 38120 26000 38176
rect 25221 38118 26000 38120
rect 25221 38115 25287 38118
rect 6880 38112 7196 38113
rect 6880 38048 6886 38112
rect 6950 38048 6966 38112
rect 7030 38048 7046 38112
rect 7110 38048 7126 38112
rect 7190 38048 7196 38112
rect 6880 38047 7196 38048
rect 12814 38112 13130 38113
rect 12814 38048 12820 38112
rect 12884 38048 12900 38112
rect 12964 38048 12980 38112
rect 13044 38048 13060 38112
rect 13124 38048 13130 38112
rect 12814 38047 13130 38048
rect 18748 38112 19064 38113
rect 18748 38048 18754 38112
rect 18818 38048 18834 38112
rect 18898 38048 18914 38112
rect 18978 38048 18994 38112
rect 19058 38048 19064 38112
rect 18748 38047 19064 38048
rect 24682 38112 24998 38113
rect 24682 38048 24688 38112
rect 24752 38048 24768 38112
rect 24832 38048 24848 38112
rect 24912 38048 24928 38112
rect 24992 38048 24998 38112
rect 25840 38088 26000 38118
rect 24682 38047 24998 38048
rect 0 37906 160 37936
rect 749 37906 815 37909
rect 3417 37906 3483 37909
rect 0 37904 815 37906
rect 0 37848 754 37904
rect 810 37848 815 37904
rect 0 37846 815 37848
rect 0 37816 160 37846
rect 749 37843 815 37846
rect 1396 37904 3483 37906
rect 1396 37848 3422 37904
rect 3478 37848 3483 37904
rect 1396 37846 3483 37848
rect 0 37634 160 37664
rect 1396 37634 1456 37846
rect 3417 37843 3483 37846
rect 2221 37770 2287 37773
rect 14457 37770 14523 37773
rect 2221 37768 14523 37770
rect 2221 37712 2226 37768
rect 2282 37712 14462 37768
rect 14518 37712 14523 37768
rect 2221 37710 14523 37712
rect 2221 37707 2287 37710
rect 6686 37637 6746 37710
rect 14457 37707 14523 37710
rect 0 37574 1456 37634
rect 6637 37632 6746 37637
rect 6637 37576 6642 37632
rect 6698 37576 6746 37632
rect 6637 37574 6746 37576
rect 24393 37634 24459 37637
rect 25840 37634 26000 37664
rect 24393 37632 26000 37634
rect 24393 37576 24398 37632
rect 24454 37576 26000 37632
rect 24393 37574 26000 37576
rect 0 37544 160 37574
rect 6637 37571 6703 37574
rect 24393 37571 24459 37574
rect 3913 37568 4229 37569
rect 3913 37504 3919 37568
rect 3983 37504 3999 37568
rect 4063 37504 4079 37568
rect 4143 37504 4159 37568
rect 4223 37504 4229 37568
rect 3913 37503 4229 37504
rect 9847 37568 10163 37569
rect 9847 37504 9853 37568
rect 9917 37504 9933 37568
rect 9997 37504 10013 37568
rect 10077 37504 10093 37568
rect 10157 37504 10163 37568
rect 9847 37503 10163 37504
rect 15781 37568 16097 37569
rect 15781 37504 15787 37568
rect 15851 37504 15867 37568
rect 15931 37504 15947 37568
rect 16011 37504 16027 37568
rect 16091 37504 16097 37568
rect 15781 37503 16097 37504
rect 21715 37568 22031 37569
rect 21715 37504 21721 37568
rect 21785 37504 21801 37568
rect 21865 37504 21881 37568
rect 21945 37504 21961 37568
rect 22025 37504 22031 37568
rect 25840 37544 26000 37574
rect 21715 37503 22031 37504
rect 3182 37436 3188 37500
rect 3252 37498 3258 37500
rect 3417 37498 3483 37501
rect 5349 37498 5415 37501
rect 3252 37496 3483 37498
rect 3252 37440 3422 37496
rect 3478 37440 3483 37496
rect 3252 37438 3483 37440
rect 3252 37436 3258 37438
rect 3417 37435 3483 37438
rect 4478 37496 5415 37498
rect 4478 37440 5354 37496
rect 5410 37440 5415 37496
rect 4478 37438 5415 37440
rect 0 37362 160 37392
rect 4478 37362 4538 37438
rect 5349 37435 5415 37438
rect 0 37302 4538 37362
rect 5533 37362 5599 37365
rect 5942 37362 5948 37364
rect 5533 37360 5948 37362
rect 5533 37304 5538 37360
rect 5594 37304 5948 37360
rect 5533 37302 5948 37304
rect 0 37272 160 37302
rect 5533 37299 5599 37302
rect 5942 37300 5948 37302
rect 6012 37300 6018 37364
rect 2773 37226 2839 37229
rect 12249 37226 12315 37229
rect 2773 37224 12315 37226
rect 2773 37168 2778 37224
rect 2834 37168 12254 37224
rect 12310 37168 12315 37224
rect 2773 37166 12315 37168
rect 2773 37163 2839 37166
rect 12249 37163 12315 37166
rect 24117 37226 24183 37229
rect 24117 37224 25146 37226
rect 24117 37168 24122 37224
rect 24178 37168 25146 37224
rect 24117 37166 25146 37168
rect 24117 37163 24183 37166
rect 0 37090 160 37120
rect 3877 37090 3943 37093
rect 0 37088 3943 37090
rect 0 37032 3882 37088
rect 3938 37032 3943 37088
rect 0 37030 3943 37032
rect 0 37000 160 37030
rect 3877 37027 3943 37030
rect 5390 37028 5396 37092
rect 5460 37090 5466 37092
rect 6545 37090 6611 37093
rect 5460 37088 6611 37090
rect 5460 37032 6550 37088
rect 6606 37032 6611 37088
rect 5460 37030 6611 37032
rect 25086 37090 25146 37166
rect 25840 37090 26000 37120
rect 25086 37030 26000 37090
rect 5460 37028 5466 37030
rect 3141 36954 3207 36957
rect 5398 36954 5458 37028
rect 6545 37027 6611 37030
rect 6880 37024 7196 37025
rect 6880 36960 6886 37024
rect 6950 36960 6966 37024
rect 7030 36960 7046 37024
rect 7110 36960 7126 37024
rect 7190 36960 7196 37024
rect 6880 36959 7196 36960
rect 12814 37024 13130 37025
rect 12814 36960 12820 37024
rect 12884 36960 12900 37024
rect 12964 36960 12980 37024
rect 13044 36960 13060 37024
rect 13124 36960 13130 37024
rect 12814 36959 13130 36960
rect 18748 37024 19064 37025
rect 18748 36960 18754 37024
rect 18818 36960 18834 37024
rect 18898 36960 18914 37024
rect 18978 36960 18994 37024
rect 19058 36960 19064 37024
rect 18748 36959 19064 36960
rect 24682 37024 24998 37025
rect 24682 36960 24688 37024
rect 24752 36960 24768 37024
rect 24832 36960 24848 37024
rect 24912 36960 24928 37024
rect 24992 36960 24998 37024
rect 25840 37000 26000 37030
rect 24682 36959 24998 36960
rect 3141 36952 5458 36954
rect 3141 36896 3146 36952
rect 3202 36896 5458 36952
rect 3141 36894 5458 36896
rect 7649 36954 7715 36957
rect 12065 36954 12131 36957
rect 7649 36952 12131 36954
rect 7649 36896 7654 36952
rect 7710 36896 12070 36952
rect 12126 36896 12131 36952
rect 7649 36894 12131 36896
rect 3141 36891 3207 36894
rect 7649 36891 7715 36894
rect 12065 36891 12131 36894
rect 0 36818 160 36848
rect 3233 36818 3299 36821
rect 0 36816 3299 36818
rect 0 36760 3238 36816
rect 3294 36760 3299 36816
rect 0 36758 3299 36760
rect 0 36728 160 36758
rect 3233 36755 3299 36758
rect 5257 36818 5323 36821
rect 8518 36818 8524 36820
rect 5257 36816 8524 36818
rect 5257 36760 5262 36816
rect 5318 36760 8524 36816
rect 5257 36758 8524 36760
rect 5257 36755 5323 36758
rect 8518 36756 8524 36758
rect 8588 36818 8594 36820
rect 9121 36818 9187 36821
rect 8588 36816 9187 36818
rect 8588 36760 9126 36816
rect 9182 36760 9187 36816
rect 8588 36758 9187 36760
rect 8588 36756 8594 36758
rect 9121 36755 9187 36758
rect 3233 36682 3299 36685
rect 4061 36682 4127 36685
rect 7649 36682 7715 36685
rect 3233 36680 7715 36682
rect 3233 36624 3238 36680
rect 3294 36624 4066 36680
rect 4122 36624 7654 36680
rect 7710 36624 7715 36680
rect 3233 36622 7715 36624
rect 3233 36619 3299 36622
rect 4061 36619 4127 36622
rect 7649 36619 7715 36622
rect 0 36546 160 36576
rect 1025 36546 1091 36549
rect 0 36544 1091 36546
rect 0 36488 1030 36544
rect 1086 36488 1091 36544
rect 0 36486 1091 36488
rect 0 36456 160 36486
rect 1025 36483 1091 36486
rect 6085 36546 6151 36549
rect 8334 36546 8340 36548
rect 6085 36544 8340 36546
rect 6085 36488 6090 36544
rect 6146 36488 8340 36544
rect 6085 36486 8340 36488
rect 6085 36483 6151 36486
rect 8334 36484 8340 36486
rect 8404 36484 8410 36548
rect 24393 36546 24459 36549
rect 25840 36546 26000 36576
rect 24393 36544 26000 36546
rect 24393 36488 24398 36544
rect 24454 36488 26000 36544
rect 24393 36486 26000 36488
rect 24393 36483 24459 36486
rect 3913 36480 4229 36481
rect 3913 36416 3919 36480
rect 3983 36416 3999 36480
rect 4063 36416 4079 36480
rect 4143 36416 4159 36480
rect 4223 36416 4229 36480
rect 3913 36415 4229 36416
rect 9847 36480 10163 36481
rect 9847 36416 9853 36480
rect 9917 36416 9933 36480
rect 9997 36416 10013 36480
rect 10077 36416 10093 36480
rect 10157 36416 10163 36480
rect 9847 36415 10163 36416
rect 15781 36480 16097 36481
rect 15781 36416 15787 36480
rect 15851 36416 15867 36480
rect 15931 36416 15947 36480
rect 16011 36416 16027 36480
rect 16091 36416 16097 36480
rect 15781 36415 16097 36416
rect 21715 36480 22031 36481
rect 21715 36416 21721 36480
rect 21785 36416 21801 36480
rect 21865 36416 21881 36480
rect 21945 36416 21961 36480
rect 22025 36416 22031 36480
rect 25840 36456 26000 36486
rect 21715 36415 22031 36416
rect 0 36274 160 36304
rect 1301 36274 1367 36277
rect 0 36272 1367 36274
rect 0 36216 1306 36272
rect 1362 36216 1367 36272
rect 0 36214 1367 36216
rect 0 36184 160 36214
rect 1301 36211 1367 36214
rect 3233 36274 3299 36277
rect 5022 36274 5028 36276
rect 3233 36272 5028 36274
rect 3233 36216 3238 36272
rect 3294 36216 5028 36272
rect 3233 36214 5028 36216
rect 3233 36211 3299 36214
rect 5022 36212 5028 36214
rect 5092 36274 5098 36276
rect 9397 36274 9463 36277
rect 5092 36272 9463 36274
rect 5092 36216 9402 36272
rect 9458 36216 9463 36272
rect 5092 36214 9463 36216
rect 5092 36212 5098 36214
rect 9397 36211 9463 36214
rect 10593 36274 10659 36277
rect 11237 36276 11303 36277
rect 11237 36274 11284 36276
rect 10593 36272 11284 36274
rect 10593 36216 10598 36272
rect 10654 36216 11242 36272
rect 10593 36214 11284 36216
rect 10593 36211 10659 36214
rect 11237 36212 11284 36214
rect 11348 36212 11354 36276
rect 11237 36211 11303 36212
rect 5441 36138 5507 36141
rect 14273 36138 14339 36141
rect 5441 36136 14339 36138
rect 5441 36080 5446 36136
rect 5502 36080 14278 36136
rect 14334 36080 14339 36136
rect 5441 36078 14339 36080
rect 5441 36075 5507 36078
rect 14273 36075 14339 36078
rect 0 36002 160 36032
rect 3417 36002 3483 36005
rect 0 36000 3483 36002
rect 0 35944 3422 36000
rect 3478 35944 3483 36000
rect 0 35942 3483 35944
rect 0 35912 160 35942
rect 3417 35939 3483 35942
rect 4061 36002 4127 36005
rect 5349 36002 5415 36005
rect 4061 36000 5415 36002
rect 4061 35944 4066 36000
rect 4122 35944 5354 36000
rect 5410 35944 5415 36000
rect 4061 35942 5415 35944
rect 4061 35939 4127 35942
rect 5349 35939 5415 35942
rect 22737 36002 22803 36005
rect 22870 36002 22876 36004
rect 22737 36000 22876 36002
rect 22737 35944 22742 36000
rect 22798 35944 22876 36000
rect 22737 35942 22876 35944
rect 22737 35939 22803 35942
rect 22870 35940 22876 35942
rect 22940 35940 22946 36004
rect 25129 36002 25195 36005
rect 25840 36002 26000 36032
rect 25129 36000 26000 36002
rect 25129 35944 25134 36000
rect 25190 35944 26000 36000
rect 25129 35942 26000 35944
rect 25129 35939 25195 35942
rect 6880 35936 7196 35937
rect 6880 35872 6886 35936
rect 6950 35872 6966 35936
rect 7030 35872 7046 35936
rect 7110 35872 7126 35936
rect 7190 35872 7196 35936
rect 6880 35871 7196 35872
rect 12814 35936 13130 35937
rect 12814 35872 12820 35936
rect 12884 35872 12900 35936
rect 12964 35872 12980 35936
rect 13044 35872 13060 35936
rect 13124 35872 13130 35936
rect 12814 35871 13130 35872
rect 18748 35936 19064 35937
rect 18748 35872 18754 35936
rect 18818 35872 18834 35936
rect 18898 35872 18914 35936
rect 18978 35872 18994 35936
rect 19058 35872 19064 35936
rect 18748 35871 19064 35872
rect 24682 35936 24998 35937
rect 24682 35872 24688 35936
rect 24752 35872 24768 35936
rect 24832 35872 24848 35936
rect 24912 35872 24928 35936
rect 24992 35872 24998 35936
rect 25840 35912 26000 35942
rect 24682 35871 24998 35872
rect 1025 35866 1091 35869
rect 2957 35866 3023 35869
rect 1025 35864 3023 35866
rect 1025 35808 1030 35864
rect 1086 35808 2962 35864
rect 3018 35808 3023 35864
rect 1025 35806 3023 35808
rect 1025 35803 1091 35806
rect 2957 35803 3023 35806
rect 3693 35866 3759 35869
rect 4286 35866 4292 35868
rect 3693 35864 4292 35866
rect 3693 35808 3698 35864
rect 3754 35808 4292 35864
rect 3693 35806 4292 35808
rect 3693 35803 3759 35806
rect 4286 35804 4292 35806
rect 4356 35804 4362 35868
rect 11513 35866 11579 35869
rect 12433 35866 12499 35869
rect 18321 35868 18387 35869
rect 18270 35866 18276 35868
rect 11513 35864 12499 35866
rect 11513 35808 11518 35864
rect 11574 35808 12438 35864
rect 12494 35808 12499 35864
rect 11513 35806 12499 35808
rect 18230 35806 18276 35866
rect 18340 35864 18387 35868
rect 18382 35808 18387 35864
rect 11513 35803 11579 35806
rect 12433 35803 12499 35806
rect 18270 35804 18276 35806
rect 18340 35804 18387 35808
rect 18321 35803 18387 35804
rect 0 35730 160 35760
rect 2865 35730 2931 35733
rect 0 35728 2931 35730
rect 0 35672 2870 35728
rect 2926 35672 2931 35728
rect 0 35670 2931 35672
rect 0 35640 160 35670
rect 2865 35667 2931 35670
rect 9397 35730 9463 35733
rect 10317 35730 10383 35733
rect 20989 35730 21055 35733
rect 9397 35728 21055 35730
rect 9397 35672 9402 35728
rect 9458 35672 10322 35728
rect 10378 35672 20994 35728
rect 21050 35672 21055 35728
rect 9397 35670 21055 35672
rect 9397 35667 9463 35670
rect 10317 35667 10383 35670
rect 20989 35667 21055 35670
rect 2037 35594 2103 35597
rect 4521 35594 4587 35597
rect 2037 35592 4587 35594
rect 2037 35536 2042 35592
rect 2098 35536 4526 35592
rect 4582 35536 4587 35592
rect 2037 35534 4587 35536
rect 2037 35531 2103 35534
rect 4521 35531 4587 35534
rect 5942 35532 5948 35596
rect 6012 35594 6018 35596
rect 8845 35594 8911 35597
rect 6012 35592 8911 35594
rect 6012 35536 8850 35592
rect 8906 35536 8911 35592
rect 6012 35534 8911 35536
rect 6012 35532 6018 35534
rect 8845 35531 8911 35534
rect 12985 35594 13051 35597
rect 22318 35594 22324 35596
rect 12985 35592 22324 35594
rect 12985 35536 12990 35592
rect 13046 35536 22324 35592
rect 12985 35534 22324 35536
rect 12985 35531 13051 35534
rect 22318 35532 22324 35534
rect 22388 35532 22394 35596
rect 0 35458 160 35488
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35368 160 35398
rect 1577 35395 1643 35398
rect 13445 35460 13511 35461
rect 13445 35456 13492 35460
rect 13556 35458 13562 35460
rect 24393 35458 24459 35461
rect 25840 35458 26000 35488
rect 13445 35400 13450 35456
rect 13445 35396 13492 35400
rect 13556 35398 13602 35458
rect 24393 35456 26000 35458
rect 24393 35400 24398 35456
rect 24454 35400 26000 35456
rect 24393 35398 26000 35400
rect 13556 35396 13562 35398
rect 13445 35395 13511 35396
rect 24393 35395 24459 35398
rect 3913 35392 4229 35393
rect 3913 35328 3919 35392
rect 3983 35328 3999 35392
rect 4063 35328 4079 35392
rect 4143 35328 4159 35392
rect 4223 35328 4229 35392
rect 3913 35327 4229 35328
rect 9847 35392 10163 35393
rect 9847 35328 9853 35392
rect 9917 35328 9933 35392
rect 9997 35328 10013 35392
rect 10077 35328 10093 35392
rect 10157 35328 10163 35392
rect 9847 35327 10163 35328
rect 15781 35392 16097 35393
rect 15781 35328 15787 35392
rect 15851 35328 15867 35392
rect 15931 35328 15947 35392
rect 16011 35328 16027 35392
rect 16091 35328 16097 35392
rect 15781 35327 16097 35328
rect 21715 35392 22031 35393
rect 21715 35328 21721 35392
rect 21785 35328 21801 35392
rect 21865 35328 21881 35392
rect 21945 35328 21961 35392
rect 22025 35328 22031 35392
rect 25840 35368 26000 35398
rect 21715 35327 22031 35328
rect 0 35186 160 35216
rect 3785 35186 3851 35189
rect 0 35184 3851 35186
rect 0 35128 3790 35184
rect 3846 35128 3851 35184
rect 0 35126 3851 35128
rect 0 35096 160 35126
rect 3785 35123 3851 35126
rect 8937 35186 9003 35189
rect 13353 35186 13419 35189
rect 8937 35184 13419 35186
rect 8937 35128 8942 35184
rect 8998 35128 13358 35184
rect 13414 35128 13419 35184
rect 8937 35126 13419 35128
rect 8937 35123 9003 35126
rect 13353 35123 13419 35126
rect 1393 35048 1459 35053
rect 12065 35052 12131 35053
rect 12014 35050 12020 35052
rect 1393 34992 1398 35048
rect 1454 34992 1459 35048
rect 1393 34987 1459 34992
rect 11938 34990 12020 35050
rect 12084 35050 12131 35052
rect 21265 35050 21331 35053
rect 12084 35048 21331 35050
rect 12126 34992 21270 35048
rect 21326 34992 21331 35048
rect 12014 34988 12020 34990
rect 12084 34990 21331 34992
rect 12084 34988 12131 34990
rect 12065 34987 12131 34988
rect 21265 34987 21331 34990
rect 0 34914 160 34944
rect 1396 34914 1456 34987
rect 0 34854 1456 34914
rect 25221 34914 25287 34917
rect 25840 34914 26000 34944
rect 25221 34912 26000 34914
rect 25221 34856 25226 34912
rect 25282 34856 26000 34912
rect 25221 34854 26000 34856
rect 0 34824 160 34854
rect 25221 34851 25287 34854
rect 6880 34848 7196 34849
rect 6880 34784 6886 34848
rect 6950 34784 6966 34848
rect 7030 34784 7046 34848
rect 7110 34784 7126 34848
rect 7190 34784 7196 34848
rect 6880 34783 7196 34784
rect 12814 34848 13130 34849
rect 12814 34784 12820 34848
rect 12884 34784 12900 34848
rect 12964 34784 12980 34848
rect 13044 34784 13060 34848
rect 13124 34784 13130 34848
rect 12814 34783 13130 34784
rect 18748 34848 19064 34849
rect 18748 34784 18754 34848
rect 18818 34784 18834 34848
rect 18898 34784 18914 34848
rect 18978 34784 18994 34848
rect 19058 34784 19064 34848
rect 18748 34783 19064 34784
rect 24682 34848 24998 34849
rect 24682 34784 24688 34848
rect 24752 34784 24768 34848
rect 24832 34784 24848 34848
rect 24912 34784 24928 34848
rect 24992 34784 24998 34848
rect 25840 34824 26000 34854
rect 24682 34783 24998 34784
rect 3325 34778 3391 34781
rect 4889 34778 4955 34781
rect 3325 34776 4955 34778
rect 3325 34720 3330 34776
rect 3386 34720 4894 34776
rect 4950 34720 4955 34776
rect 3325 34718 4955 34720
rect 3325 34715 3391 34718
rect 4889 34715 4955 34718
rect 13261 34778 13327 34781
rect 13261 34776 14842 34778
rect 13261 34720 13266 34776
rect 13322 34720 14842 34776
rect 13261 34718 14842 34720
rect 13261 34715 13327 34718
rect 0 34642 160 34672
rect 749 34642 815 34645
rect 0 34640 815 34642
rect 0 34584 754 34640
rect 810 34584 815 34640
rect 0 34582 815 34584
rect 0 34552 160 34582
rect 749 34579 815 34582
rect 1669 34642 1735 34645
rect 5165 34642 5231 34645
rect 1669 34640 5231 34642
rect 1669 34584 1674 34640
rect 1730 34584 5170 34640
rect 5226 34584 5231 34640
rect 1669 34582 5231 34584
rect 1669 34579 1735 34582
rect 5165 34579 5231 34582
rect 12198 34580 12204 34644
rect 12268 34642 12274 34644
rect 14549 34642 14615 34645
rect 12268 34640 14615 34642
rect 12268 34584 14554 34640
rect 14610 34584 14615 34640
rect 12268 34582 14615 34584
rect 14782 34642 14842 34718
rect 20713 34642 20779 34645
rect 14782 34640 20779 34642
rect 14782 34584 20718 34640
rect 20774 34584 20779 34640
rect 14782 34582 20779 34584
rect 12268 34580 12274 34582
rect 14549 34579 14615 34582
rect 20713 34579 20779 34582
rect 4061 34506 4127 34509
rect 2730 34504 4127 34506
rect 2730 34448 4066 34504
rect 4122 34448 4127 34504
rect 2730 34446 4127 34448
rect 0 34370 160 34400
rect 2730 34370 2790 34446
rect 4061 34443 4127 34446
rect 5349 34506 5415 34509
rect 13077 34506 13143 34509
rect 15009 34506 15075 34509
rect 18965 34506 19031 34509
rect 5349 34504 19031 34506
rect 5349 34448 5354 34504
rect 5410 34448 13082 34504
rect 13138 34448 15014 34504
rect 15070 34448 18970 34504
rect 19026 34448 19031 34504
rect 5349 34446 19031 34448
rect 5349 34443 5415 34446
rect 13077 34443 13143 34446
rect 15009 34443 15075 34446
rect 18965 34443 19031 34446
rect 24393 34506 24459 34509
rect 24393 34504 25146 34506
rect 24393 34448 24398 34504
rect 24454 34448 25146 34504
rect 24393 34446 25146 34448
rect 24393 34443 24459 34446
rect 0 34310 2790 34370
rect 25086 34370 25146 34446
rect 25840 34370 26000 34400
rect 25086 34310 26000 34370
rect 0 34280 160 34310
rect 3913 34304 4229 34305
rect 3913 34240 3919 34304
rect 3983 34240 3999 34304
rect 4063 34240 4079 34304
rect 4143 34240 4159 34304
rect 4223 34240 4229 34304
rect 3913 34239 4229 34240
rect 9847 34304 10163 34305
rect 9847 34240 9853 34304
rect 9917 34240 9933 34304
rect 9997 34240 10013 34304
rect 10077 34240 10093 34304
rect 10157 34240 10163 34304
rect 9847 34239 10163 34240
rect 15781 34304 16097 34305
rect 15781 34240 15787 34304
rect 15851 34240 15867 34304
rect 15931 34240 15947 34304
rect 16011 34240 16027 34304
rect 16091 34240 16097 34304
rect 15781 34239 16097 34240
rect 21715 34304 22031 34305
rect 21715 34240 21721 34304
rect 21785 34240 21801 34304
rect 21865 34240 21881 34304
rect 21945 34240 21961 34304
rect 22025 34240 22031 34304
rect 25840 34280 26000 34310
rect 21715 34239 22031 34240
rect 6177 34234 6243 34237
rect 8845 34234 8911 34237
rect 6177 34232 8911 34234
rect 6177 34176 6182 34232
rect 6238 34176 8850 34232
rect 8906 34176 8911 34232
rect 6177 34174 8911 34176
rect 6177 34171 6243 34174
rect 8845 34171 8911 34174
rect 9029 34234 9095 34237
rect 9489 34234 9555 34237
rect 9029 34232 9555 34234
rect 9029 34176 9034 34232
rect 9090 34176 9494 34232
rect 9550 34176 9555 34232
rect 9029 34174 9555 34176
rect 9029 34171 9095 34174
rect 9489 34171 9555 34174
rect 10777 34232 10843 34237
rect 10777 34176 10782 34232
rect 10838 34176 10843 34232
rect 10777 34171 10843 34176
rect 0 34098 160 34128
rect 3417 34098 3483 34101
rect 0 34096 3483 34098
rect 0 34040 3422 34096
rect 3478 34040 3483 34096
rect 0 34038 3483 34040
rect 0 34008 160 34038
rect 3417 34035 3483 34038
rect 6821 34098 6887 34101
rect 10542 34098 10548 34100
rect 6821 34096 10548 34098
rect 6821 34040 6826 34096
rect 6882 34040 10548 34096
rect 6821 34038 10548 34040
rect 6821 34035 6887 34038
rect 10542 34036 10548 34038
rect 10612 34098 10618 34100
rect 10780 34098 10840 34171
rect 10612 34038 10840 34098
rect 12525 34098 12591 34101
rect 17769 34098 17835 34101
rect 12525 34096 17835 34098
rect 12525 34040 12530 34096
rect 12586 34040 17774 34096
rect 17830 34040 17835 34096
rect 12525 34038 17835 34040
rect 10612 34036 10618 34038
rect 12525 34035 12591 34038
rect 17769 34035 17835 34038
rect 4061 33962 4127 33965
rect 8845 33962 8911 33965
rect 9397 33962 9463 33965
rect 4061 33960 9463 33962
rect 4061 33904 4066 33960
rect 4122 33904 8850 33960
rect 8906 33904 9402 33960
rect 9458 33904 9463 33960
rect 4061 33902 9463 33904
rect 4061 33899 4127 33902
rect 8845 33899 8911 33902
rect 9397 33899 9463 33902
rect 12341 33962 12407 33965
rect 12525 33962 12591 33965
rect 12341 33960 12591 33962
rect 12341 33904 12346 33960
rect 12402 33904 12530 33960
rect 12586 33904 12591 33960
rect 12341 33902 12591 33904
rect 12341 33899 12407 33902
rect 12525 33899 12591 33902
rect 13905 33962 13971 33965
rect 17033 33962 17099 33965
rect 13905 33960 17099 33962
rect 13905 33904 13910 33960
rect 13966 33904 17038 33960
rect 17094 33904 17099 33960
rect 13905 33902 17099 33904
rect 13905 33899 13971 33902
rect 17033 33899 17099 33902
rect 0 33826 160 33856
rect 1025 33826 1091 33829
rect 0 33824 1091 33826
rect 0 33768 1030 33824
rect 1086 33768 1091 33824
rect 0 33766 1091 33768
rect 0 33736 160 33766
rect 1025 33763 1091 33766
rect 25221 33826 25287 33829
rect 25840 33826 26000 33856
rect 25221 33824 26000 33826
rect 25221 33768 25226 33824
rect 25282 33768 26000 33824
rect 25221 33766 26000 33768
rect 25221 33763 25287 33766
rect 6880 33760 7196 33761
rect 6880 33696 6886 33760
rect 6950 33696 6966 33760
rect 7030 33696 7046 33760
rect 7110 33696 7126 33760
rect 7190 33696 7196 33760
rect 6880 33695 7196 33696
rect 12814 33760 13130 33761
rect 12814 33696 12820 33760
rect 12884 33696 12900 33760
rect 12964 33696 12980 33760
rect 13044 33696 13060 33760
rect 13124 33696 13130 33760
rect 12814 33695 13130 33696
rect 18748 33760 19064 33761
rect 18748 33696 18754 33760
rect 18818 33696 18834 33760
rect 18898 33696 18914 33760
rect 18978 33696 18994 33760
rect 19058 33696 19064 33760
rect 18748 33695 19064 33696
rect 24682 33760 24998 33761
rect 24682 33696 24688 33760
rect 24752 33696 24768 33760
rect 24832 33696 24848 33760
rect 24912 33696 24928 33760
rect 24992 33696 24998 33760
rect 25840 33736 26000 33766
rect 24682 33695 24998 33696
rect 2221 33690 2287 33693
rect 2221 33688 2790 33690
rect 2221 33632 2226 33688
rect 2282 33632 2790 33688
rect 2221 33630 2790 33632
rect 2221 33627 2287 33630
rect 0 33554 160 33584
rect 1301 33554 1367 33557
rect 0 33552 1367 33554
rect 0 33496 1306 33552
rect 1362 33496 1367 33552
rect 0 33494 1367 33496
rect 2730 33554 2790 33630
rect 7465 33554 7531 33557
rect 2730 33552 7531 33554
rect 2730 33496 7470 33552
rect 7526 33496 7531 33552
rect 2730 33494 7531 33496
rect 0 33464 160 33494
rect 1301 33491 1367 33494
rect 7465 33491 7531 33494
rect 7833 33554 7899 33557
rect 9765 33554 9831 33557
rect 7833 33552 9831 33554
rect 7833 33496 7838 33552
rect 7894 33496 9770 33552
rect 9826 33496 9831 33552
rect 7833 33494 9831 33496
rect 7833 33491 7899 33494
rect 9765 33491 9831 33494
rect 18965 33554 19031 33557
rect 22737 33554 22803 33557
rect 18965 33552 22803 33554
rect 18965 33496 18970 33552
rect 19026 33496 22742 33552
rect 22798 33496 22803 33552
rect 18965 33494 22803 33496
rect 18965 33491 19031 33494
rect 22737 33491 22803 33494
rect 4337 33418 4403 33421
rect 19333 33418 19399 33421
rect 4337 33416 19399 33418
rect 4337 33360 4342 33416
rect 4398 33360 19338 33416
rect 19394 33360 19399 33416
rect 4337 33358 19399 33360
rect 4337 33355 4403 33358
rect 19333 33355 19399 33358
rect 0 33282 160 33312
rect 2865 33282 2931 33285
rect 0 33280 2931 33282
rect 0 33224 2870 33280
rect 2926 33224 2931 33280
rect 0 33222 2931 33224
rect 0 33192 160 33222
rect 2865 33219 2931 33222
rect 17953 33282 18019 33285
rect 18413 33282 18479 33285
rect 17953 33280 18479 33282
rect 17953 33224 17958 33280
rect 18014 33224 18418 33280
rect 18474 33224 18479 33280
rect 17953 33222 18479 33224
rect 17953 33219 18019 33222
rect 18413 33219 18479 33222
rect 22553 33282 22619 33285
rect 22686 33282 22692 33284
rect 22553 33280 22692 33282
rect 22553 33224 22558 33280
rect 22614 33224 22692 33280
rect 22553 33222 22692 33224
rect 22553 33219 22619 33222
rect 22686 33220 22692 33222
rect 22756 33220 22762 33284
rect 24393 33282 24459 33285
rect 25840 33282 26000 33312
rect 24393 33280 26000 33282
rect 24393 33224 24398 33280
rect 24454 33224 26000 33280
rect 24393 33222 26000 33224
rect 24393 33219 24459 33222
rect 3913 33216 4229 33217
rect 3913 33152 3919 33216
rect 3983 33152 3999 33216
rect 4063 33152 4079 33216
rect 4143 33152 4159 33216
rect 4223 33152 4229 33216
rect 3913 33151 4229 33152
rect 9847 33216 10163 33217
rect 9847 33152 9853 33216
rect 9917 33152 9933 33216
rect 9997 33152 10013 33216
rect 10077 33152 10093 33216
rect 10157 33152 10163 33216
rect 9847 33151 10163 33152
rect 15781 33216 16097 33217
rect 15781 33152 15787 33216
rect 15851 33152 15867 33216
rect 15931 33152 15947 33216
rect 16011 33152 16027 33216
rect 16091 33152 16097 33216
rect 15781 33151 16097 33152
rect 21715 33216 22031 33217
rect 21715 33152 21721 33216
rect 21785 33152 21801 33216
rect 21865 33152 21881 33216
rect 21945 33152 21961 33216
rect 22025 33152 22031 33216
rect 25840 33192 26000 33222
rect 21715 33151 22031 33152
rect 18086 33084 18092 33148
rect 18156 33146 18162 33148
rect 19701 33146 19767 33149
rect 18156 33144 19767 33146
rect 18156 33088 19706 33144
rect 19762 33088 19767 33144
rect 18156 33086 19767 33088
rect 18156 33084 18162 33086
rect 19701 33083 19767 33086
rect 0 33010 160 33040
rect 1485 33010 1551 33013
rect 0 33008 1551 33010
rect 0 32952 1490 33008
rect 1546 32952 1551 33008
rect 0 32950 1551 32952
rect 0 32920 160 32950
rect 1485 32947 1551 32950
rect 3049 33010 3115 33013
rect 5257 33010 5323 33013
rect 3049 33008 5323 33010
rect 3049 32952 3054 33008
rect 3110 32952 5262 33008
rect 5318 32952 5323 33008
rect 3049 32950 5323 32952
rect 3049 32947 3115 32950
rect 5257 32947 5323 32950
rect 6361 33010 6427 33013
rect 11646 33010 11652 33012
rect 6361 33008 11652 33010
rect 6361 32952 6366 33008
rect 6422 32952 11652 33008
rect 6361 32950 11652 32952
rect 6361 32947 6427 32950
rect 11646 32948 11652 32950
rect 11716 32948 11722 33012
rect 2037 32874 2103 32877
rect 6913 32874 6979 32877
rect 2037 32872 6979 32874
rect 2037 32816 2042 32872
rect 2098 32816 6918 32872
rect 6974 32816 6979 32872
rect 2037 32814 6979 32816
rect 2037 32811 2103 32814
rect 6913 32811 6979 32814
rect 7649 32874 7715 32877
rect 13537 32874 13603 32877
rect 15377 32874 15443 32877
rect 7649 32872 15443 32874
rect 7649 32816 7654 32872
rect 7710 32816 13542 32872
rect 13598 32816 15382 32872
rect 15438 32816 15443 32872
rect 7649 32814 15443 32816
rect 7649 32811 7715 32814
rect 13537 32811 13603 32814
rect 15377 32811 15443 32814
rect 0 32738 160 32768
rect 2773 32738 2839 32741
rect 0 32736 2839 32738
rect 0 32680 2778 32736
rect 2834 32680 2839 32736
rect 0 32678 2839 32680
rect 0 32648 160 32678
rect 2773 32675 2839 32678
rect 4521 32738 4587 32741
rect 4654 32738 4660 32740
rect 4521 32736 4660 32738
rect 4521 32680 4526 32736
rect 4582 32680 4660 32736
rect 4521 32678 4660 32680
rect 4521 32675 4587 32678
rect 4654 32676 4660 32678
rect 4724 32676 4730 32740
rect 7281 32738 7347 32741
rect 11237 32740 11303 32741
rect 11237 32738 11284 32740
rect 7281 32736 11284 32738
rect 11348 32738 11354 32740
rect 25221 32738 25287 32741
rect 25840 32738 26000 32768
rect 7281 32680 7286 32736
rect 7342 32680 11242 32736
rect 7281 32678 11284 32680
rect 7281 32675 7347 32678
rect 11237 32676 11284 32678
rect 11348 32678 11430 32738
rect 25221 32736 26000 32738
rect 25221 32680 25226 32736
rect 25282 32680 26000 32736
rect 25221 32678 26000 32680
rect 11348 32676 11354 32678
rect 11237 32675 11303 32676
rect 25221 32675 25287 32678
rect 6880 32672 7196 32673
rect 6880 32608 6886 32672
rect 6950 32608 6966 32672
rect 7030 32608 7046 32672
rect 7110 32608 7126 32672
rect 7190 32608 7196 32672
rect 6880 32607 7196 32608
rect 12814 32672 13130 32673
rect 12814 32608 12820 32672
rect 12884 32608 12900 32672
rect 12964 32608 12980 32672
rect 13044 32608 13060 32672
rect 13124 32608 13130 32672
rect 12814 32607 13130 32608
rect 18748 32672 19064 32673
rect 18748 32608 18754 32672
rect 18818 32608 18834 32672
rect 18898 32608 18914 32672
rect 18978 32608 18994 32672
rect 19058 32608 19064 32672
rect 18748 32607 19064 32608
rect 24682 32672 24998 32673
rect 24682 32608 24688 32672
rect 24752 32608 24768 32672
rect 24832 32608 24848 32672
rect 24912 32608 24928 32672
rect 24992 32608 24998 32672
rect 25840 32648 26000 32678
rect 24682 32607 24998 32608
rect 2630 32540 2636 32604
rect 2700 32602 2706 32604
rect 3601 32602 3667 32605
rect 2700 32600 3667 32602
rect 2700 32544 3606 32600
rect 3662 32544 3667 32600
rect 2700 32542 3667 32544
rect 2700 32540 2706 32542
rect 3601 32539 3667 32542
rect 8569 32602 8635 32605
rect 9489 32602 9555 32605
rect 8569 32600 9555 32602
rect 8569 32544 8574 32600
rect 8630 32544 9494 32600
rect 9550 32544 9555 32600
rect 8569 32542 9555 32544
rect 8569 32539 8635 32542
rect 9489 32539 9555 32542
rect 0 32466 160 32496
rect 1301 32466 1367 32469
rect 0 32464 1367 32466
rect 0 32408 1306 32464
rect 1362 32408 1367 32464
rect 0 32406 1367 32408
rect 0 32376 160 32406
rect 1301 32403 1367 32406
rect 2405 32466 2471 32469
rect 3182 32466 3188 32468
rect 2405 32464 3188 32466
rect 2405 32408 2410 32464
rect 2466 32408 3188 32464
rect 2405 32406 3188 32408
rect 2405 32403 2471 32406
rect 3182 32404 3188 32406
rect 3252 32404 3258 32468
rect 3550 32268 3556 32332
rect 3620 32330 3626 32332
rect 4061 32330 4127 32333
rect 3620 32328 4127 32330
rect 3620 32272 4066 32328
rect 4122 32272 4127 32328
rect 3620 32270 4127 32272
rect 3620 32268 3626 32270
rect 4061 32267 4127 32270
rect 5625 32330 5691 32333
rect 11830 32330 11836 32332
rect 5625 32328 11836 32330
rect 5625 32272 5630 32328
rect 5686 32272 11836 32328
rect 5625 32270 11836 32272
rect 5625 32267 5691 32270
rect 11830 32268 11836 32270
rect 11900 32268 11906 32332
rect 0 32194 160 32224
rect 1209 32194 1275 32197
rect 0 32192 1275 32194
rect 0 32136 1214 32192
rect 1270 32136 1275 32192
rect 0 32134 1275 32136
rect 0 32104 160 32134
rect 1209 32131 1275 32134
rect 24393 32194 24459 32197
rect 25840 32194 26000 32224
rect 24393 32192 26000 32194
rect 24393 32136 24398 32192
rect 24454 32136 26000 32192
rect 24393 32134 26000 32136
rect 24393 32131 24459 32134
rect 3913 32128 4229 32129
rect 3913 32064 3919 32128
rect 3983 32064 3999 32128
rect 4063 32064 4079 32128
rect 4143 32064 4159 32128
rect 4223 32064 4229 32128
rect 3913 32063 4229 32064
rect 9847 32128 10163 32129
rect 9847 32064 9853 32128
rect 9917 32064 9933 32128
rect 9997 32064 10013 32128
rect 10077 32064 10093 32128
rect 10157 32064 10163 32128
rect 9847 32063 10163 32064
rect 15781 32128 16097 32129
rect 15781 32064 15787 32128
rect 15851 32064 15867 32128
rect 15931 32064 15947 32128
rect 16011 32064 16027 32128
rect 16091 32064 16097 32128
rect 15781 32063 16097 32064
rect 21715 32128 22031 32129
rect 21715 32064 21721 32128
rect 21785 32064 21801 32128
rect 21865 32064 21881 32128
rect 21945 32064 21961 32128
rect 22025 32064 22031 32128
rect 25840 32104 26000 32134
rect 21715 32063 22031 32064
rect 0 31922 160 31952
rect 3325 31922 3391 31925
rect 0 31920 3391 31922
rect 0 31864 3330 31920
rect 3386 31864 3391 31920
rect 0 31862 3391 31864
rect 0 31832 160 31862
rect 3325 31859 3391 31862
rect 4286 31860 4292 31924
rect 4356 31922 4362 31924
rect 5390 31922 5396 31924
rect 4356 31862 5396 31922
rect 4356 31860 4362 31862
rect 5390 31860 5396 31862
rect 5460 31922 5466 31924
rect 9673 31922 9739 31925
rect 5460 31920 9739 31922
rect 5460 31864 9678 31920
rect 9734 31864 9739 31920
rect 5460 31862 9739 31864
rect 5460 31860 5466 31862
rect 9673 31859 9739 31862
rect 2129 31786 2195 31789
rect 8477 31786 8543 31789
rect 16021 31786 16087 31789
rect 23197 31788 23263 31789
rect 23197 31786 23244 31788
rect 2129 31784 8402 31786
rect 2129 31728 2134 31784
rect 2190 31728 8402 31784
rect 2129 31726 8402 31728
rect 2129 31723 2195 31726
rect 0 31650 160 31680
rect 3785 31650 3851 31653
rect 6637 31650 6703 31653
rect 0 31648 3851 31650
rect 0 31592 3790 31648
rect 3846 31592 3851 31648
rect 0 31590 3851 31592
rect 0 31560 160 31590
rect 3785 31587 3851 31590
rect 3926 31648 6703 31650
rect 3926 31592 6642 31648
rect 6698 31592 6703 31648
rect 3926 31590 6703 31592
rect 8342 31650 8402 31726
rect 8477 31784 16087 31786
rect 8477 31728 8482 31784
rect 8538 31728 16026 31784
rect 16082 31728 16087 31784
rect 8477 31726 16087 31728
rect 23152 31784 23244 31786
rect 23152 31728 23202 31784
rect 23152 31726 23244 31728
rect 8477 31723 8543 31726
rect 16021 31723 16087 31726
rect 23197 31724 23244 31726
rect 23308 31724 23314 31788
rect 23197 31723 23263 31724
rect 8518 31650 8524 31652
rect 8342 31590 8524 31650
rect 2221 31514 2287 31517
rect 3926 31514 3986 31590
rect 6637 31587 6703 31590
rect 8518 31588 8524 31590
rect 8588 31588 8594 31652
rect 13905 31650 13971 31653
rect 15285 31650 15351 31653
rect 13905 31648 15351 31650
rect 13905 31592 13910 31648
rect 13966 31592 15290 31648
rect 15346 31592 15351 31648
rect 13905 31590 15351 31592
rect 13905 31587 13971 31590
rect 15285 31587 15351 31590
rect 25129 31650 25195 31653
rect 25840 31650 26000 31680
rect 25129 31648 26000 31650
rect 25129 31592 25134 31648
rect 25190 31592 26000 31648
rect 25129 31590 26000 31592
rect 25129 31587 25195 31590
rect 6880 31584 7196 31585
rect 6880 31520 6886 31584
rect 6950 31520 6966 31584
rect 7030 31520 7046 31584
rect 7110 31520 7126 31584
rect 7190 31520 7196 31584
rect 6880 31519 7196 31520
rect 12814 31584 13130 31585
rect 12814 31520 12820 31584
rect 12884 31520 12900 31584
rect 12964 31520 12980 31584
rect 13044 31520 13060 31584
rect 13124 31520 13130 31584
rect 12814 31519 13130 31520
rect 18748 31584 19064 31585
rect 18748 31520 18754 31584
rect 18818 31520 18834 31584
rect 18898 31520 18914 31584
rect 18978 31520 18994 31584
rect 19058 31520 19064 31584
rect 18748 31519 19064 31520
rect 24682 31584 24998 31585
rect 24682 31520 24688 31584
rect 24752 31520 24768 31584
rect 24832 31520 24848 31584
rect 24912 31520 24928 31584
rect 24992 31520 24998 31584
rect 25840 31560 26000 31590
rect 24682 31519 24998 31520
rect 2221 31512 3986 31514
rect 2221 31456 2226 31512
rect 2282 31456 3986 31512
rect 2221 31454 3986 31456
rect 4153 31514 4219 31517
rect 4613 31514 4679 31517
rect 6453 31514 6519 31517
rect 12617 31514 12683 31517
rect 4153 31512 6519 31514
rect 4153 31456 4158 31512
rect 4214 31456 4618 31512
rect 4674 31456 6458 31512
rect 6514 31456 6519 31512
rect 4153 31454 6519 31456
rect 2221 31451 2287 31454
rect 4153 31451 4219 31454
rect 4613 31451 4679 31454
rect 6453 31451 6519 31454
rect 12574 31512 12683 31514
rect 12574 31456 12622 31512
rect 12678 31456 12683 31512
rect 12574 31451 12683 31456
rect 0 31378 160 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 160 31318
rect 1393 31315 1459 31318
rect 4153 31378 4219 31381
rect 11145 31378 11211 31381
rect 4153 31376 11211 31378
rect 4153 31320 4158 31376
rect 4214 31320 11150 31376
rect 11206 31320 11211 31376
rect 4153 31318 11211 31320
rect 4153 31315 4219 31318
rect 11145 31315 11211 31318
rect 12574 31245 12634 31451
rect 4981 31242 5047 31245
rect 9765 31242 9831 31245
rect 4981 31240 12450 31242
rect 4981 31184 4986 31240
rect 5042 31184 9770 31240
rect 9826 31184 12450 31240
rect 4981 31182 12450 31184
rect 12574 31240 12683 31245
rect 12574 31184 12622 31240
rect 12678 31184 12683 31240
rect 12574 31182 12683 31184
rect 4981 31179 5047 31182
rect 9765 31179 9831 31182
rect 0 31106 160 31136
rect 2773 31106 2839 31109
rect 0 31104 2839 31106
rect 0 31048 2778 31104
rect 2834 31048 2839 31104
rect 0 31046 2839 31048
rect 0 31016 160 31046
rect 2773 31043 2839 31046
rect 10501 31106 10567 31109
rect 10501 31104 10978 31106
rect 10501 31048 10506 31104
rect 10562 31048 10978 31104
rect 10501 31046 10978 31048
rect 10501 31043 10567 31046
rect 3913 31040 4229 31041
rect 3913 30976 3919 31040
rect 3983 30976 3999 31040
rect 4063 30976 4079 31040
rect 4143 30976 4159 31040
rect 4223 30976 4229 31040
rect 3913 30975 4229 30976
rect 9847 31040 10163 31041
rect 9847 30976 9853 31040
rect 9917 30976 9933 31040
rect 9997 30976 10013 31040
rect 10077 30976 10093 31040
rect 10157 30976 10163 31040
rect 9847 30975 10163 30976
rect 0 30834 160 30864
rect 1301 30834 1367 30837
rect 0 30832 1367 30834
rect 0 30776 1306 30832
rect 1362 30776 1367 30832
rect 0 30774 1367 30776
rect 0 30744 160 30774
rect 1301 30771 1367 30774
rect 1894 30772 1900 30836
rect 1964 30834 1970 30836
rect 4889 30834 4955 30837
rect 10133 30834 10199 30837
rect 10777 30834 10843 30837
rect 1964 30832 4955 30834
rect 1964 30776 4894 30832
rect 4950 30776 4955 30832
rect 1964 30774 4955 30776
rect 1964 30772 1970 30774
rect 4889 30771 4955 30774
rect 8342 30832 10843 30834
rect 8342 30776 10138 30832
rect 10194 30776 10782 30832
rect 10838 30776 10843 30832
rect 8342 30774 10843 30776
rect 2589 30700 2655 30701
rect 2589 30698 2636 30700
rect 2508 30696 2636 30698
rect 2700 30698 2706 30700
rect 8342 30698 8402 30774
rect 10133 30771 10199 30774
rect 10777 30771 10843 30774
rect 10918 30701 10978 31046
rect 12390 30834 12450 31182
rect 12617 31179 12683 31182
rect 15377 31242 15443 31245
rect 15745 31242 15811 31245
rect 15377 31240 15811 31242
rect 15377 31184 15382 31240
rect 15438 31184 15750 31240
rect 15806 31184 15811 31240
rect 15377 31182 15811 31184
rect 15377 31179 15443 31182
rect 15745 31179 15811 31182
rect 13261 31106 13327 31109
rect 13486 31106 13492 31108
rect 13261 31104 13492 31106
rect 13261 31048 13266 31104
rect 13322 31048 13492 31104
rect 13261 31046 13492 31048
rect 13261 31043 13327 31046
rect 13486 31044 13492 31046
rect 13556 31044 13562 31108
rect 24393 31106 24459 31109
rect 25840 31106 26000 31136
rect 24393 31104 26000 31106
rect 24393 31048 24398 31104
rect 24454 31048 26000 31104
rect 24393 31046 26000 31048
rect 24393 31043 24459 31046
rect 15781 31040 16097 31041
rect 15781 30976 15787 31040
rect 15851 30976 15867 31040
rect 15931 30976 15947 31040
rect 16011 30976 16027 31040
rect 16091 30976 16097 31040
rect 15781 30975 16097 30976
rect 21715 31040 22031 31041
rect 21715 30976 21721 31040
rect 21785 30976 21801 31040
rect 21865 30976 21881 31040
rect 21945 30976 21961 31040
rect 22025 30976 22031 31040
rect 25840 31016 26000 31046
rect 21715 30975 22031 30976
rect 14222 30834 14228 30836
rect 12390 30774 14228 30834
rect 14222 30772 14228 30774
rect 14292 30772 14298 30836
rect 16982 30772 16988 30836
rect 17052 30834 17058 30836
rect 24577 30834 24643 30837
rect 17052 30832 24643 30834
rect 17052 30776 24582 30832
rect 24638 30776 24643 30832
rect 17052 30774 24643 30776
rect 17052 30772 17058 30774
rect 24577 30771 24643 30774
rect 9213 30700 9279 30701
rect 10593 30700 10659 30701
rect 2508 30640 2594 30696
rect 2508 30638 2636 30640
rect 2589 30636 2636 30638
rect 2700 30638 8402 30698
rect 2700 30636 2706 30638
rect 8518 30636 8524 30700
rect 8588 30698 8594 30700
rect 9213 30698 9260 30700
rect 8588 30696 9260 30698
rect 8588 30640 9218 30696
rect 8588 30638 9260 30640
rect 8588 30636 8594 30638
rect 9213 30636 9260 30638
rect 9324 30636 9330 30700
rect 9438 30636 9444 30700
rect 9508 30698 9514 30700
rect 10358 30698 10364 30700
rect 9508 30638 10364 30698
rect 9508 30636 9514 30638
rect 10358 30636 10364 30638
rect 10428 30636 10434 30700
rect 10542 30636 10548 30700
rect 10612 30698 10659 30700
rect 10612 30696 10704 30698
rect 10654 30640 10704 30696
rect 10612 30638 10704 30640
rect 10918 30696 11027 30701
rect 10918 30640 10966 30696
rect 11022 30640 11027 30696
rect 10918 30638 11027 30640
rect 10612 30636 10659 30638
rect 2589 30635 2655 30636
rect 9213 30635 9279 30636
rect 10593 30635 10659 30636
rect 10961 30635 11027 30638
rect 11605 30698 11671 30701
rect 16982 30698 16988 30700
rect 11605 30696 16988 30698
rect 11605 30640 11610 30696
rect 11666 30640 16988 30696
rect 11605 30638 16988 30640
rect 11605 30635 11671 30638
rect 16982 30636 16988 30638
rect 17052 30636 17058 30700
rect 0 30562 160 30592
rect 3417 30562 3483 30565
rect 6085 30562 6151 30565
rect 0 30560 3483 30562
rect 0 30504 3422 30560
rect 3478 30504 3483 30560
rect 0 30502 3483 30504
rect 0 30472 160 30502
rect 3417 30499 3483 30502
rect 3558 30560 6151 30562
rect 3558 30504 6090 30560
rect 6146 30504 6151 30560
rect 3558 30502 6151 30504
rect 1301 30426 1367 30429
rect 2078 30426 2084 30428
rect 1301 30424 2084 30426
rect 1301 30368 1306 30424
rect 1362 30368 2084 30424
rect 1301 30366 2084 30368
rect 1301 30363 1367 30366
rect 2078 30364 2084 30366
rect 2148 30364 2154 30428
rect 2221 30426 2287 30429
rect 3558 30426 3618 30502
rect 6085 30499 6151 30502
rect 7833 30562 7899 30565
rect 11881 30562 11947 30565
rect 7833 30560 11947 30562
rect 7833 30504 7838 30560
rect 7894 30504 11886 30560
rect 11942 30504 11947 30560
rect 7833 30502 11947 30504
rect 7833 30499 7899 30502
rect 11881 30499 11947 30502
rect 25129 30562 25195 30565
rect 25840 30562 26000 30592
rect 25129 30560 26000 30562
rect 25129 30504 25134 30560
rect 25190 30504 26000 30560
rect 25129 30502 26000 30504
rect 25129 30499 25195 30502
rect 6880 30496 7196 30497
rect 6880 30432 6886 30496
rect 6950 30432 6966 30496
rect 7030 30432 7046 30496
rect 7110 30432 7126 30496
rect 7190 30432 7196 30496
rect 6880 30431 7196 30432
rect 12814 30496 13130 30497
rect 12814 30432 12820 30496
rect 12884 30432 12900 30496
rect 12964 30432 12980 30496
rect 13044 30432 13060 30496
rect 13124 30432 13130 30496
rect 12814 30431 13130 30432
rect 18748 30496 19064 30497
rect 18748 30432 18754 30496
rect 18818 30432 18834 30496
rect 18898 30432 18914 30496
rect 18978 30432 18994 30496
rect 19058 30432 19064 30496
rect 18748 30431 19064 30432
rect 24682 30496 24998 30497
rect 24682 30432 24688 30496
rect 24752 30432 24768 30496
rect 24832 30432 24848 30496
rect 24912 30432 24928 30496
rect 24992 30432 24998 30496
rect 25840 30472 26000 30502
rect 24682 30431 24998 30432
rect 2221 30424 3618 30426
rect 2221 30368 2226 30424
rect 2282 30368 3618 30424
rect 2221 30366 3618 30368
rect 4245 30426 4311 30429
rect 5809 30426 5875 30429
rect 4245 30424 5875 30426
rect 4245 30368 4250 30424
rect 4306 30368 5814 30424
rect 5870 30368 5875 30424
rect 4245 30366 5875 30368
rect 2221 30363 2287 30366
rect 4245 30363 4311 30366
rect 5809 30363 5875 30366
rect 8109 30426 8175 30429
rect 8334 30426 8340 30428
rect 8109 30424 8340 30426
rect 8109 30368 8114 30424
rect 8170 30368 8340 30424
rect 8109 30366 8340 30368
rect 8109 30363 8175 30366
rect 8334 30364 8340 30366
rect 8404 30364 8410 30428
rect 8702 30364 8708 30428
rect 8772 30426 8778 30428
rect 9397 30426 9463 30429
rect 8772 30424 9463 30426
rect 8772 30368 9402 30424
rect 9458 30368 9463 30424
rect 8772 30366 9463 30368
rect 8772 30364 8778 30366
rect 9397 30363 9463 30366
rect 9581 30426 9647 30429
rect 12617 30426 12683 30429
rect 9581 30424 12683 30426
rect 9581 30368 9586 30424
rect 9642 30368 12622 30424
rect 12678 30368 12683 30424
rect 9581 30366 12683 30368
rect 9581 30363 9647 30366
rect 12617 30363 12683 30366
rect 0 30290 160 30320
rect 3785 30290 3851 30293
rect 0 30288 3851 30290
rect 0 30232 3790 30288
rect 3846 30232 3851 30288
rect 0 30230 3851 30232
rect 0 30200 160 30230
rect 3785 30227 3851 30230
rect 5257 30290 5323 30293
rect 6453 30290 6519 30293
rect 5257 30288 6519 30290
rect 5257 30232 5262 30288
rect 5318 30232 6458 30288
rect 6514 30232 6519 30288
rect 5257 30230 6519 30232
rect 5257 30227 5323 30230
rect 6453 30227 6519 30230
rect 6729 30290 6795 30293
rect 10910 30290 10916 30292
rect 6729 30288 10916 30290
rect 6729 30232 6734 30288
rect 6790 30232 10916 30288
rect 6729 30230 10916 30232
rect 6729 30227 6795 30230
rect 10910 30228 10916 30230
rect 10980 30290 10986 30292
rect 11053 30290 11119 30293
rect 10980 30288 11119 30290
rect 10980 30232 11058 30288
rect 11114 30232 11119 30288
rect 10980 30230 11119 30232
rect 10980 30228 10986 30230
rect 11053 30227 11119 30230
rect 11789 30290 11855 30293
rect 14917 30290 14983 30293
rect 11789 30288 14983 30290
rect 11789 30232 11794 30288
rect 11850 30232 14922 30288
rect 14978 30232 14983 30288
rect 11789 30230 14983 30232
rect 11789 30227 11855 30230
rect 14917 30227 14983 30230
rect 3417 30154 3483 30157
rect 11237 30154 11303 30157
rect 3417 30152 11303 30154
rect 3417 30096 3422 30152
rect 3478 30096 11242 30152
rect 11298 30096 11303 30152
rect 3417 30094 11303 30096
rect 3417 30091 3483 30094
rect 0 30018 160 30048
rect 1485 30018 1551 30021
rect 0 30016 1551 30018
rect 0 29960 1490 30016
rect 1546 29960 1551 30016
rect 0 29958 1551 29960
rect 0 29928 160 29958
rect 1485 29955 1551 29958
rect 0 29746 160 29776
rect 933 29746 999 29749
rect 0 29744 999 29746
rect 0 29688 938 29744
rect 994 29688 999 29744
rect 0 29686 999 29688
rect 0 29656 160 29686
rect 933 29683 999 29686
rect 1577 29746 1643 29749
rect 3742 29746 3802 30094
rect 11237 30091 11303 30094
rect 6126 29956 6132 30020
rect 6196 30018 6202 30020
rect 6545 30018 6611 30021
rect 6196 30016 6611 30018
rect 6196 29960 6550 30016
rect 6606 29960 6611 30016
rect 6196 29958 6611 29960
rect 6196 29956 6202 29958
rect 6545 29955 6611 29958
rect 24393 30018 24459 30021
rect 25840 30018 26000 30048
rect 24393 30016 26000 30018
rect 24393 29960 24398 30016
rect 24454 29960 26000 30016
rect 24393 29958 26000 29960
rect 24393 29955 24459 29958
rect 3913 29952 4229 29953
rect 3913 29888 3919 29952
rect 3983 29888 3999 29952
rect 4063 29888 4079 29952
rect 4143 29888 4159 29952
rect 4223 29888 4229 29952
rect 3913 29887 4229 29888
rect 9847 29952 10163 29953
rect 9847 29888 9853 29952
rect 9917 29888 9933 29952
rect 9997 29888 10013 29952
rect 10077 29888 10093 29952
rect 10157 29888 10163 29952
rect 9847 29887 10163 29888
rect 15781 29952 16097 29953
rect 15781 29888 15787 29952
rect 15851 29888 15867 29952
rect 15931 29888 15947 29952
rect 16011 29888 16027 29952
rect 16091 29888 16097 29952
rect 15781 29887 16097 29888
rect 21715 29952 22031 29953
rect 21715 29888 21721 29952
rect 21785 29888 21801 29952
rect 21865 29888 21881 29952
rect 21945 29888 21961 29952
rect 22025 29888 22031 29952
rect 25840 29928 26000 29958
rect 21715 29887 22031 29888
rect 3877 29746 3943 29749
rect 1577 29744 2790 29746
rect 1577 29688 1582 29744
rect 1638 29688 2790 29744
rect 1577 29686 2790 29688
rect 3742 29744 3943 29746
rect 3742 29688 3882 29744
rect 3938 29688 3943 29744
rect 3742 29686 3943 29688
rect 1577 29683 1643 29686
rect 2730 29610 2790 29686
rect 3877 29683 3943 29686
rect 7465 29746 7531 29749
rect 9489 29746 9555 29749
rect 7465 29744 17050 29746
rect 7465 29688 7470 29744
rect 7526 29688 9494 29744
rect 9550 29688 17050 29744
rect 7465 29686 17050 29688
rect 7465 29683 7531 29686
rect 9489 29683 9555 29686
rect 16757 29610 16823 29613
rect 2730 29608 16823 29610
rect 2730 29552 16762 29608
rect 16818 29552 16823 29608
rect 2730 29550 16823 29552
rect 16757 29547 16823 29550
rect 0 29474 160 29504
rect 1117 29474 1183 29477
rect 0 29472 1183 29474
rect 0 29416 1122 29472
rect 1178 29416 1183 29472
rect 0 29414 1183 29416
rect 0 29384 160 29414
rect 1117 29411 1183 29414
rect 1761 29474 1827 29477
rect 6453 29474 6519 29477
rect 1761 29472 6519 29474
rect 1761 29416 1766 29472
rect 1822 29416 6458 29472
rect 6514 29416 6519 29472
rect 1761 29414 6519 29416
rect 1761 29411 1827 29414
rect 6453 29411 6519 29414
rect 7281 29474 7347 29477
rect 7281 29472 12450 29474
rect 7281 29416 7286 29472
rect 7342 29416 12450 29472
rect 7281 29414 12450 29416
rect 7281 29411 7347 29414
rect 6880 29408 7196 29409
rect 6880 29344 6886 29408
rect 6950 29344 6966 29408
rect 7030 29344 7046 29408
rect 7110 29344 7126 29408
rect 7190 29344 7196 29408
rect 6880 29343 7196 29344
rect 3601 29338 3667 29341
rect 6085 29338 6151 29341
rect 3601 29336 6151 29338
rect 3601 29280 3606 29336
rect 3662 29280 6090 29336
rect 6146 29280 6151 29336
rect 3601 29278 6151 29280
rect 3601 29275 3667 29278
rect 6085 29275 6151 29278
rect 8201 29338 8267 29341
rect 8753 29338 8819 29341
rect 8201 29336 8819 29338
rect 8201 29280 8206 29336
rect 8262 29280 8758 29336
rect 8814 29280 8819 29336
rect 8201 29278 8819 29280
rect 8201 29275 8267 29278
rect 8753 29275 8819 29278
rect 10133 29338 10199 29341
rect 10133 29336 12312 29338
rect 10133 29280 10138 29336
rect 10194 29280 12312 29336
rect 10133 29278 12312 29280
rect 10133 29275 10199 29278
rect 0 29202 160 29232
rect 1301 29202 1367 29205
rect 0 29200 1367 29202
rect 0 29144 1306 29200
rect 1362 29144 1367 29200
rect 0 29142 1367 29144
rect 0 29112 160 29142
rect 1301 29139 1367 29142
rect 3141 29202 3207 29205
rect 4286 29202 4292 29204
rect 3141 29200 4292 29202
rect 3141 29144 3146 29200
rect 3202 29144 4292 29200
rect 3141 29142 4292 29144
rect 3141 29139 3207 29142
rect 4286 29140 4292 29142
rect 4356 29140 4362 29204
rect 4981 29202 5047 29205
rect 11053 29202 11119 29205
rect 4981 29200 11119 29202
rect 4981 29144 4986 29200
rect 5042 29144 11058 29200
rect 11114 29144 11119 29200
rect 4981 29142 11119 29144
rect 4981 29139 5047 29142
rect 11053 29139 11119 29142
rect 2037 29066 2103 29069
rect 5073 29068 5139 29069
rect 2037 29064 4906 29066
rect 2037 29008 2042 29064
rect 2098 29008 4906 29064
rect 2037 29006 4906 29008
rect 2037 29003 2103 29006
rect 0 28930 160 28960
rect 3601 28930 3667 28933
rect 0 28928 3667 28930
rect 0 28872 3606 28928
rect 3662 28872 3667 28928
rect 0 28870 3667 28872
rect 4846 28930 4906 29006
rect 5022 29004 5028 29068
rect 5092 29066 5139 29068
rect 8753 29066 8819 29069
rect 9581 29066 9647 29069
rect 5092 29064 5184 29066
rect 5134 29008 5184 29064
rect 5092 29006 5184 29008
rect 5398 29064 9647 29066
rect 5398 29008 8758 29064
rect 8814 29008 9586 29064
rect 9642 29008 9647 29064
rect 5398 29006 9647 29008
rect 5092 29004 5139 29006
rect 5073 29003 5139 29004
rect 5398 28930 5458 29006
rect 8753 29003 8819 29006
rect 9581 29003 9647 29006
rect 11789 29068 11855 29069
rect 11789 29064 11836 29068
rect 11900 29066 11906 29068
rect 12252 29066 12312 29278
rect 12390 29202 12450 29414
rect 16614 29412 16620 29476
rect 16684 29474 16690 29476
rect 16849 29474 16915 29477
rect 16990 29474 17050 29686
rect 17718 29684 17724 29748
rect 17788 29746 17794 29748
rect 22093 29746 22159 29749
rect 17788 29744 22159 29746
rect 17788 29688 22098 29744
rect 22154 29688 22159 29744
rect 17788 29686 22159 29688
rect 17788 29684 17794 29686
rect 22093 29683 22159 29686
rect 16684 29472 17050 29474
rect 16684 29416 16854 29472
rect 16910 29416 17050 29472
rect 16684 29414 17050 29416
rect 25129 29474 25195 29477
rect 25840 29474 26000 29504
rect 25129 29472 26000 29474
rect 25129 29416 25134 29472
rect 25190 29416 26000 29472
rect 25129 29414 26000 29416
rect 16684 29412 16690 29414
rect 16849 29411 16915 29414
rect 25129 29411 25195 29414
rect 12814 29408 13130 29409
rect 12814 29344 12820 29408
rect 12884 29344 12900 29408
rect 12964 29344 12980 29408
rect 13044 29344 13060 29408
rect 13124 29344 13130 29408
rect 12814 29343 13130 29344
rect 18748 29408 19064 29409
rect 18748 29344 18754 29408
rect 18818 29344 18834 29408
rect 18898 29344 18914 29408
rect 18978 29344 18994 29408
rect 19058 29344 19064 29408
rect 18748 29343 19064 29344
rect 24682 29408 24998 29409
rect 24682 29344 24688 29408
rect 24752 29344 24768 29408
rect 24832 29344 24848 29408
rect 24912 29344 24928 29408
rect 24992 29344 24998 29408
rect 25840 29384 26000 29414
rect 24682 29343 24998 29344
rect 15837 29338 15903 29341
rect 17585 29338 17651 29341
rect 15837 29336 17651 29338
rect 15837 29280 15842 29336
rect 15898 29280 17590 29336
rect 17646 29280 17651 29336
rect 15837 29278 17651 29280
rect 15837 29275 15903 29278
rect 17585 29275 17651 29278
rect 15469 29202 15535 29205
rect 12390 29200 15535 29202
rect 12390 29144 15474 29200
rect 15530 29144 15535 29200
rect 12390 29142 15535 29144
rect 15469 29139 15535 29142
rect 13813 29066 13879 29069
rect 11789 29008 11794 29064
rect 11789 29004 11836 29008
rect 11900 29006 11946 29066
rect 12252 29064 13879 29066
rect 12252 29008 13818 29064
rect 13874 29008 13879 29064
rect 12252 29006 13879 29008
rect 11900 29004 11906 29006
rect 11789 29003 11855 29004
rect 13813 29003 13879 29006
rect 20069 29066 20135 29069
rect 20846 29066 20852 29068
rect 20069 29064 20852 29066
rect 20069 29008 20074 29064
rect 20130 29008 20852 29064
rect 20069 29006 20852 29008
rect 20069 29003 20135 29006
rect 20846 29004 20852 29006
rect 20916 29004 20922 29068
rect 4846 28870 5458 28930
rect 0 28840 160 28870
rect 3601 28867 3667 28870
rect 10910 28868 10916 28932
rect 10980 28930 10986 28932
rect 12525 28930 12591 28933
rect 10980 28928 12591 28930
rect 10980 28872 12530 28928
rect 12586 28872 12591 28928
rect 10980 28870 12591 28872
rect 10980 28868 10986 28870
rect 12525 28867 12591 28870
rect 24393 28930 24459 28933
rect 25840 28930 26000 28960
rect 24393 28928 26000 28930
rect 24393 28872 24398 28928
rect 24454 28872 26000 28928
rect 24393 28870 26000 28872
rect 24393 28867 24459 28870
rect 3913 28864 4229 28865
rect 3913 28800 3919 28864
rect 3983 28800 3999 28864
rect 4063 28800 4079 28864
rect 4143 28800 4159 28864
rect 4223 28800 4229 28864
rect 3913 28799 4229 28800
rect 9847 28864 10163 28865
rect 9847 28800 9853 28864
rect 9917 28800 9933 28864
rect 9997 28800 10013 28864
rect 10077 28800 10093 28864
rect 10157 28800 10163 28864
rect 9847 28799 10163 28800
rect 15781 28864 16097 28865
rect 15781 28800 15787 28864
rect 15851 28800 15867 28864
rect 15931 28800 15947 28864
rect 16011 28800 16027 28864
rect 16091 28800 16097 28864
rect 15781 28799 16097 28800
rect 21715 28864 22031 28865
rect 21715 28800 21721 28864
rect 21785 28800 21801 28864
rect 21865 28800 21881 28864
rect 21945 28800 21961 28864
rect 22025 28800 22031 28864
rect 25840 28840 26000 28870
rect 21715 28799 22031 28800
rect 1117 28794 1183 28797
rect 3049 28794 3115 28797
rect 1117 28792 3115 28794
rect 1117 28736 1122 28792
rect 1178 28736 3054 28792
rect 3110 28736 3115 28792
rect 1117 28734 3115 28736
rect 1117 28731 1183 28734
rect 3049 28731 3115 28734
rect 4470 28732 4476 28796
rect 4540 28794 4546 28796
rect 7189 28794 7255 28797
rect 4540 28792 7255 28794
rect 4540 28736 7194 28792
rect 7250 28736 7255 28792
rect 4540 28734 7255 28736
rect 4540 28732 4546 28734
rect 7189 28731 7255 28734
rect 0 28658 160 28688
rect 933 28658 999 28661
rect 0 28656 999 28658
rect 0 28600 938 28656
rect 994 28600 999 28656
rect 0 28598 999 28600
rect 0 28568 160 28598
rect 933 28595 999 28598
rect 2078 28596 2084 28660
rect 2148 28658 2154 28660
rect 2497 28658 2563 28661
rect 2148 28656 2563 28658
rect 2148 28600 2502 28656
rect 2558 28600 2563 28656
rect 2148 28598 2563 28600
rect 2148 28596 2154 28598
rect 2497 28595 2563 28598
rect 4654 28596 4660 28660
rect 4724 28658 4730 28660
rect 15101 28658 15167 28661
rect 23197 28658 23263 28661
rect 4724 28656 23263 28658
rect 4724 28600 15106 28656
rect 15162 28600 23202 28656
rect 23258 28600 23263 28656
rect 4724 28598 23263 28600
rect 4724 28596 4730 28598
rect 15101 28595 15167 28598
rect 23197 28595 23263 28598
rect 749 28522 815 28525
rect 2446 28522 2452 28524
rect 749 28520 2452 28522
rect 749 28464 754 28520
rect 810 28464 2452 28520
rect 749 28462 2452 28464
rect 749 28459 815 28462
rect 2446 28460 2452 28462
rect 2516 28460 2522 28524
rect 4889 28522 4955 28525
rect 8886 28522 8892 28524
rect 4889 28520 8892 28522
rect 4889 28464 4894 28520
rect 4950 28464 8892 28520
rect 4889 28462 8892 28464
rect 4889 28459 4955 28462
rect 8886 28460 8892 28462
rect 8956 28522 8962 28524
rect 9489 28522 9555 28525
rect 13670 28522 13676 28524
rect 8956 28520 13676 28522
rect 8956 28464 9494 28520
rect 9550 28464 13676 28520
rect 8956 28462 13676 28464
rect 8956 28460 8962 28462
rect 9489 28459 9555 28462
rect 13670 28460 13676 28462
rect 13740 28522 13746 28524
rect 20713 28522 20779 28525
rect 13740 28520 20779 28522
rect 13740 28464 20718 28520
rect 20774 28464 20779 28520
rect 13740 28462 20779 28464
rect 13740 28460 13746 28462
rect 20713 28459 20779 28462
rect 0 28386 160 28416
rect 1485 28386 1551 28389
rect 0 28384 1551 28386
rect 0 28328 1490 28384
rect 1546 28328 1551 28384
rect 0 28326 1551 28328
rect 0 28296 160 28326
rect 1485 28323 1551 28326
rect 25129 28386 25195 28389
rect 25840 28386 26000 28416
rect 25129 28384 26000 28386
rect 25129 28328 25134 28384
rect 25190 28328 26000 28384
rect 25129 28326 26000 28328
rect 25129 28323 25195 28326
rect 6880 28320 7196 28321
rect 6880 28256 6886 28320
rect 6950 28256 6966 28320
rect 7030 28256 7046 28320
rect 7110 28256 7126 28320
rect 7190 28256 7196 28320
rect 6880 28255 7196 28256
rect 12814 28320 13130 28321
rect 12814 28256 12820 28320
rect 12884 28256 12900 28320
rect 12964 28256 12980 28320
rect 13044 28256 13060 28320
rect 13124 28256 13130 28320
rect 12814 28255 13130 28256
rect 18748 28320 19064 28321
rect 18748 28256 18754 28320
rect 18818 28256 18834 28320
rect 18898 28256 18914 28320
rect 18978 28256 18994 28320
rect 19058 28256 19064 28320
rect 18748 28255 19064 28256
rect 24682 28320 24998 28321
rect 24682 28256 24688 28320
rect 24752 28256 24768 28320
rect 24832 28256 24848 28320
rect 24912 28256 24928 28320
rect 24992 28256 24998 28320
rect 25840 28296 26000 28326
rect 24682 28255 24998 28256
rect 1945 28250 2011 28253
rect 3877 28250 3943 28253
rect 1945 28248 3943 28250
rect 1945 28192 1950 28248
rect 2006 28192 3882 28248
rect 3938 28192 3943 28248
rect 1945 28190 3943 28192
rect 1945 28187 2011 28190
rect 3877 28187 3943 28190
rect 10041 28250 10107 28253
rect 12065 28250 12131 28253
rect 10041 28248 12131 28250
rect 10041 28192 10046 28248
rect 10102 28192 12070 28248
rect 12126 28192 12131 28248
rect 10041 28190 12131 28192
rect 10041 28187 10107 28190
rect 12065 28187 12131 28190
rect 0 28114 160 28144
rect 841 28114 907 28117
rect 0 28112 907 28114
rect 0 28056 846 28112
rect 902 28056 907 28112
rect 0 28054 907 28056
rect 0 28024 160 28054
rect 841 28051 907 28054
rect 1853 28114 1919 28117
rect 8845 28114 8911 28117
rect 1853 28112 8911 28114
rect 1853 28056 1858 28112
rect 1914 28056 8850 28112
rect 8906 28056 8911 28112
rect 1853 28054 8911 28056
rect 1853 28051 1919 28054
rect 8845 28051 8911 28054
rect 12433 28114 12499 28117
rect 17493 28114 17559 28117
rect 12433 28112 17559 28114
rect 12433 28056 12438 28112
rect 12494 28056 17498 28112
rect 17554 28056 17559 28112
rect 12433 28054 17559 28056
rect 12433 28051 12499 28054
rect 17493 28051 17559 28054
rect 1710 27916 1716 27980
rect 1780 27978 1786 27980
rect 2405 27978 2471 27981
rect 1780 27976 2471 27978
rect 1780 27920 2410 27976
rect 2466 27920 2471 27976
rect 1780 27918 2471 27920
rect 1780 27916 1786 27918
rect 2405 27915 2471 27918
rect 2681 27978 2747 27981
rect 17125 27978 17191 27981
rect 2681 27976 17191 27978
rect 2681 27920 2686 27976
rect 2742 27920 17130 27976
rect 17186 27920 17191 27976
rect 2681 27918 17191 27920
rect 2681 27915 2747 27918
rect 17125 27915 17191 27918
rect 0 27842 160 27872
rect 749 27842 815 27845
rect 0 27840 815 27842
rect 0 27784 754 27840
rect 810 27784 815 27840
rect 0 27782 815 27784
rect 0 27752 160 27782
rect 749 27779 815 27782
rect 4981 27842 5047 27845
rect 6085 27842 6151 27845
rect 4981 27840 6151 27842
rect 4981 27784 4986 27840
rect 5042 27784 6090 27840
rect 6146 27784 6151 27840
rect 4981 27782 6151 27784
rect 4981 27779 5047 27782
rect 6085 27779 6151 27782
rect 14089 27842 14155 27845
rect 14457 27842 14523 27845
rect 14089 27840 14523 27842
rect 14089 27784 14094 27840
rect 14150 27784 14462 27840
rect 14518 27784 14523 27840
rect 14089 27782 14523 27784
rect 14089 27779 14155 27782
rect 14457 27779 14523 27782
rect 24393 27842 24459 27845
rect 25840 27842 26000 27872
rect 24393 27840 26000 27842
rect 24393 27784 24398 27840
rect 24454 27784 26000 27840
rect 24393 27782 26000 27784
rect 24393 27779 24459 27782
rect 3913 27776 4229 27777
rect 3913 27712 3919 27776
rect 3983 27712 3999 27776
rect 4063 27712 4079 27776
rect 4143 27712 4159 27776
rect 4223 27712 4229 27776
rect 3913 27711 4229 27712
rect 9847 27776 10163 27777
rect 9847 27712 9853 27776
rect 9917 27712 9933 27776
rect 9997 27712 10013 27776
rect 10077 27712 10093 27776
rect 10157 27712 10163 27776
rect 9847 27711 10163 27712
rect 15781 27776 16097 27777
rect 15781 27712 15787 27776
rect 15851 27712 15867 27776
rect 15931 27712 15947 27776
rect 16011 27712 16027 27776
rect 16091 27712 16097 27776
rect 15781 27711 16097 27712
rect 21715 27776 22031 27777
rect 21715 27712 21721 27776
rect 21785 27712 21801 27776
rect 21865 27712 21881 27776
rect 21945 27712 21961 27776
rect 22025 27712 22031 27776
rect 25840 27752 26000 27782
rect 21715 27711 22031 27712
rect 1393 27706 1459 27709
rect 982 27704 1459 27706
rect 982 27648 1398 27704
rect 1454 27648 1459 27704
rect 982 27646 1459 27648
rect 0 27570 160 27600
rect 982 27570 1042 27646
rect 1393 27643 1459 27646
rect 7557 27706 7623 27709
rect 14917 27706 14983 27709
rect 7557 27704 7666 27706
rect 7557 27648 7562 27704
rect 7618 27648 7666 27704
rect 7557 27643 7666 27648
rect 2313 27570 2379 27573
rect 0 27510 1042 27570
rect 1166 27568 2379 27570
rect 1166 27512 2318 27568
rect 2374 27512 2379 27568
rect 1166 27510 2379 27512
rect 0 27480 160 27510
rect 0 27298 160 27328
rect 1166 27298 1226 27510
rect 2313 27507 2379 27510
rect 6085 27570 6151 27573
rect 7606 27570 7666 27643
rect 12390 27704 14983 27706
rect 12390 27648 14922 27704
rect 14978 27648 14983 27704
rect 12390 27646 14983 27648
rect 12390 27570 12450 27646
rect 14917 27643 14983 27646
rect 16573 27706 16639 27709
rect 17534 27706 17540 27708
rect 16573 27704 17540 27706
rect 16573 27648 16578 27704
rect 16634 27648 17540 27704
rect 16573 27646 17540 27648
rect 16573 27643 16639 27646
rect 17534 27644 17540 27646
rect 17604 27644 17610 27708
rect 6085 27568 12450 27570
rect 6085 27512 6090 27568
rect 6146 27512 12450 27568
rect 6085 27510 12450 27512
rect 16205 27570 16271 27573
rect 17309 27570 17375 27573
rect 16205 27568 17375 27570
rect 16205 27512 16210 27568
rect 16266 27512 17314 27568
rect 17370 27512 17375 27568
rect 16205 27510 17375 27512
rect 6085 27507 6151 27510
rect 16205 27507 16271 27510
rect 17309 27507 17375 27510
rect 10777 27434 10843 27437
rect 13169 27434 13235 27437
rect 0 27238 1226 27298
rect 1534 27432 10843 27434
rect 1534 27376 10782 27432
rect 10838 27376 10843 27432
rect 1534 27374 10843 27376
rect 0 27208 160 27238
rect 473 27162 539 27165
rect 1534 27162 1594 27374
rect 10777 27371 10843 27374
rect 12390 27432 13235 27434
rect 12390 27376 13174 27432
rect 13230 27376 13235 27432
rect 12390 27374 13235 27376
rect 2589 27298 2655 27301
rect 6361 27298 6427 27301
rect 2589 27296 6427 27298
rect 2589 27240 2594 27296
rect 2650 27240 6366 27296
rect 6422 27240 6427 27296
rect 2589 27238 6427 27240
rect 2589 27235 2655 27238
rect 6361 27235 6427 27238
rect 7414 27236 7420 27300
rect 7484 27298 7490 27300
rect 12390 27298 12450 27374
rect 13169 27371 13235 27374
rect 15326 27372 15332 27436
rect 15396 27434 15402 27436
rect 17217 27434 17283 27437
rect 15396 27432 17283 27434
rect 15396 27376 17222 27432
rect 17278 27376 17283 27432
rect 15396 27374 17283 27376
rect 15396 27372 15402 27374
rect 17217 27371 17283 27374
rect 16481 27300 16547 27301
rect 7484 27238 12450 27298
rect 7484 27236 7490 27238
rect 16430 27236 16436 27300
rect 16500 27298 16547 27300
rect 25129 27298 25195 27301
rect 25840 27298 26000 27328
rect 16500 27296 16592 27298
rect 16542 27240 16592 27296
rect 16500 27238 16592 27240
rect 25129 27296 26000 27298
rect 25129 27240 25134 27296
rect 25190 27240 26000 27296
rect 25129 27238 26000 27240
rect 16500 27236 16547 27238
rect 16481 27235 16547 27236
rect 25129 27235 25195 27238
rect 6880 27232 7196 27233
rect 6880 27168 6886 27232
rect 6950 27168 6966 27232
rect 7030 27168 7046 27232
rect 7110 27168 7126 27232
rect 7190 27168 7196 27232
rect 6880 27167 7196 27168
rect 12814 27232 13130 27233
rect 12814 27168 12820 27232
rect 12884 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13130 27232
rect 12814 27167 13130 27168
rect 18748 27232 19064 27233
rect 18748 27168 18754 27232
rect 18818 27168 18834 27232
rect 18898 27168 18914 27232
rect 18978 27168 18994 27232
rect 19058 27168 19064 27232
rect 18748 27167 19064 27168
rect 24682 27232 24998 27233
rect 24682 27168 24688 27232
rect 24752 27168 24768 27232
rect 24832 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 24998 27232
rect 25840 27208 26000 27238
rect 24682 27167 24998 27168
rect 473 27160 1594 27162
rect 473 27104 478 27160
rect 534 27104 1594 27160
rect 473 27102 1594 27104
rect 473 27099 539 27102
rect 0 27026 160 27056
rect 1301 27026 1367 27029
rect 0 27024 1367 27026
rect 0 26968 1306 27024
rect 1362 26968 1367 27024
rect 0 26966 1367 26968
rect 0 26936 160 26966
rect 1301 26963 1367 26966
rect 6126 26964 6132 27028
rect 6196 27026 6202 27028
rect 9949 27026 10015 27029
rect 11094 27026 11100 27028
rect 6196 26966 7850 27026
rect 6196 26964 6202 26966
rect 473 26890 539 26893
rect 7649 26890 7715 26893
rect 473 26888 7715 26890
rect 473 26832 478 26888
rect 534 26832 7654 26888
rect 7710 26832 7715 26888
rect 473 26830 7715 26832
rect 7790 26890 7850 26966
rect 9949 27024 11100 27026
rect 9949 26968 9954 27024
rect 10010 26968 11100 27024
rect 9949 26966 11100 26968
rect 9949 26963 10015 26966
rect 11094 26964 11100 26966
rect 11164 26964 11170 27028
rect 13629 27026 13695 27029
rect 20069 27026 20135 27029
rect 21265 27028 21331 27029
rect 21214 27026 21220 27028
rect 13629 27024 20135 27026
rect 13629 26968 13634 27024
rect 13690 26968 20074 27024
rect 20130 26968 20135 27024
rect 13629 26966 20135 26968
rect 21174 26966 21220 27026
rect 21284 27024 21331 27028
rect 21326 26968 21331 27024
rect 13629 26963 13695 26966
rect 20069 26963 20135 26966
rect 21214 26964 21220 26966
rect 21284 26964 21331 26968
rect 21265 26963 21331 26964
rect 15101 26890 15167 26893
rect 7790 26888 15167 26890
rect 7790 26832 15106 26888
rect 15162 26832 15167 26888
rect 7790 26830 15167 26832
rect 473 26827 539 26830
rect 7649 26827 7715 26830
rect 15101 26827 15167 26830
rect 15510 26828 15516 26892
rect 15580 26890 15586 26892
rect 20294 26890 20300 26892
rect 15580 26830 20300 26890
rect 15580 26828 15586 26830
rect 20294 26828 20300 26830
rect 20364 26828 20370 26892
rect 0 26754 160 26784
rect 1209 26754 1275 26757
rect 17309 26756 17375 26757
rect 17309 26754 17356 26756
rect 0 26752 1275 26754
rect 0 26696 1214 26752
rect 1270 26696 1275 26752
rect 0 26694 1275 26696
rect 17264 26752 17356 26754
rect 17264 26696 17314 26752
rect 17264 26694 17356 26696
rect 0 26664 160 26694
rect 1209 26691 1275 26694
rect 17309 26692 17356 26694
rect 17420 26692 17426 26756
rect 24393 26754 24459 26757
rect 25840 26754 26000 26784
rect 24393 26752 26000 26754
rect 24393 26696 24398 26752
rect 24454 26696 26000 26752
rect 24393 26694 26000 26696
rect 17309 26691 17375 26692
rect 24393 26691 24459 26694
rect 3913 26688 4229 26689
rect 3913 26624 3919 26688
rect 3983 26624 3999 26688
rect 4063 26624 4079 26688
rect 4143 26624 4159 26688
rect 4223 26624 4229 26688
rect 3913 26623 4229 26624
rect 9847 26688 10163 26689
rect 9847 26624 9853 26688
rect 9917 26624 9933 26688
rect 9997 26624 10013 26688
rect 10077 26624 10093 26688
rect 10157 26624 10163 26688
rect 9847 26623 10163 26624
rect 15781 26688 16097 26689
rect 15781 26624 15787 26688
rect 15851 26624 15867 26688
rect 15931 26624 15947 26688
rect 16011 26624 16027 26688
rect 16091 26624 16097 26688
rect 15781 26623 16097 26624
rect 21715 26688 22031 26689
rect 21715 26624 21721 26688
rect 21785 26624 21801 26688
rect 21865 26624 21881 26688
rect 21945 26624 21961 26688
rect 22025 26624 22031 26688
rect 25840 26664 26000 26694
rect 21715 26623 22031 26624
rect 6085 26618 6151 26621
rect 9581 26618 9647 26621
rect 6085 26616 9647 26618
rect 6085 26560 6090 26616
rect 6146 26560 9586 26616
rect 9642 26560 9647 26616
rect 6085 26558 9647 26560
rect 6085 26555 6151 26558
rect 9581 26555 9647 26558
rect 0 26482 160 26512
rect 1117 26482 1183 26485
rect 0 26480 1183 26482
rect 0 26424 1122 26480
rect 1178 26424 1183 26480
rect 0 26422 1183 26424
rect 0 26392 160 26422
rect 1117 26419 1183 26422
rect 1853 26482 1919 26485
rect 6821 26482 6887 26485
rect 1853 26480 6887 26482
rect 1853 26424 1858 26480
rect 1914 26424 6826 26480
rect 6882 26424 6887 26480
rect 1853 26422 6887 26424
rect 1853 26419 1919 26422
rect 6821 26419 6887 26422
rect 10133 26482 10199 26485
rect 10777 26482 10843 26485
rect 10133 26480 10843 26482
rect 10133 26424 10138 26480
rect 10194 26424 10782 26480
rect 10838 26424 10843 26480
rect 10133 26422 10843 26424
rect 10133 26419 10199 26422
rect 10777 26419 10843 26422
rect 11329 26482 11395 26485
rect 18689 26482 18755 26485
rect 11329 26480 18755 26482
rect 11329 26424 11334 26480
rect 11390 26424 18694 26480
rect 18750 26424 18755 26480
rect 11329 26422 18755 26424
rect 11329 26419 11395 26422
rect 18689 26419 18755 26422
rect 1894 26284 1900 26348
rect 1964 26346 1970 26348
rect 2037 26346 2103 26349
rect 1964 26344 2103 26346
rect 1964 26288 2042 26344
rect 2098 26288 2103 26344
rect 1964 26286 2103 26288
rect 1964 26284 1970 26286
rect 2037 26283 2103 26286
rect 0 26210 160 26240
rect 2589 26210 2655 26213
rect 11697 26212 11763 26213
rect 11646 26210 11652 26212
rect 0 26208 2655 26210
rect 0 26152 2594 26208
rect 2650 26152 2655 26208
rect 0 26150 2655 26152
rect 11606 26150 11652 26210
rect 11716 26208 11763 26212
rect 11758 26152 11763 26208
rect 0 26120 160 26150
rect 2589 26147 2655 26150
rect 11646 26148 11652 26150
rect 11716 26148 11763 26152
rect 11697 26147 11763 26148
rect 21633 26210 21699 26213
rect 24209 26210 24275 26213
rect 21633 26208 24275 26210
rect 21633 26152 21638 26208
rect 21694 26152 24214 26208
rect 24270 26152 24275 26208
rect 21633 26150 24275 26152
rect 21633 26147 21699 26150
rect 24209 26147 24275 26150
rect 25129 26210 25195 26213
rect 25840 26210 26000 26240
rect 25129 26208 26000 26210
rect 25129 26152 25134 26208
rect 25190 26152 26000 26208
rect 25129 26150 26000 26152
rect 25129 26147 25195 26150
rect 6880 26144 7196 26145
rect 6880 26080 6886 26144
rect 6950 26080 6966 26144
rect 7030 26080 7046 26144
rect 7110 26080 7126 26144
rect 7190 26080 7196 26144
rect 6880 26079 7196 26080
rect 12814 26144 13130 26145
rect 12814 26080 12820 26144
rect 12884 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13130 26144
rect 12814 26079 13130 26080
rect 18748 26144 19064 26145
rect 18748 26080 18754 26144
rect 18818 26080 18834 26144
rect 18898 26080 18914 26144
rect 18978 26080 18994 26144
rect 19058 26080 19064 26144
rect 18748 26079 19064 26080
rect 24682 26144 24998 26145
rect 24682 26080 24688 26144
rect 24752 26080 24768 26144
rect 24832 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 24998 26144
rect 25840 26120 26000 26150
rect 24682 26079 24998 26080
rect 1853 26074 1919 26077
rect 2262 26074 2268 26076
rect 1853 26072 2268 26074
rect 1853 26016 1858 26072
rect 1914 26016 2268 26072
rect 1853 26014 2268 26016
rect 1853 26011 1919 26014
rect 2262 26012 2268 26014
rect 2332 26012 2338 26076
rect 11881 26074 11947 26077
rect 12014 26074 12020 26076
rect 11881 26072 12020 26074
rect 11881 26016 11886 26072
rect 11942 26016 12020 26072
rect 11881 26014 12020 26016
rect 11881 26011 11947 26014
rect 12014 26012 12020 26014
rect 12084 26012 12090 26076
rect 0 25938 160 25968
rect 3509 25938 3575 25941
rect 0 25936 3575 25938
rect 0 25880 3514 25936
rect 3570 25880 3575 25936
rect 0 25878 3575 25880
rect 0 25848 160 25878
rect 3509 25875 3575 25878
rect 3969 25938 4035 25941
rect 8477 25938 8543 25941
rect 3969 25936 8543 25938
rect 3969 25880 3974 25936
rect 4030 25880 8482 25936
rect 8538 25880 8543 25936
rect 3969 25878 8543 25880
rect 3969 25875 4035 25878
rect 8477 25875 8543 25878
rect 10317 25938 10383 25941
rect 14089 25938 14155 25941
rect 10317 25936 14155 25938
rect 10317 25880 10322 25936
rect 10378 25880 14094 25936
rect 14150 25880 14155 25936
rect 10317 25878 14155 25880
rect 10317 25875 10383 25878
rect 14089 25875 14155 25878
rect 15929 25938 15995 25941
rect 16246 25938 16252 25940
rect 15929 25936 16252 25938
rect 15929 25880 15934 25936
rect 15990 25880 16252 25936
rect 15929 25878 16252 25880
rect 15929 25875 15995 25878
rect 16246 25876 16252 25878
rect 16316 25938 16322 25940
rect 16481 25938 16547 25941
rect 16316 25936 16547 25938
rect 16316 25880 16486 25936
rect 16542 25880 16547 25936
rect 16316 25878 16547 25880
rect 16316 25876 16322 25878
rect 16481 25875 16547 25878
rect 4061 25802 4127 25805
rect 2730 25800 4127 25802
rect 2730 25744 4066 25800
rect 4122 25744 4127 25800
rect 2730 25742 4127 25744
rect 0 25666 160 25696
rect 2730 25666 2790 25742
rect 4061 25739 4127 25742
rect 5993 25802 6059 25805
rect 8334 25802 8340 25804
rect 5993 25800 8340 25802
rect 5993 25744 5998 25800
rect 6054 25744 8340 25800
rect 5993 25742 8340 25744
rect 5993 25739 6059 25742
rect 8334 25740 8340 25742
rect 8404 25740 8410 25804
rect 0 25606 2790 25666
rect 0 25576 160 25606
rect 17166 25604 17172 25668
rect 17236 25666 17242 25668
rect 17585 25666 17651 25669
rect 17236 25664 17651 25666
rect 17236 25608 17590 25664
rect 17646 25608 17651 25664
rect 17236 25606 17651 25608
rect 17236 25604 17242 25606
rect 17585 25603 17651 25606
rect 24393 25666 24459 25669
rect 25840 25666 26000 25696
rect 24393 25664 26000 25666
rect 24393 25608 24398 25664
rect 24454 25608 26000 25664
rect 24393 25606 26000 25608
rect 24393 25603 24459 25606
rect 3913 25600 4229 25601
rect 3913 25536 3919 25600
rect 3983 25536 3999 25600
rect 4063 25536 4079 25600
rect 4143 25536 4159 25600
rect 4223 25536 4229 25600
rect 3913 25535 4229 25536
rect 9847 25600 10163 25601
rect 9847 25536 9853 25600
rect 9917 25536 9933 25600
rect 9997 25536 10013 25600
rect 10077 25536 10093 25600
rect 10157 25536 10163 25600
rect 9847 25535 10163 25536
rect 15781 25600 16097 25601
rect 15781 25536 15787 25600
rect 15851 25536 15867 25600
rect 15931 25536 15947 25600
rect 16011 25536 16027 25600
rect 16091 25536 16097 25600
rect 15781 25535 16097 25536
rect 21715 25600 22031 25601
rect 21715 25536 21721 25600
rect 21785 25536 21801 25600
rect 21865 25536 21881 25600
rect 21945 25536 21961 25600
rect 22025 25536 22031 25600
rect 25840 25576 26000 25606
rect 21715 25535 22031 25536
rect 2681 25532 2747 25533
rect 2630 25530 2636 25532
rect 2590 25470 2636 25530
rect 2700 25528 2747 25532
rect 2742 25472 2747 25528
rect 2630 25468 2636 25470
rect 2700 25468 2747 25472
rect 2681 25467 2747 25468
rect 0 25394 160 25424
rect 1301 25394 1367 25397
rect 0 25392 1367 25394
rect 0 25336 1306 25392
rect 1362 25336 1367 25392
rect 0 25334 1367 25336
rect 0 25304 160 25334
rect 1301 25331 1367 25334
rect 2957 25394 3023 25397
rect 6913 25394 6979 25397
rect 2957 25392 6979 25394
rect 2957 25336 2962 25392
rect 3018 25336 6918 25392
rect 6974 25336 6979 25392
rect 2957 25334 6979 25336
rect 2957 25331 3023 25334
rect 6913 25331 6979 25334
rect 7281 25394 7347 25397
rect 11789 25394 11855 25397
rect 7281 25392 11855 25394
rect 7281 25336 7286 25392
rect 7342 25336 11794 25392
rect 11850 25336 11855 25392
rect 7281 25334 11855 25336
rect 7281 25331 7347 25334
rect 11789 25331 11855 25334
rect 1853 25258 1919 25261
rect 15929 25258 15995 25261
rect 17585 25260 17651 25261
rect 1853 25256 15995 25258
rect 1853 25200 1858 25256
rect 1914 25200 15934 25256
rect 15990 25200 15995 25256
rect 1853 25198 15995 25200
rect 1853 25195 1919 25198
rect 15929 25195 15995 25198
rect 17534 25196 17540 25260
rect 17604 25258 17651 25260
rect 20621 25258 20687 25261
rect 17604 25256 17696 25258
rect 17646 25200 17696 25256
rect 17604 25198 17696 25200
rect 18462 25256 20687 25258
rect 18462 25200 20626 25256
rect 20682 25200 20687 25256
rect 18462 25198 20687 25200
rect 17604 25196 17651 25198
rect 17585 25195 17651 25196
rect 0 25122 160 25152
rect 1209 25122 1275 25125
rect 0 25120 1275 25122
rect 0 25064 1214 25120
rect 1270 25064 1275 25120
rect 0 25062 1275 25064
rect 0 25032 160 25062
rect 1209 25059 1275 25062
rect 11973 25122 12039 25125
rect 12198 25122 12204 25124
rect 11973 25120 12204 25122
rect 11973 25064 11978 25120
rect 12034 25064 12204 25120
rect 11973 25062 12204 25064
rect 11973 25059 12039 25062
rect 12198 25060 12204 25062
rect 12268 25060 12274 25124
rect 14222 25060 14228 25124
rect 14292 25122 14298 25124
rect 16113 25122 16179 25125
rect 18462 25122 18522 25198
rect 20621 25195 20687 25198
rect 14292 25120 16179 25122
rect 14292 25064 16118 25120
rect 16174 25064 16179 25120
rect 14292 25062 16179 25064
rect 14292 25060 14298 25062
rect 16113 25059 16179 25062
rect 16622 25062 18522 25122
rect 25129 25122 25195 25125
rect 25840 25122 26000 25152
rect 25129 25120 26000 25122
rect 25129 25064 25134 25120
rect 25190 25064 26000 25120
rect 25129 25062 26000 25064
rect 6880 25056 7196 25057
rect 6880 24992 6886 25056
rect 6950 24992 6966 25056
rect 7030 24992 7046 25056
rect 7110 24992 7126 25056
rect 7190 24992 7196 25056
rect 6880 24991 7196 24992
rect 12814 25056 13130 25057
rect 12814 24992 12820 25056
rect 12884 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13130 25056
rect 12814 24991 13130 24992
rect 2773 24986 2839 24989
rect 3734 24986 3740 24988
rect 2773 24984 3740 24986
rect 2773 24928 2778 24984
rect 2834 24928 3740 24984
rect 2773 24926 3740 24928
rect 2773 24923 2839 24926
rect 3734 24924 3740 24926
rect 3804 24986 3810 24988
rect 5165 24986 5231 24989
rect 3804 24984 5231 24986
rect 3804 24928 5170 24984
rect 5226 24928 5231 24984
rect 3804 24926 5231 24928
rect 3804 24924 3810 24926
rect 5165 24923 5231 24926
rect 15285 24986 15351 24989
rect 16622 24988 16682 25062
rect 25129 25059 25195 25062
rect 18748 25056 19064 25057
rect 18748 24992 18754 25056
rect 18818 24992 18834 25056
rect 18898 24992 18914 25056
rect 18978 24992 18994 25056
rect 19058 24992 19064 25056
rect 18748 24991 19064 24992
rect 24682 25056 24998 25057
rect 24682 24992 24688 25056
rect 24752 24992 24768 25056
rect 24832 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 24998 25056
rect 25840 25032 26000 25062
rect 24682 24991 24998 24992
rect 16614 24986 16620 24988
rect 15285 24984 16620 24986
rect 15285 24928 15290 24984
rect 15346 24928 16620 24984
rect 15285 24926 16620 24928
rect 15285 24923 15351 24926
rect 16614 24924 16620 24926
rect 16684 24924 16690 24988
rect 0 24850 160 24880
rect 2129 24850 2195 24853
rect 0 24848 2195 24850
rect 0 24792 2134 24848
rect 2190 24792 2195 24848
rect 0 24790 2195 24792
rect 0 24760 160 24790
rect 2129 24787 2195 24790
rect 2630 24788 2636 24852
rect 2700 24850 2706 24852
rect 3141 24850 3207 24853
rect 2700 24848 3207 24850
rect 2700 24792 3146 24848
rect 3202 24792 3207 24848
rect 2700 24790 3207 24792
rect 2700 24788 2706 24790
rect 3141 24787 3207 24790
rect 4153 24850 4219 24853
rect 22093 24850 22159 24853
rect 4153 24848 22159 24850
rect 4153 24792 4158 24848
rect 4214 24792 22098 24848
rect 22154 24792 22159 24848
rect 4153 24790 22159 24792
rect 4153 24787 4219 24790
rect 22093 24787 22159 24790
rect 22502 24788 22508 24852
rect 22572 24850 22578 24852
rect 22921 24850 22987 24853
rect 22572 24848 22987 24850
rect 22572 24792 22926 24848
rect 22982 24792 22987 24848
rect 22572 24790 22987 24792
rect 22572 24788 22578 24790
rect 22921 24787 22987 24790
rect 3693 24714 3759 24717
rect 4286 24714 4292 24716
rect 3693 24712 4292 24714
rect 3693 24656 3698 24712
rect 3754 24656 4292 24712
rect 3693 24654 4292 24656
rect 3693 24651 3759 24654
rect 4286 24652 4292 24654
rect 4356 24652 4362 24716
rect 13721 24714 13787 24717
rect 15377 24714 15443 24717
rect 13721 24712 15443 24714
rect 13721 24656 13726 24712
rect 13782 24656 15382 24712
rect 15438 24656 15443 24712
rect 13721 24654 15443 24656
rect 13721 24651 13787 24654
rect 15377 24651 15443 24654
rect 0 24578 160 24608
rect 1117 24578 1183 24581
rect 0 24576 1183 24578
rect 0 24520 1122 24576
rect 1178 24520 1183 24576
rect 0 24518 1183 24520
rect 0 24488 160 24518
rect 1117 24515 1183 24518
rect 15101 24578 15167 24581
rect 15326 24578 15332 24580
rect 15101 24576 15332 24578
rect 15101 24520 15106 24576
rect 15162 24520 15332 24576
rect 15101 24518 15332 24520
rect 15101 24515 15167 24518
rect 15326 24516 15332 24518
rect 15396 24516 15402 24580
rect 19609 24578 19675 24581
rect 19926 24578 19932 24580
rect 19609 24576 19932 24578
rect 19609 24520 19614 24576
rect 19670 24520 19932 24576
rect 19609 24518 19932 24520
rect 19609 24515 19675 24518
rect 19926 24516 19932 24518
rect 19996 24516 20002 24580
rect 24393 24578 24459 24581
rect 25840 24578 26000 24608
rect 24393 24576 26000 24578
rect 24393 24520 24398 24576
rect 24454 24520 26000 24576
rect 24393 24518 26000 24520
rect 24393 24515 24459 24518
rect 3913 24512 4229 24513
rect 3913 24448 3919 24512
rect 3983 24448 3999 24512
rect 4063 24448 4079 24512
rect 4143 24448 4159 24512
rect 4223 24448 4229 24512
rect 3913 24447 4229 24448
rect 9847 24512 10163 24513
rect 9847 24448 9853 24512
rect 9917 24448 9933 24512
rect 9997 24448 10013 24512
rect 10077 24448 10093 24512
rect 10157 24448 10163 24512
rect 9847 24447 10163 24448
rect 15781 24512 16097 24513
rect 15781 24448 15787 24512
rect 15851 24448 15867 24512
rect 15931 24448 15947 24512
rect 16011 24448 16027 24512
rect 16091 24448 16097 24512
rect 15781 24447 16097 24448
rect 21715 24512 22031 24513
rect 21715 24448 21721 24512
rect 21785 24448 21801 24512
rect 21865 24448 21881 24512
rect 21945 24448 21961 24512
rect 22025 24448 22031 24512
rect 25840 24488 26000 24518
rect 21715 24447 22031 24448
rect 0 24306 160 24336
rect 1669 24306 1735 24309
rect 0 24304 1735 24306
rect 0 24248 1674 24304
rect 1730 24248 1735 24304
rect 0 24246 1735 24248
rect 0 24216 160 24246
rect 1669 24243 1735 24246
rect 1853 24306 1919 24309
rect 4470 24306 4476 24308
rect 1853 24304 4476 24306
rect 1853 24248 1858 24304
rect 1914 24248 4476 24304
rect 1853 24246 4476 24248
rect 1853 24243 1919 24246
rect 4470 24244 4476 24246
rect 4540 24244 4546 24308
rect 8293 24306 8359 24309
rect 10593 24306 10659 24309
rect 11881 24306 11947 24309
rect 16430 24306 16436 24308
rect 8293 24304 10659 24306
rect 8293 24248 8298 24304
rect 8354 24248 10598 24304
rect 10654 24248 10659 24304
rect 8293 24246 10659 24248
rect 8293 24243 8359 24246
rect 10593 24243 10659 24246
rect 10734 24304 16436 24306
rect 10734 24248 11886 24304
rect 11942 24248 16436 24304
rect 10734 24246 16436 24248
rect 289 24170 355 24173
rect 10133 24170 10199 24173
rect 289 24168 10199 24170
rect 289 24112 294 24168
rect 350 24112 10138 24168
rect 10194 24112 10199 24168
rect 289 24110 10199 24112
rect 289 24107 355 24110
rect 10133 24107 10199 24110
rect 0 24034 160 24064
rect 1393 24034 1459 24037
rect 0 24032 1459 24034
rect 0 23976 1398 24032
rect 1454 23976 1459 24032
rect 0 23974 1459 23976
rect 0 23944 160 23974
rect 1393 23971 1459 23974
rect 2865 24034 2931 24037
rect 6126 24034 6132 24036
rect 2865 24032 6132 24034
rect 2865 23976 2870 24032
rect 2926 23976 6132 24032
rect 2865 23974 6132 23976
rect 2865 23971 2931 23974
rect 6126 23972 6132 23974
rect 6196 23972 6202 24036
rect 9581 24034 9647 24037
rect 10734 24034 10794 24246
rect 11881 24243 11947 24246
rect 16430 24244 16436 24246
rect 16500 24244 16506 24308
rect 22870 24244 22876 24308
rect 22940 24306 22946 24308
rect 23841 24306 23907 24309
rect 22940 24304 23907 24306
rect 22940 24248 23846 24304
rect 23902 24248 23907 24304
rect 22940 24246 23907 24248
rect 22940 24244 22946 24246
rect 23841 24243 23907 24246
rect 11329 24170 11395 24173
rect 12617 24170 12683 24173
rect 11329 24168 12683 24170
rect 11329 24112 11334 24168
rect 11390 24112 12622 24168
rect 12678 24112 12683 24168
rect 11329 24110 12683 24112
rect 11329 24107 11395 24110
rect 12617 24107 12683 24110
rect 15193 24170 15259 24173
rect 17309 24170 17375 24173
rect 15193 24168 17375 24170
rect 15193 24112 15198 24168
rect 15254 24112 17314 24168
rect 17370 24112 17375 24168
rect 15193 24110 17375 24112
rect 15193 24107 15259 24110
rect 17309 24107 17375 24110
rect 17718 24108 17724 24172
rect 17788 24170 17794 24172
rect 25497 24170 25563 24173
rect 17788 24168 25563 24170
rect 17788 24112 25502 24168
rect 25558 24112 25563 24168
rect 17788 24110 25563 24112
rect 17788 24108 17794 24110
rect 25497 24107 25563 24110
rect 9581 24032 10794 24034
rect 9581 23976 9586 24032
rect 9642 23976 10794 24032
rect 9581 23974 10794 23976
rect 25129 24034 25195 24037
rect 25840 24034 26000 24064
rect 25129 24032 26000 24034
rect 25129 23976 25134 24032
rect 25190 23976 26000 24032
rect 25129 23974 26000 23976
rect 9581 23971 9647 23974
rect 25129 23971 25195 23974
rect 6880 23968 7196 23969
rect 6880 23904 6886 23968
rect 6950 23904 6966 23968
rect 7030 23904 7046 23968
rect 7110 23904 7126 23968
rect 7190 23904 7196 23968
rect 6880 23903 7196 23904
rect 12814 23968 13130 23969
rect 12814 23904 12820 23968
rect 12884 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13130 23968
rect 12814 23903 13130 23904
rect 18748 23968 19064 23969
rect 18748 23904 18754 23968
rect 18818 23904 18834 23968
rect 18898 23904 18914 23968
rect 18978 23904 18994 23968
rect 19058 23904 19064 23968
rect 18748 23903 19064 23904
rect 24682 23968 24998 23969
rect 24682 23904 24688 23968
rect 24752 23904 24768 23968
rect 24832 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 24998 23968
rect 25840 23944 26000 23974
rect 24682 23903 24998 23904
rect 841 23898 907 23901
rect 4061 23898 4127 23901
rect 841 23896 4127 23898
rect 841 23840 846 23896
rect 902 23840 4066 23896
rect 4122 23840 4127 23896
rect 841 23838 4127 23840
rect 841 23835 907 23838
rect 4061 23835 4127 23838
rect 10726 23836 10732 23900
rect 10796 23898 10802 23900
rect 10869 23898 10935 23901
rect 10796 23896 10935 23898
rect 10796 23840 10874 23896
rect 10930 23840 10935 23896
rect 10796 23838 10935 23840
rect 10796 23836 10802 23838
rect 10869 23835 10935 23838
rect 0 23762 160 23792
rect 1301 23762 1367 23765
rect 0 23760 1367 23762
rect 0 23704 1306 23760
rect 1362 23704 1367 23760
rect 0 23702 1367 23704
rect 0 23672 160 23702
rect 1301 23699 1367 23702
rect 6085 23762 6151 23765
rect 21633 23762 21699 23765
rect 6085 23760 21699 23762
rect 6085 23704 6090 23760
rect 6146 23704 21638 23760
rect 21694 23704 21699 23760
rect 6085 23702 21699 23704
rect 6085 23699 6151 23702
rect 21633 23699 21699 23702
rect 381 23626 447 23629
rect 7414 23626 7420 23628
rect 381 23624 7420 23626
rect 381 23568 386 23624
rect 442 23568 7420 23624
rect 381 23566 7420 23568
rect 381 23563 447 23566
rect 7414 23564 7420 23566
rect 7484 23564 7490 23628
rect 8753 23626 8819 23629
rect 12065 23626 12131 23629
rect 8753 23624 12131 23626
rect 8753 23568 8758 23624
rect 8814 23568 12070 23624
rect 12126 23568 12131 23624
rect 8753 23566 12131 23568
rect 8753 23563 8819 23566
rect 12065 23563 12131 23566
rect 13261 23626 13327 23629
rect 13813 23626 13879 23629
rect 13261 23624 13879 23626
rect 13261 23568 13266 23624
rect 13322 23568 13818 23624
rect 13874 23568 13879 23624
rect 13261 23566 13879 23568
rect 13261 23563 13327 23566
rect 13813 23563 13879 23566
rect 19517 23626 19583 23629
rect 22686 23626 22692 23628
rect 19517 23624 22692 23626
rect 19517 23568 19522 23624
rect 19578 23568 22692 23624
rect 19517 23566 22692 23568
rect 19517 23563 19583 23566
rect 22686 23564 22692 23566
rect 22756 23564 22762 23628
rect 0 23490 160 23520
rect 749 23490 815 23493
rect 0 23488 815 23490
rect 0 23432 754 23488
rect 810 23432 815 23488
rect 0 23430 815 23432
rect 0 23400 160 23430
rect 749 23427 815 23430
rect 10869 23490 10935 23493
rect 14457 23490 14523 23493
rect 10869 23488 14523 23490
rect 10869 23432 10874 23488
rect 10930 23432 14462 23488
rect 14518 23432 14523 23488
rect 10869 23430 14523 23432
rect 10869 23427 10935 23430
rect 14457 23427 14523 23430
rect 22185 23490 22251 23493
rect 22686 23490 22692 23492
rect 22185 23488 22692 23490
rect 22185 23432 22190 23488
rect 22246 23432 22692 23488
rect 22185 23430 22692 23432
rect 22185 23427 22251 23430
rect 22686 23428 22692 23430
rect 22756 23428 22762 23492
rect 24393 23490 24459 23493
rect 25840 23490 26000 23520
rect 24393 23488 26000 23490
rect 24393 23432 24398 23488
rect 24454 23432 26000 23488
rect 24393 23430 26000 23432
rect 24393 23427 24459 23430
rect 3913 23424 4229 23425
rect 3913 23360 3919 23424
rect 3983 23360 3999 23424
rect 4063 23360 4079 23424
rect 4143 23360 4159 23424
rect 4223 23360 4229 23424
rect 3913 23359 4229 23360
rect 9847 23424 10163 23425
rect 9847 23360 9853 23424
rect 9917 23360 9933 23424
rect 9997 23360 10013 23424
rect 10077 23360 10093 23424
rect 10157 23360 10163 23424
rect 9847 23359 10163 23360
rect 15781 23424 16097 23425
rect 15781 23360 15787 23424
rect 15851 23360 15867 23424
rect 15931 23360 15947 23424
rect 16011 23360 16027 23424
rect 16091 23360 16097 23424
rect 15781 23359 16097 23360
rect 21715 23424 22031 23425
rect 21715 23360 21721 23424
rect 21785 23360 21801 23424
rect 21865 23360 21881 23424
rect 21945 23360 21961 23424
rect 22025 23360 22031 23424
rect 25840 23400 26000 23430
rect 21715 23359 22031 23360
rect 0 23218 160 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 160 23158
rect 1485 23155 1551 23158
rect 3049 23218 3115 23221
rect 3366 23218 3372 23220
rect 3049 23216 3372 23218
rect 3049 23160 3054 23216
rect 3110 23160 3372 23216
rect 3049 23158 3372 23160
rect 3049 23155 3115 23158
rect 3366 23156 3372 23158
rect 3436 23156 3442 23220
rect 3785 23218 3851 23221
rect 5574 23218 5580 23220
rect 3785 23216 5580 23218
rect 3785 23160 3790 23216
rect 3846 23160 5580 23216
rect 3785 23158 5580 23160
rect 3785 23155 3851 23158
rect 5574 23156 5580 23158
rect 5644 23218 5650 23220
rect 11513 23218 11579 23221
rect 5644 23216 11579 23218
rect 5644 23160 11518 23216
rect 11574 23160 11579 23216
rect 5644 23158 11579 23160
rect 5644 23156 5650 23158
rect 11513 23155 11579 23158
rect 1117 23082 1183 23085
rect 12617 23082 12683 23085
rect 1117 23080 12683 23082
rect 1117 23024 1122 23080
rect 1178 23024 12622 23080
rect 12678 23024 12683 23080
rect 1117 23022 12683 23024
rect 1117 23019 1183 23022
rect 12617 23019 12683 23022
rect 0 22946 160 22976
rect 1025 22946 1091 22949
rect 0 22944 1091 22946
rect 0 22888 1030 22944
rect 1086 22888 1091 22944
rect 0 22886 1091 22888
rect 0 22856 160 22886
rect 1025 22883 1091 22886
rect 2262 22884 2268 22948
rect 2332 22946 2338 22948
rect 2497 22946 2563 22949
rect 2332 22944 2563 22946
rect 2332 22888 2502 22944
rect 2558 22888 2563 22944
rect 2332 22886 2563 22888
rect 2332 22884 2338 22886
rect 2497 22883 2563 22886
rect 7925 22946 7991 22949
rect 11145 22946 11211 22949
rect 7925 22944 11211 22946
rect 7925 22888 7930 22944
rect 7986 22888 11150 22944
rect 11206 22888 11211 22944
rect 7925 22886 11211 22888
rect 7925 22883 7991 22886
rect 11145 22883 11211 22886
rect 25129 22946 25195 22949
rect 25840 22946 26000 22976
rect 25129 22944 26000 22946
rect 25129 22888 25134 22944
rect 25190 22888 26000 22944
rect 25129 22886 26000 22888
rect 25129 22883 25195 22886
rect 2500 22810 2560 22883
rect 6880 22880 7196 22881
rect 6880 22816 6886 22880
rect 6950 22816 6966 22880
rect 7030 22816 7046 22880
rect 7110 22816 7126 22880
rect 7190 22816 7196 22880
rect 6880 22815 7196 22816
rect 12814 22880 13130 22881
rect 12814 22816 12820 22880
rect 12884 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13130 22880
rect 12814 22815 13130 22816
rect 18748 22880 19064 22881
rect 18748 22816 18754 22880
rect 18818 22816 18834 22880
rect 18898 22816 18914 22880
rect 18978 22816 18994 22880
rect 19058 22816 19064 22880
rect 18748 22815 19064 22816
rect 24682 22880 24998 22881
rect 24682 22816 24688 22880
rect 24752 22816 24768 22880
rect 24832 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 24998 22880
rect 25840 22856 26000 22886
rect 24682 22815 24998 22816
rect 5390 22810 5396 22812
rect 2500 22750 5396 22810
rect 5390 22748 5396 22750
rect 5460 22810 5466 22812
rect 6545 22810 6611 22813
rect 5460 22808 6611 22810
rect 5460 22752 6550 22808
rect 6606 22752 6611 22808
rect 5460 22750 6611 22752
rect 5460 22748 5466 22750
rect 6545 22747 6611 22750
rect 10041 22810 10107 22813
rect 11789 22810 11855 22813
rect 10041 22808 11855 22810
rect 10041 22752 10046 22808
rect 10102 22752 11794 22808
rect 11850 22752 11855 22808
rect 10041 22750 11855 22752
rect 10041 22747 10107 22750
rect 11789 22747 11855 22750
rect 0 22674 160 22704
rect 1301 22674 1367 22677
rect 0 22672 1367 22674
rect 0 22616 1306 22672
rect 1362 22616 1367 22672
rect 0 22614 1367 22616
rect 0 22584 160 22614
rect 1301 22611 1367 22614
rect 9581 22674 9647 22677
rect 14273 22674 14339 22677
rect 9581 22672 14339 22674
rect 9581 22616 9586 22672
rect 9642 22616 14278 22672
rect 14334 22616 14339 22672
rect 9581 22614 14339 22616
rect 9581 22611 9647 22614
rect 14273 22611 14339 22614
rect 11329 22538 11395 22541
rect 11462 22538 11468 22540
rect 11329 22536 11468 22538
rect 11329 22480 11334 22536
rect 11390 22480 11468 22536
rect 11329 22478 11468 22480
rect 11329 22475 11395 22478
rect 11462 22476 11468 22478
rect 11532 22476 11538 22540
rect 21633 22538 21699 22541
rect 22461 22538 22527 22541
rect 21633 22536 22527 22538
rect 21633 22480 21638 22536
rect 21694 22480 22466 22536
rect 22522 22480 22527 22536
rect 21633 22478 22527 22480
rect 21633 22475 21699 22478
rect 22461 22475 22527 22478
rect 0 22402 160 22432
rect 1485 22402 1551 22405
rect 0 22400 1551 22402
rect 0 22344 1490 22400
rect 1546 22344 1551 22400
rect 0 22342 1551 22344
rect 0 22312 160 22342
rect 1485 22339 1551 22342
rect 14549 22400 14615 22405
rect 14549 22344 14554 22400
rect 14610 22344 14615 22400
rect 14549 22339 14615 22344
rect 24485 22402 24551 22405
rect 25840 22402 26000 22432
rect 24485 22400 26000 22402
rect 24485 22344 24490 22400
rect 24546 22344 26000 22400
rect 24485 22342 26000 22344
rect 24485 22339 24551 22342
rect 3913 22336 4229 22337
rect 3913 22272 3919 22336
rect 3983 22272 3999 22336
rect 4063 22272 4079 22336
rect 4143 22272 4159 22336
rect 4223 22272 4229 22336
rect 3913 22271 4229 22272
rect 9847 22336 10163 22337
rect 9847 22272 9853 22336
rect 9917 22272 9933 22336
rect 9997 22272 10013 22336
rect 10077 22272 10093 22336
rect 10157 22272 10163 22336
rect 9847 22271 10163 22272
rect 0 22130 160 22160
rect 3233 22130 3299 22133
rect 0 22128 3299 22130
rect 0 22072 3238 22128
rect 3294 22072 3299 22128
rect 0 22070 3299 22072
rect 14552 22130 14612 22339
rect 15781 22336 16097 22337
rect 15781 22272 15787 22336
rect 15851 22272 15867 22336
rect 15931 22272 15947 22336
rect 16011 22272 16027 22336
rect 16091 22272 16097 22336
rect 15781 22271 16097 22272
rect 21715 22336 22031 22337
rect 21715 22272 21721 22336
rect 21785 22272 21801 22336
rect 21865 22272 21881 22336
rect 21945 22272 21961 22336
rect 22025 22272 22031 22336
rect 25840 22312 26000 22342
rect 21715 22271 22031 22272
rect 15745 22130 15811 22133
rect 14552 22128 15811 22130
rect 14552 22072 15750 22128
rect 15806 22072 15811 22128
rect 14552 22070 15811 22072
rect 0 22040 160 22070
rect 3233 22067 3299 22070
rect 15745 22067 15811 22070
rect 18413 22130 18479 22133
rect 20989 22130 21055 22133
rect 21357 22130 21423 22133
rect 18413 22128 18522 22130
rect 18413 22072 18418 22128
rect 18474 22072 18522 22128
rect 18413 22067 18522 22072
rect 20989 22128 21423 22130
rect 20989 22072 20994 22128
rect 21050 22072 21362 22128
rect 21418 22072 21423 22128
rect 20989 22070 21423 22072
rect 20989 22067 21055 22070
rect 21357 22067 21423 22070
rect 4153 21994 4219 21997
rect 9765 21994 9831 21997
rect 4153 21992 9831 21994
rect 4153 21936 4158 21992
rect 4214 21936 9770 21992
rect 9826 21936 9831 21992
rect 4153 21934 9831 21936
rect 4153 21931 4219 21934
rect 9765 21931 9831 21934
rect 11053 21994 11119 21997
rect 13854 21994 13860 21996
rect 11053 21992 13860 21994
rect 11053 21936 11058 21992
rect 11114 21936 13860 21992
rect 11053 21934 13860 21936
rect 11053 21931 11119 21934
rect 13854 21932 13860 21934
rect 13924 21932 13930 21996
rect 0 21858 160 21888
rect 18462 21861 18522 22067
rect 1301 21858 1367 21861
rect 0 21856 1367 21858
rect 0 21800 1306 21856
rect 1362 21800 1367 21856
rect 0 21798 1367 21800
rect 0 21768 160 21798
rect 1301 21795 1367 21798
rect 4613 21858 4679 21861
rect 5625 21858 5691 21861
rect 4613 21856 5691 21858
rect 4613 21800 4618 21856
rect 4674 21800 5630 21856
rect 5686 21800 5691 21856
rect 4613 21798 5691 21800
rect 4613 21795 4679 21798
rect 5625 21795 5691 21798
rect 16849 21858 16915 21861
rect 17166 21858 17172 21860
rect 16849 21856 17172 21858
rect 16849 21800 16854 21856
rect 16910 21800 17172 21856
rect 16849 21798 17172 21800
rect 16849 21795 16915 21798
rect 17166 21796 17172 21798
rect 17236 21796 17242 21860
rect 18413 21856 18522 21861
rect 18413 21800 18418 21856
rect 18474 21800 18522 21856
rect 18413 21798 18522 21800
rect 25129 21858 25195 21861
rect 25840 21858 26000 21888
rect 25129 21856 26000 21858
rect 25129 21800 25134 21856
rect 25190 21800 26000 21856
rect 25129 21798 26000 21800
rect 18413 21795 18479 21798
rect 25129 21795 25195 21798
rect 6880 21792 7196 21793
rect 6880 21728 6886 21792
rect 6950 21728 6966 21792
rect 7030 21728 7046 21792
rect 7110 21728 7126 21792
rect 7190 21728 7196 21792
rect 6880 21727 7196 21728
rect 12814 21792 13130 21793
rect 12814 21728 12820 21792
rect 12884 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13130 21792
rect 12814 21727 13130 21728
rect 18748 21792 19064 21793
rect 18748 21728 18754 21792
rect 18818 21728 18834 21792
rect 18898 21728 18914 21792
rect 18978 21728 18994 21792
rect 19058 21728 19064 21792
rect 18748 21727 19064 21728
rect 24682 21792 24998 21793
rect 24682 21728 24688 21792
rect 24752 21728 24768 21792
rect 24832 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 24998 21792
rect 25840 21768 26000 21798
rect 24682 21727 24998 21728
rect 9121 21722 9187 21725
rect 9581 21722 9647 21725
rect 9121 21720 9647 21722
rect 9121 21664 9126 21720
rect 9182 21664 9586 21720
rect 9642 21664 9647 21720
rect 9121 21662 9647 21664
rect 9121 21659 9187 21662
rect 9581 21659 9647 21662
rect 17953 21722 18019 21725
rect 18321 21722 18387 21725
rect 17953 21720 18387 21722
rect 17953 21664 17958 21720
rect 18014 21664 18326 21720
rect 18382 21664 18387 21720
rect 17953 21662 18387 21664
rect 17953 21659 18019 21662
rect 18321 21659 18387 21662
rect 0 21586 160 21616
rect 1209 21586 1275 21589
rect 0 21584 1275 21586
rect 0 21528 1214 21584
rect 1270 21528 1275 21584
rect 0 21526 1275 21528
rect 0 21496 160 21526
rect 1209 21523 1275 21526
rect 1761 21586 1827 21589
rect 7649 21586 7715 21589
rect 10869 21586 10935 21589
rect 16481 21586 16547 21589
rect 1761 21584 7715 21586
rect 1761 21528 1766 21584
rect 1822 21528 7654 21584
rect 7710 21528 7715 21584
rect 1761 21526 7715 21528
rect 1761 21523 1827 21526
rect 7649 21523 7715 21526
rect 7790 21584 16547 21586
rect 7790 21528 10874 21584
rect 10930 21528 16486 21584
rect 16542 21528 16547 21584
rect 7790 21526 16547 21528
rect 5022 21450 5028 21452
rect 3742 21390 5028 21450
rect 0 21314 160 21344
rect 1209 21314 1275 21317
rect 0 21312 1275 21314
rect 0 21256 1214 21312
rect 1270 21256 1275 21312
rect 0 21254 1275 21256
rect 0 21224 160 21254
rect 1209 21251 1275 21254
rect 0 21042 160 21072
rect 1301 21042 1367 21045
rect 0 21040 1367 21042
rect 0 20984 1306 21040
rect 1362 20984 1367 21040
rect 0 20982 1367 20984
rect 0 20952 160 20982
rect 1301 20979 1367 20982
rect 2313 21042 2379 21045
rect 3742 21042 3802 21390
rect 5022 21388 5028 21390
rect 5092 21450 5098 21452
rect 7790 21450 7850 21526
rect 10869 21523 10935 21526
rect 16481 21523 16547 21526
rect 17534 21524 17540 21588
rect 17604 21586 17610 21588
rect 17769 21586 17835 21589
rect 17604 21584 17835 21586
rect 17604 21528 17774 21584
rect 17830 21528 17835 21584
rect 17604 21526 17835 21528
rect 17604 21524 17610 21526
rect 17769 21523 17835 21526
rect 5092 21390 7850 21450
rect 8201 21450 8267 21453
rect 11697 21450 11763 21453
rect 16481 21450 16547 21453
rect 8201 21448 10426 21450
rect 8201 21392 8206 21448
rect 8262 21392 10426 21448
rect 8201 21390 10426 21392
rect 5092 21388 5098 21390
rect 8201 21387 8267 21390
rect 9254 21252 9260 21316
rect 9324 21314 9330 21316
rect 9397 21314 9463 21317
rect 9324 21312 9463 21314
rect 9324 21256 9402 21312
rect 9458 21256 9463 21312
rect 9324 21254 9463 21256
rect 10366 21314 10426 21390
rect 11697 21448 16547 21450
rect 11697 21392 11702 21448
rect 11758 21392 16486 21448
rect 16542 21392 16547 21448
rect 11697 21390 16547 21392
rect 11697 21387 11763 21390
rect 16481 21387 16547 21390
rect 16614 21388 16620 21452
rect 16684 21450 16690 21452
rect 18137 21450 18203 21453
rect 16684 21448 18203 21450
rect 16684 21392 18142 21448
rect 18198 21392 18203 21448
rect 16684 21390 18203 21392
rect 16684 21388 16690 21390
rect 18137 21387 18203 21390
rect 10366 21254 12450 21314
rect 9324 21252 9330 21254
rect 9397 21251 9463 21254
rect 3913 21248 4229 21249
rect 3913 21184 3919 21248
rect 3983 21184 3999 21248
rect 4063 21184 4079 21248
rect 4143 21184 4159 21248
rect 4223 21184 4229 21248
rect 3913 21183 4229 21184
rect 9847 21248 10163 21249
rect 9847 21184 9853 21248
rect 9917 21184 9933 21248
rect 9997 21184 10013 21248
rect 10077 21184 10093 21248
rect 10157 21184 10163 21248
rect 9847 21183 10163 21184
rect 3969 21042 4035 21045
rect 2313 21040 4035 21042
rect 2313 20984 2318 21040
rect 2374 20984 3974 21040
rect 4030 20984 4035 21040
rect 2313 20982 4035 20984
rect 2313 20979 2379 20982
rect 3969 20979 4035 20982
rect 4337 21042 4403 21045
rect 4705 21042 4771 21045
rect 9857 21042 9923 21045
rect 4337 21040 9923 21042
rect 4337 20984 4342 21040
rect 4398 20984 4710 21040
rect 4766 20984 9862 21040
rect 9918 20984 9923 21040
rect 4337 20982 9923 20984
rect 4337 20979 4403 20982
rect 4705 20979 4771 20982
rect 9857 20979 9923 20982
rect 10133 21042 10199 21045
rect 11789 21042 11855 21045
rect 10133 21040 11855 21042
rect 10133 20984 10138 21040
rect 10194 20984 11794 21040
rect 11850 20984 11855 21040
rect 10133 20982 11855 20984
rect 12390 21042 12450 21254
rect 16430 21252 16436 21316
rect 16500 21314 16506 21316
rect 20253 21314 20319 21317
rect 16500 21312 20319 21314
rect 16500 21256 20258 21312
rect 20314 21256 20319 21312
rect 16500 21254 20319 21256
rect 16500 21252 16506 21254
rect 20253 21251 20319 21254
rect 23841 21314 23907 21317
rect 25840 21314 26000 21344
rect 23841 21312 26000 21314
rect 23841 21256 23846 21312
rect 23902 21256 26000 21312
rect 23841 21254 26000 21256
rect 23841 21251 23907 21254
rect 15781 21248 16097 21249
rect 15781 21184 15787 21248
rect 15851 21184 15867 21248
rect 15931 21184 15947 21248
rect 16011 21184 16027 21248
rect 16091 21184 16097 21248
rect 15781 21183 16097 21184
rect 21715 21248 22031 21249
rect 21715 21184 21721 21248
rect 21785 21184 21801 21248
rect 21865 21184 21881 21248
rect 21945 21184 21961 21248
rect 22025 21184 22031 21248
rect 25840 21224 26000 21254
rect 21715 21183 22031 21184
rect 17309 21180 17375 21181
rect 17309 21176 17356 21180
rect 17420 21178 17426 21180
rect 19149 21178 19215 21181
rect 19977 21180 20043 21181
rect 19558 21178 19564 21180
rect 17309 21120 17314 21176
rect 17309 21116 17356 21120
rect 17420 21118 17466 21178
rect 19149 21176 19564 21178
rect 19149 21120 19154 21176
rect 19210 21120 19564 21176
rect 19149 21118 19564 21120
rect 17420 21116 17426 21118
rect 17309 21115 17375 21116
rect 19149 21115 19215 21118
rect 19558 21116 19564 21118
rect 19628 21116 19634 21180
rect 19926 21116 19932 21180
rect 19996 21178 20043 21180
rect 19996 21176 20088 21178
rect 20038 21120 20088 21176
rect 19996 21118 20088 21120
rect 19996 21116 20043 21118
rect 19977 21115 20043 21116
rect 20805 21042 20871 21045
rect 12390 21040 20871 21042
rect 12390 20984 20810 21040
rect 20866 20984 20871 21040
rect 12390 20982 20871 20984
rect 10133 20979 10199 20982
rect 11789 20979 11855 20982
rect 20805 20979 20871 20982
rect 6678 20844 6684 20908
rect 6748 20906 6754 20908
rect 9622 20906 9628 20908
rect 6748 20846 9628 20906
rect 6748 20844 6754 20846
rect 9622 20844 9628 20846
rect 9692 20844 9698 20908
rect 12566 20844 12572 20908
rect 12636 20906 12642 20908
rect 13169 20906 13235 20909
rect 12636 20904 13235 20906
rect 12636 20848 13174 20904
rect 13230 20848 13235 20904
rect 12636 20846 13235 20848
rect 12636 20844 12642 20846
rect 13169 20843 13235 20846
rect 0 20770 160 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 160 20710
rect 1301 20707 1367 20710
rect 2446 20708 2452 20772
rect 2516 20770 2522 20772
rect 3182 20770 3188 20772
rect 2516 20710 3188 20770
rect 2516 20708 2522 20710
rect 3182 20708 3188 20710
rect 3252 20708 3258 20772
rect 6310 20708 6316 20772
rect 6380 20770 6386 20772
rect 6545 20770 6611 20773
rect 6380 20768 6611 20770
rect 6380 20712 6550 20768
rect 6606 20712 6611 20768
rect 6380 20710 6611 20712
rect 6380 20708 6386 20710
rect 6545 20707 6611 20710
rect 7557 20772 7623 20773
rect 7557 20768 7604 20772
rect 7668 20770 7674 20772
rect 8017 20770 8083 20773
rect 12617 20770 12683 20773
rect 19333 20772 19399 20773
rect 19333 20770 19380 20772
rect 7557 20712 7562 20768
rect 7557 20708 7604 20712
rect 7668 20710 7714 20770
rect 8017 20768 12683 20770
rect 8017 20712 8022 20768
rect 8078 20712 12622 20768
rect 12678 20712 12683 20768
rect 8017 20710 12683 20712
rect 19288 20768 19380 20770
rect 19288 20712 19338 20768
rect 19288 20710 19380 20712
rect 7668 20708 7674 20710
rect 7557 20707 7623 20708
rect 8017 20707 8083 20710
rect 12617 20707 12683 20710
rect 19333 20708 19380 20710
rect 19444 20708 19450 20772
rect 25129 20770 25195 20773
rect 25840 20770 26000 20800
rect 25129 20768 26000 20770
rect 25129 20712 25134 20768
rect 25190 20712 26000 20768
rect 25129 20710 26000 20712
rect 19333 20707 19399 20708
rect 25129 20707 25195 20710
rect 6880 20704 7196 20705
rect 6880 20640 6886 20704
rect 6950 20640 6966 20704
rect 7030 20640 7046 20704
rect 7110 20640 7126 20704
rect 7190 20640 7196 20704
rect 6880 20639 7196 20640
rect 12814 20704 13130 20705
rect 12814 20640 12820 20704
rect 12884 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13130 20704
rect 12814 20639 13130 20640
rect 18748 20704 19064 20705
rect 18748 20640 18754 20704
rect 18818 20640 18834 20704
rect 18898 20640 18914 20704
rect 18978 20640 18994 20704
rect 19058 20640 19064 20704
rect 18748 20639 19064 20640
rect 24682 20704 24998 20705
rect 24682 20640 24688 20704
rect 24752 20640 24768 20704
rect 24832 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 24998 20704
rect 25840 20680 26000 20710
rect 24682 20639 24998 20640
rect 2037 20634 2103 20637
rect 6361 20634 6427 20637
rect 2037 20632 6427 20634
rect 2037 20576 2042 20632
rect 2098 20576 6366 20632
rect 6422 20576 6427 20632
rect 2037 20574 6427 20576
rect 2037 20571 2103 20574
rect 6361 20571 6427 20574
rect 0 20498 160 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 160 20438
rect 1393 20435 1459 20438
rect 2773 20498 2839 20501
rect 3734 20498 3740 20500
rect 2773 20496 3740 20498
rect 2773 20440 2778 20496
rect 2834 20440 3740 20496
rect 2773 20438 3740 20440
rect 2773 20435 2839 20438
rect 3734 20436 3740 20438
rect 3804 20498 3810 20500
rect 3877 20498 3943 20501
rect 3804 20496 3943 20498
rect 3804 20440 3882 20496
rect 3938 20440 3943 20496
rect 3804 20438 3943 20440
rect 3804 20436 3810 20438
rect 3877 20435 3943 20438
rect 9949 20498 10015 20501
rect 13261 20498 13327 20501
rect 9949 20496 13327 20498
rect 9949 20440 9954 20496
rect 10010 20440 13266 20496
rect 13322 20440 13327 20496
rect 9949 20438 13327 20440
rect 9949 20435 10015 20438
rect 13261 20435 13327 20438
rect 841 20362 907 20365
rect 11237 20362 11303 20365
rect 841 20360 11303 20362
rect 841 20304 846 20360
rect 902 20304 11242 20360
rect 11298 20304 11303 20360
rect 841 20302 11303 20304
rect 841 20299 907 20302
rect 11237 20299 11303 20302
rect 0 20226 160 20256
rect 749 20226 815 20229
rect 0 20224 815 20226
rect 0 20168 754 20224
rect 810 20168 815 20224
rect 0 20166 815 20168
rect 0 20136 160 20166
rect 749 20163 815 20166
rect 6361 20226 6427 20229
rect 8845 20226 8911 20229
rect 6361 20224 8911 20226
rect 6361 20168 6366 20224
rect 6422 20168 8850 20224
rect 8906 20168 8911 20224
rect 6361 20166 8911 20168
rect 6361 20163 6427 20166
rect 8845 20163 8911 20166
rect 24025 20226 24091 20229
rect 25840 20226 26000 20256
rect 24025 20224 26000 20226
rect 24025 20168 24030 20224
rect 24086 20168 26000 20224
rect 24025 20166 26000 20168
rect 24025 20163 24091 20166
rect 3913 20160 4229 20161
rect 3913 20096 3919 20160
rect 3983 20096 3999 20160
rect 4063 20096 4079 20160
rect 4143 20096 4159 20160
rect 4223 20096 4229 20160
rect 3913 20095 4229 20096
rect 9847 20160 10163 20161
rect 9847 20096 9853 20160
rect 9917 20096 9933 20160
rect 9997 20096 10013 20160
rect 10077 20096 10093 20160
rect 10157 20096 10163 20160
rect 9847 20095 10163 20096
rect 15781 20160 16097 20161
rect 15781 20096 15787 20160
rect 15851 20096 15867 20160
rect 15931 20096 15947 20160
rect 16011 20096 16027 20160
rect 16091 20096 16097 20160
rect 15781 20095 16097 20096
rect 21715 20160 22031 20161
rect 21715 20096 21721 20160
rect 21785 20096 21801 20160
rect 21865 20096 21881 20160
rect 21945 20096 21961 20160
rect 22025 20096 22031 20160
rect 25840 20136 26000 20166
rect 21715 20095 22031 20096
rect 0 19954 160 19984
rect 841 19954 907 19957
rect 0 19952 907 19954
rect 0 19896 846 19952
rect 902 19896 907 19952
rect 0 19894 907 19896
rect 0 19864 160 19894
rect 841 19891 907 19894
rect 2221 19954 2287 19957
rect 2630 19954 2636 19956
rect 2221 19952 2636 19954
rect 2221 19896 2226 19952
rect 2282 19896 2636 19952
rect 2221 19894 2636 19896
rect 2221 19891 2287 19894
rect 2630 19892 2636 19894
rect 2700 19954 2706 19956
rect 8201 19954 8267 19957
rect 9857 19954 9923 19957
rect 2700 19952 9923 19954
rect 2700 19896 8206 19952
rect 8262 19896 9862 19952
rect 9918 19896 9923 19952
rect 2700 19894 9923 19896
rect 2700 19892 2706 19894
rect 8201 19891 8267 19894
rect 9857 19891 9923 19894
rect 12525 19954 12591 19957
rect 14958 19954 14964 19956
rect 12525 19952 14964 19954
rect 12525 19896 12530 19952
rect 12586 19896 14964 19952
rect 12525 19894 14964 19896
rect 12525 19891 12591 19894
rect 14958 19892 14964 19894
rect 15028 19892 15034 19956
rect 1577 19818 1643 19821
rect 2865 19818 2931 19821
rect 6821 19818 6887 19821
rect 1577 19816 6887 19818
rect 1577 19760 1582 19816
rect 1638 19760 2870 19816
rect 2926 19760 6826 19816
rect 6882 19760 6887 19816
rect 1577 19758 6887 19760
rect 1577 19755 1643 19758
rect 2865 19755 2931 19758
rect 6821 19755 6887 19758
rect 7465 19818 7531 19821
rect 8150 19818 8156 19820
rect 7465 19816 8156 19818
rect 7465 19760 7470 19816
rect 7526 19760 8156 19816
rect 7465 19758 8156 19760
rect 7465 19755 7531 19758
rect 8150 19756 8156 19758
rect 8220 19756 8226 19820
rect 10593 19818 10659 19821
rect 10726 19818 10732 19820
rect 10593 19816 10732 19818
rect 10593 19760 10598 19816
rect 10654 19760 10732 19816
rect 10593 19758 10732 19760
rect 10593 19755 10659 19758
rect 10726 19756 10732 19758
rect 10796 19756 10802 19820
rect 13537 19818 13603 19821
rect 13670 19818 13676 19820
rect 13537 19816 13676 19818
rect 13537 19760 13542 19816
rect 13598 19760 13676 19816
rect 13537 19758 13676 19760
rect 13537 19755 13603 19758
rect 13670 19756 13676 19758
rect 13740 19756 13746 19820
rect 0 19682 160 19712
rect 1301 19682 1367 19685
rect 0 19680 1367 19682
rect 0 19624 1306 19680
rect 1362 19624 1367 19680
rect 0 19622 1367 19624
rect 0 19592 160 19622
rect 1301 19619 1367 19622
rect 21214 19620 21220 19684
rect 21284 19620 21290 19684
rect 25313 19682 25379 19685
rect 25840 19682 26000 19712
rect 25313 19680 26000 19682
rect 25313 19624 25318 19680
rect 25374 19624 26000 19680
rect 25313 19622 26000 19624
rect 6880 19616 7196 19617
rect 6880 19552 6886 19616
rect 6950 19552 6966 19616
rect 7030 19552 7046 19616
rect 7110 19552 7126 19616
rect 7190 19552 7196 19616
rect 6880 19551 7196 19552
rect 12814 19616 13130 19617
rect 12814 19552 12820 19616
rect 12884 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13130 19616
rect 12814 19551 13130 19552
rect 18748 19616 19064 19617
rect 18748 19552 18754 19616
rect 18818 19552 18834 19616
rect 18898 19552 18914 19616
rect 18978 19552 18994 19616
rect 19058 19552 19064 19616
rect 18748 19551 19064 19552
rect 15142 19484 15148 19548
rect 15212 19546 15218 19548
rect 15212 19486 17050 19546
rect 15212 19484 15218 19486
rect 0 19410 160 19440
rect 1761 19410 1827 19413
rect 0 19408 1827 19410
rect 0 19352 1766 19408
rect 1822 19352 1827 19408
rect 0 19350 1827 19352
rect 0 19320 160 19350
rect 1761 19347 1827 19350
rect 7189 19410 7255 19413
rect 9254 19410 9260 19412
rect 7189 19408 9260 19410
rect 7189 19352 7194 19408
rect 7250 19352 9260 19408
rect 7189 19350 9260 19352
rect 7189 19347 7255 19350
rect 9254 19348 9260 19350
rect 9324 19410 9330 19412
rect 9489 19410 9555 19413
rect 9324 19408 9555 19410
rect 9324 19352 9494 19408
rect 9550 19352 9555 19408
rect 9324 19350 9555 19352
rect 9324 19348 9330 19350
rect 9489 19347 9555 19350
rect 10225 19410 10291 19413
rect 11421 19410 11487 19413
rect 10225 19408 11487 19410
rect 10225 19352 10230 19408
rect 10286 19352 11426 19408
rect 11482 19352 11487 19408
rect 10225 19350 11487 19352
rect 10225 19347 10291 19350
rect 11421 19347 11487 19350
rect 12341 19410 12407 19413
rect 13905 19410 13971 19413
rect 12341 19408 13971 19410
rect 12341 19352 12346 19408
rect 12402 19352 13910 19408
rect 13966 19352 13971 19408
rect 12341 19350 13971 19352
rect 12341 19347 12407 19350
rect 13905 19347 13971 19350
rect 16205 19410 16271 19413
rect 16798 19410 16804 19412
rect 16205 19408 16804 19410
rect 16205 19352 16210 19408
rect 16266 19352 16804 19408
rect 16205 19350 16804 19352
rect 16205 19347 16271 19350
rect 16798 19348 16804 19350
rect 16868 19348 16874 19412
rect 16990 19410 17050 19486
rect 19425 19410 19491 19413
rect 16990 19408 19491 19410
rect 16990 19352 19430 19408
rect 19486 19352 19491 19408
rect 16990 19350 19491 19352
rect 19425 19347 19491 19350
rect 21081 19410 21147 19413
rect 21222 19410 21282 19620
rect 25313 19619 25379 19622
rect 24682 19616 24998 19617
rect 24682 19552 24688 19616
rect 24752 19552 24768 19616
rect 24832 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 24998 19616
rect 25840 19592 26000 19622
rect 24682 19551 24998 19552
rect 21081 19408 21282 19410
rect 21081 19352 21086 19408
rect 21142 19352 21282 19408
rect 21081 19350 21282 19352
rect 21081 19347 21147 19350
rect 3785 19274 3851 19277
rect 4286 19274 4292 19276
rect 3785 19272 4292 19274
rect 3785 19216 3790 19272
rect 3846 19216 4292 19272
rect 3785 19214 4292 19216
rect 3785 19211 3851 19214
rect 4286 19212 4292 19214
rect 4356 19212 4362 19276
rect 9622 19212 9628 19276
rect 9692 19274 9698 19276
rect 10409 19274 10475 19277
rect 9692 19272 10475 19274
rect 9692 19216 10414 19272
rect 10470 19216 10475 19272
rect 9692 19214 10475 19216
rect 9692 19212 9698 19214
rect 10409 19211 10475 19214
rect 11421 19274 11487 19277
rect 16982 19274 16988 19276
rect 11421 19272 16988 19274
rect 11421 19216 11426 19272
rect 11482 19216 16988 19272
rect 11421 19214 16988 19216
rect 11421 19211 11487 19214
rect 16982 19212 16988 19214
rect 17052 19212 17058 19276
rect 0 19138 160 19168
rect 3325 19138 3391 19141
rect 0 19136 3391 19138
rect 0 19080 3330 19136
rect 3386 19080 3391 19136
rect 0 19078 3391 19080
rect 0 19048 160 19078
rect 3325 19075 3391 19078
rect 23841 19138 23907 19141
rect 25840 19138 26000 19168
rect 23841 19136 26000 19138
rect 23841 19080 23846 19136
rect 23902 19080 26000 19136
rect 23841 19078 26000 19080
rect 23841 19075 23907 19078
rect 3913 19072 4229 19073
rect 3913 19008 3919 19072
rect 3983 19008 3999 19072
rect 4063 19008 4079 19072
rect 4143 19008 4159 19072
rect 4223 19008 4229 19072
rect 3913 19007 4229 19008
rect 9847 19072 10163 19073
rect 9847 19008 9853 19072
rect 9917 19008 9933 19072
rect 9997 19008 10013 19072
rect 10077 19008 10093 19072
rect 10157 19008 10163 19072
rect 9847 19007 10163 19008
rect 15781 19072 16097 19073
rect 15781 19008 15787 19072
rect 15851 19008 15867 19072
rect 15931 19008 15947 19072
rect 16011 19008 16027 19072
rect 16091 19008 16097 19072
rect 15781 19007 16097 19008
rect 21715 19072 22031 19073
rect 21715 19008 21721 19072
rect 21785 19008 21801 19072
rect 21865 19008 21881 19072
rect 21945 19008 21961 19072
rect 22025 19008 22031 19072
rect 25840 19048 26000 19078
rect 21715 19007 22031 19008
rect 6453 19002 6519 19005
rect 8937 19002 9003 19005
rect 6453 19000 9003 19002
rect 6453 18944 6458 19000
rect 6514 18944 8942 19000
rect 8998 18944 9003 19000
rect 6453 18942 9003 18944
rect 6453 18939 6519 18942
rect 8937 18939 9003 18942
rect 0 18866 160 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 160 18806
rect 1393 18803 1459 18806
rect 2078 18804 2084 18868
rect 2148 18866 2154 18868
rect 3969 18866 4035 18869
rect 2148 18864 4035 18866
rect 2148 18808 3974 18864
rect 4030 18808 4035 18864
rect 2148 18806 4035 18808
rect 2148 18804 2154 18806
rect 3969 18803 4035 18806
rect 8385 18866 8451 18869
rect 17166 18866 17172 18868
rect 8385 18864 17172 18866
rect 8385 18808 8390 18864
rect 8446 18808 17172 18864
rect 8385 18806 17172 18808
rect 8385 18803 8451 18806
rect 17166 18804 17172 18806
rect 17236 18804 17242 18868
rect 5993 18730 6059 18733
rect 14406 18730 14412 18732
rect 5993 18728 14412 18730
rect 5993 18672 5998 18728
rect 6054 18672 14412 18728
rect 5993 18670 14412 18672
rect 5993 18667 6059 18670
rect 14406 18668 14412 18670
rect 14476 18668 14482 18732
rect 15326 18668 15332 18732
rect 15396 18730 15402 18732
rect 16205 18730 16271 18733
rect 16430 18730 16436 18732
rect 15396 18728 16436 18730
rect 15396 18672 16210 18728
rect 16266 18672 16436 18728
rect 15396 18670 16436 18672
rect 15396 18668 15402 18670
rect 16205 18667 16271 18670
rect 16430 18668 16436 18670
rect 16500 18668 16506 18732
rect 0 18594 160 18624
rect 1669 18594 1735 18597
rect 0 18592 1735 18594
rect 0 18536 1674 18592
rect 1730 18536 1735 18592
rect 0 18534 1735 18536
rect 0 18504 160 18534
rect 1669 18531 1735 18534
rect 1853 18594 1919 18597
rect 5441 18594 5507 18597
rect 6085 18594 6151 18597
rect 1853 18592 6151 18594
rect 1853 18536 1858 18592
rect 1914 18536 5446 18592
rect 5502 18536 6090 18592
rect 6146 18536 6151 18592
rect 1853 18534 6151 18536
rect 1853 18531 1919 18534
rect 5441 18531 5507 18534
rect 6085 18531 6151 18534
rect 25129 18594 25195 18597
rect 25840 18594 26000 18624
rect 25129 18592 26000 18594
rect 25129 18536 25134 18592
rect 25190 18536 26000 18592
rect 25129 18534 26000 18536
rect 25129 18531 25195 18534
rect 6880 18528 7196 18529
rect 6880 18464 6886 18528
rect 6950 18464 6966 18528
rect 7030 18464 7046 18528
rect 7110 18464 7126 18528
rect 7190 18464 7196 18528
rect 6880 18463 7196 18464
rect 12814 18528 13130 18529
rect 12814 18464 12820 18528
rect 12884 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13130 18528
rect 12814 18463 13130 18464
rect 18748 18528 19064 18529
rect 18748 18464 18754 18528
rect 18818 18464 18834 18528
rect 18898 18464 18914 18528
rect 18978 18464 18994 18528
rect 19058 18464 19064 18528
rect 18748 18463 19064 18464
rect 24682 18528 24998 18529
rect 24682 18464 24688 18528
rect 24752 18464 24768 18528
rect 24832 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 24998 18528
rect 25840 18504 26000 18534
rect 24682 18463 24998 18464
rect 4153 18458 4219 18461
rect 5625 18458 5691 18461
rect 4153 18456 5691 18458
rect 4153 18400 4158 18456
rect 4214 18400 5630 18456
rect 5686 18400 5691 18456
rect 4153 18398 5691 18400
rect 4153 18395 4219 18398
rect 5625 18395 5691 18398
rect 7925 18458 7991 18461
rect 12617 18458 12683 18461
rect 7925 18456 12683 18458
rect 7925 18400 7930 18456
rect 7986 18400 12622 18456
rect 12678 18400 12683 18456
rect 7925 18398 12683 18400
rect 7925 18395 7991 18398
rect 0 18322 160 18352
rect 1301 18322 1367 18325
rect 0 18320 1367 18322
rect 0 18264 1306 18320
rect 1362 18264 1367 18320
rect 0 18262 1367 18264
rect 0 18232 160 18262
rect 1301 18259 1367 18262
rect 1710 18260 1716 18324
rect 1780 18322 1786 18324
rect 4153 18322 4219 18325
rect 1780 18320 4219 18322
rect 1780 18264 4158 18320
rect 4214 18264 4219 18320
rect 1780 18262 4219 18264
rect 1780 18260 1786 18262
rect 4153 18259 4219 18262
rect 1485 18186 1551 18189
rect 6913 18186 6979 18189
rect 1485 18184 6979 18186
rect 1485 18128 1490 18184
rect 1546 18128 6918 18184
rect 6974 18128 6979 18184
rect 1485 18126 6979 18128
rect 1485 18123 1551 18126
rect 6913 18123 6979 18126
rect 0 18050 160 18080
rect 1209 18050 1275 18053
rect 0 18048 1275 18050
rect 0 17992 1214 18048
rect 1270 17992 1275 18048
rect 0 17990 1275 17992
rect 0 17960 160 17990
rect 1209 17987 1275 17990
rect 4470 17988 4476 18052
rect 4540 18050 4546 18052
rect 7833 18050 7899 18053
rect 4540 18048 7899 18050
rect 4540 17992 7838 18048
rect 7894 17992 7899 18048
rect 4540 17990 7899 17992
rect 4540 17988 4546 17990
rect 7833 17987 7899 17990
rect 10409 18050 10475 18053
rect 10910 18050 10916 18052
rect 10409 18048 10916 18050
rect 10409 17992 10414 18048
rect 10470 17992 10916 18048
rect 10409 17990 10916 17992
rect 10409 17987 10475 17990
rect 10910 17988 10916 17990
rect 10980 17988 10986 18052
rect 12390 18050 12450 18398
rect 12617 18395 12683 18398
rect 12525 18050 12591 18053
rect 12390 18048 12591 18050
rect 12390 17992 12530 18048
rect 12586 17992 12591 18048
rect 12390 17990 12591 17992
rect 12525 17987 12591 17990
rect 13169 18050 13235 18053
rect 15009 18050 15075 18053
rect 15561 18052 15627 18053
rect 15510 18050 15516 18052
rect 13169 18048 15075 18050
rect 13169 17992 13174 18048
rect 13230 17992 15014 18048
rect 15070 17992 15075 18048
rect 13169 17990 15075 17992
rect 15470 17990 15516 18050
rect 15580 18048 15627 18052
rect 15622 17992 15627 18048
rect 13169 17987 13235 17990
rect 15009 17987 15075 17990
rect 15510 17988 15516 17990
rect 15580 17988 15627 17992
rect 15561 17987 15627 17988
rect 24393 18050 24459 18053
rect 25840 18050 26000 18080
rect 24393 18048 26000 18050
rect 24393 17992 24398 18048
rect 24454 17992 26000 18048
rect 24393 17990 26000 17992
rect 24393 17987 24459 17990
rect 3913 17984 4229 17985
rect 3913 17920 3919 17984
rect 3983 17920 3999 17984
rect 4063 17920 4079 17984
rect 4143 17920 4159 17984
rect 4223 17920 4229 17984
rect 3913 17919 4229 17920
rect 9847 17984 10163 17985
rect 9847 17920 9853 17984
rect 9917 17920 9933 17984
rect 9997 17920 10013 17984
rect 10077 17920 10093 17984
rect 10157 17920 10163 17984
rect 9847 17919 10163 17920
rect 15781 17984 16097 17985
rect 15781 17920 15787 17984
rect 15851 17920 15867 17984
rect 15931 17920 15947 17984
rect 16011 17920 16027 17984
rect 16091 17920 16097 17984
rect 15781 17919 16097 17920
rect 21715 17984 22031 17985
rect 21715 17920 21721 17984
rect 21785 17920 21801 17984
rect 21865 17920 21881 17984
rect 21945 17920 21961 17984
rect 22025 17920 22031 17984
rect 25840 17960 26000 17990
rect 21715 17919 22031 17920
rect 1577 17914 1643 17917
rect 16297 17916 16363 17917
rect 798 17912 1643 17914
rect 798 17856 1582 17912
rect 1638 17856 1643 17912
rect 798 17854 1643 17856
rect 0 17778 160 17808
rect 798 17778 858 17854
rect 1577 17851 1643 17854
rect 16246 17852 16252 17916
rect 16316 17914 16363 17916
rect 16316 17912 16408 17914
rect 16358 17856 16408 17912
rect 16316 17854 16408 17856
rect 16316 17852 16363 17854
rect 16297 17851 16363 17852
rect 0 17718 858 17778
rect 3601 17778 3667 17781
rect 5073 17778 5139 17781
rect 3601 17776 5139 17778
rect 3601 17720 3606 17776
rect 3662 17720 5078 17776
rect 5134 17720 5139 17776
rect 3601 17718 5139 17720
rect 0 17688 160 17718
rect 3601 17715 3667 17718
rect 5073 17715 5139 17718
rect 11513 17778 11579 17781
rect 21633 17778 21699 17781
rect 11513 17776 21699 17778
rect 11513 17720 11518 17776
rect 11574 17720 21638 17776
rect 21694 17720 21699 17776
rect 11513 17718 21699 17720
rect 11513 17715 11579 17718
rect 21633 17715 21699 17718
rect 289 17642 355 17645
rect 7281 17642 7347 17645
rect 289 17640 7347 17642
rect 289 17584 294 17640
rect 350 17584 7286 17640
rect 7342 17584 7347 17640
rect 289 17582 7347 17584
rect 289 17579 355 17582
rect 7281 17579 7347 17582
rect 12249 17642 12315 17645
rect 12566 17642 12572 17644
rect 12249 17640 12572 17642
rect 12249 17584 12254 17640
rect 12310 17584 12572 17640
rect 12249 17582 12572 17584
rect 12249 17579 12315 17582
rect 12566 17580 12572 17582
rect 12636 17580 12642 17644
rect 0 17506 160 17536
rect 1761 17506 1827 17509
rect 0 17504 1827 17506
rect 0 17448 1766 17504
rect 1822 17448 1827 17504
rect 0 17446 1827 17448
rect 0 17416 160 17446
rect 1761 17443 1827 17446
rect 25129 17506 25195 17509
rect 25840 17506 26000 17536
rect 25129 17504 26000 17506
rect 25129 17448 25134 17504
rect 25190 17448 26000 17504
rect 25129 17446 26000 17448
rect 25129 17443 25195 17446
rect 6880 17440 7196 17441
rect 6880 17376 6886 17440
rect 6950 17376 6966 17440
rect 7030 17376 7046 17440
rect 7110 17376 7126 17440
rect 7190 17376 7196 17440
rect 6880 17375 7196 17376
rect 12814 17440 13130 17441
rect 12814 17376 12820 17440
rect 12884 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13130 17440
rect 12814 17375 13130 17376
rect 18748 17440 19064 17441
rect 18748 17376 18754 17440
rect 18818 17376 18834 17440
rect 18898 17376 18914 17440
rect 18978 17376 18994 17440
rect 19058 17376 19064 17440
rect 18748 17375 19064 17376
rect 24682 17440 24998 17441
rect 24682 17376 24688 17440
rect 24752 17376 24768 17440
rect 24832 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 24998 17440
rect 25840 17416 26000 17446
rect 24682 17375 24998 17376
rect 1025 17370 1091 17373
rect 5901 17370 5967 17373
rect 1025 17368 5967 17370
rect 1025 17312 1030 17368
rect 1086 17312 5906 17368
rect 5962 17312 5967 17368
rect 1025 17310 5967 17312
rect 1025 17307 1091 17310
rect 5901 17307 5967 17310
rect 9581 17370 9647 17373
rect 9581 17368 11300 17370
rect 9581 17312 9586 17368
rect 9642 17312 11300 17368
rect 9581 17310 11300 17312
rect 9581 17307 9647 17310
rect 0 17234 160 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 160 17174
rect 1485 17171 1551 17174
rect 6637 17234 6703 17237
rect 11053 17234 11119 17237
rect 6637 17232 11119 17234
rect 6637 17176 6642 17232
rect 6698 17176 11058 17232
rect 11114 17176 11119 17232
rect 6637 17174 11119 17176
rect 11240 17234 11300 17310
rect 14089 17234 14155 17237
rect 11240 17232 14155 17234
rect 11240 17176 14094 17232
rect 14150 17176 14155 17232
rect 11240 17174 14155 17176
rect 6637 17171 6703 17174
rect 11053 17171 11119 17174
rect 14089 17171 14155 17174
rect 14549 17234 14615 17237
rect 16614 17234 16620 17236
rect 14549 17232 16620 17234
rect 14549 17176 14554 17232
rect 14610 17176 16620 17232
rect 14549 17174 16620 17176
rect 14549 17171 14615 17174
rect 16614 17172 16620 17174
rect 16684 17172 16690 17236
rect 16982 17172 16988 17236
rect 17052 17234 17058 17236
rect 18229 17234 18295 17237
rect 17052 17232 18295 17234
rect 17052 17176 18234 17232
rect 18290 17176 18295 17232
rect 17052 17174 18295 17176
rect 17052 17172 17058 17174
rect 18229 17171 18295 17174
rect 19149 17234 19215 17237
rect 20110 17234 20116 17236
rect 19149 17232 20116 17234
rect 19149 17176 19154 17232
rect 19210 17176 20116 17232
rect 19149 17174 20116 17176
rect 19149 17171 19215 17174
rect 20110 17172 20116 17174
rect 20180 17172 20186 17236
rect 6821 17098 6887 17101
rect 9121 17098 9187 17101
rect 20294 17098 20300 17100
rect 6821 17096 20300 17098
rect 6821 17040 6826 17096
rect 6882 17040 9126 17096
rect 9182 17040 20300 17096
rect 6821 17038 20300 17040
rect 6821 17035 6887 17038
rect 9121 17035 9187 17038
rect 20294 17036 20300 17038
rect 20364 17036 20370 17100
rect 0 16962 160 16992
rect 2037 16964 2103 16965
rect 2037 16962 2084 16964
rect 0 16902 1042 16962
rect 1992 16960 2084 16962
rect 2148 16962 2154 16964
rect 2313 16962 2379 16965
rect 2148 16960 2379 16962
rect 1992 16904 2042 16960
rect 2148 16904 2318 16960
rect 2374 16904 2379 16960
rect 1992 16902 2084 16904
rect 0 16872 160 16902
rect 982 16826 1042 16902
rect 2037 16900 2084 16902
rect 2148 16902 2379 16904
rect 2148 16900 2154 16902
rect 2037 16899 2103 16900
rect 2313 16899 2379 16902
rect 5625 16962 5691 16965
rect 7189 16962 7255 16965
rect 5625 16960 7255 16962
rect 5625 16904 5630 16960
rect 5686 16904 7194 16960
rect 7250 16904 7255 16960
rect 5625 16902 7255 16904
rect 5625 16899 5691 16902
rect 7189 16899 7255 16902
rect 8150 16900 8156 16964
rect 8220 16962 8226 16964
rect 9438 16962 9444 16964
rect 8220 16902 9444 16962
rect 8220 16900 8226 16902
rect 9438 16900 9444 16902
rect 9508 16900 9514 16964
rect 24117 16962 24183 16965
rect 25840 16962 26000 16992
rect 24117 16960 26000 16962
rect 24117 16904 24122 16960
rect 24178 16904 26000 16960
rect 24117 16902 26000 16904
rect 24117 16899 24183 16902
rect 3913 16896 4229 16897
rect 3913 16832 3919 16896
rect 3983 16832 3999 16896
rect 4063 16832 4079 16896
rect 4143 16832 4159 16896
rect 4223 16832 4229 16896
rect 3913 16831 4229 16832
rect 9847 16896 10163 16897
rect 9847 16832 9853 16896
rect 9917 16832 9933 16896
rect 9997 16832 10013 16896
rect 10077 16832 10093 16896
rect 10157 16832 10163 16896
rect 9847 16831 10163 16832
rect 15781 16896 16097 16897
rect 15781 16832 15787 16896
rect 15851 16832 15867 16896
rect 15931 16832 15947 16896
rect 16011 16832 16027 16896
rect 16091 16832 16097 16896
rect 15781 16831 16097 16832
rect 21715 16896 22031 16897
rect 21715 16832 21721 16896
rect 21785 16832 21801 16896
rect 21865 16832 21881 16896
rect 21945 16832 21961 16896
rect 22025 16832 22031 16896
rect 25840 16872 26000 16902
rect 21715 16831 22031 16832
rect 2037 16826 2103 16829
rect 982 16824 2103 16826
rect 982 16768 2042 16824
rect 2098 16768 2103 16824
rect 982 16766 2103 16768
rect 2037 16763 2103 16766
rect 0 16690 160 16720
rect 2865 16690 2931 16693
rect 0 16688 2931 16690
rect 0 16632 2870 16688
rect 2926 16632 2931 16688
rect 0 16630 2931 16632
rect 0 16600 160 16630
rect 2865 16627 2931 16630
rect 6821 16690 6887 16693
rect 8661 16690 8727 16693
rect 6821 16688 8727 16690
rect 6821 16632 6826 16688
rect 6882 16632 8666 16688
rect 8722 16632 8727 16688
rect 6821 16630 8727 16632
rect 6821 16627 6887 16630
rect 8661 16627 8727 16630
rect 12525 16692 12591 16693
rect 12525 16688 12572 16692
rect 12636 16690 12642 16692
rect 14089 16690 14155 16693
rect 12525 16632 12530 16688
rect 12525 16628 12572 16632
rect 12636 16630 12682 16690
rect 14046 16688 14155 16690
rect 14046 16632 14094 16688
rect 14150 16632 14155 16688
rect 12636 16628 12642 16630
rect 12525 16627 12591 16628
rect 14046 16627 14155 16632
rect 15009 16690 15075 16693
rect 15142 16690 15148 16692
rect 15009 16688 15148 16690
rect 15009 16632 15014 16688
rect 15070 16632 15148 16688
rect 15009 16630 15148 16632
rect 15009 16627 15075 16630
rect 15142 16628 15148 16630
rect 15212 16628 15218 16692
rect 20662 16628 20668 16692
rect 20732 16690 20738 16692
rect 20897 16690 20963 16693
rect 20732 16688 20963 16690
rect 20732 16632 20902 16688
rect 20958 16632 20963 16688
rect 20732 16630 20963 16632
rect 20732 16628 20738 16630
rect 20897 16627 20963 16630
rect 2405 16556 2471 16557
rect 2405 16552 2452 16556
rect 2516 16554 2522 16556
rect 2405 16496 2410 16552
rect 2405 16492 2452 16496
rect 2516 16494 2562 16554
rect 2516 16492 2522 16494
rect 5022 16492 5028 16556
rect 5092 16554 5098 16556
rect 8702 16554 8708 16556
rect 5092 16494 8708 16554
rect 5092 16492 5098 16494
rect 8702 16492 8708 16494
rect 8772 16492 8778 16556
rect 8845 16554 8911 16557
rect 14046 16554 14106 16627
rect 16021 16554 16087 16557
rect 8845 16552 16087 16554
rect 8845 16496 8850 16552
rect 8906 16496 16026 16552
rect 16082 16496 16087 16552
rect 8845 16494 16087 16496
rect 2405 16491 2471 16492
rect 8845 16491 8911 16494
rect 16021 16491 16087 16494
rect 19333 16556 19399 16557
rect 19333 16552 19380 16556
rect 19444 16554 19450 16556
rect 19333 16496 19338 16552
rect 19333 16492 19380 16496
rect 19444 16494 19490 16554
rect 19444 16492 19450 16494
rect 19333 16491 19399 16492
rect 0 16418 160 16448
rect 3969 16418 4035 16421
rect 0 16416 4035 16418
rect 0 16360 3974 16416
rect 4030 16360 4035 16416
rect 0 16358 4035 16360
rect 0 16328 160 16358
rect 3969 16355 4035 16358
rect 25221 16418 25287 16421
rect 25840 16418 26000 16448
rect 25221 16416 26000 16418
rect 25221 16360 25226 16416
rect 25282 16360 26000 16416
rect 25221 16358 26000 16360
rect 25221 16355 25287 16358
rect 6880 16352 7196 16353
rect 6880 16288 6886 16352
rect 6950 16288 6966 16352
rect 7030 16288 7046 16352
rect 7110 16288 7126 16352
rect 7190 16288 7196 16352
rect 6880 16287 7196 16288
rect 12814 16352 13130 16353
rect 12814 16288 12820 16352
rect 12884 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13130 16352
rect 12814 16287 13130 16288
rect 18748 16352 19064 16353
rect 18748 16288 18754 16352
rect 18818 16288 18834 16352
rect 18898 16288 18914 16352
rect 18978 16288 18994 16352
rect 19058 16288 19064 16352
rect 18748 16287 19064 16288
rect 24682 16352 24998 16353
rect 24682 16288 24688 16352
rect 24752 16288 24768 16352
rect 24832 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 24998 16352
rect 25840 16328 26000 16358
rect 24682 16287 24998 16288
rect 3325 16282 3391 16285
rect 3550 16282 3556 16284
rect 3325 16280 3556 16282
rect 3325 16224 3330 16280
rect 3386 16224 3556 16280
rect 3325 16222 3556 16224
rect 3325 16219 3391 16222
rect 3550 16220 3556 16222
rect 3620 16220 3626 16284
rect 0 16146 160 16176
rect 3049 16146 3115 16149
rect 0 16144 3115 16146
rect 0 16088 3054 16144
rect 3110 16088 3115 16144
rect 0 16086 3115 16088
rect 0 16056 160 16086
rect 3049 16083 3115 16086
rect 10910 16084 10916 16148
rect 10980 16146 10986 16148
rect 14089 16146 14155 16149
rect 10980 16144 14155 16146
rect 10980 16088 14094 16144
rect 14150 16088 14155 16144
rect 10980 16086 14155 16088
rect 10980 16084 10986 16086
rect 14089 16083 14155 16086
rect 17166 16084 17172 16148
rect 17236 16146 17242 16148
rect 22185 16146 22251 16149
rect 17236 16144 22251 16146
rect 17236 16088 22190 16144
rect 22246 16088 22251 16144
rect 17236 16086 22251 16088
rect 17236 16084 17242 16086
rect 22185 16083 22251 16086
rect 14038 15948 14044 16012
rect 14108 16010 14114 16012
rect 20069 16010 20135 16013
rect 14108 16008 20135 16010
rect 14108 15952 20074 16008
rect 20130 15952 20135 16008
rect 14108 15950 20135 15952
rect 14108 15948 14114 15950
rect 20069 15947 20135 15950
rect 0 15874 160 15904
rect 24117 15874 24183 15877
rect 25840 15874 26000 15904
rect 0 15814 3434 15874
rect 0 15784 160 15814
rect 0 15602 160 15632
rect 3049 15602 3115 15605
rect 0 15600 3115 15602
rect 0 15544 3054 15600
rect 3110 15544 3115 15600
rect 0 15542 3115 15544
rect 3374 15602 3434 15814
rect 24117 15872 26000 15874
rect 24117 15816 24122 15872
rect 24178 15816 26000 15872
rect 24117 15814 26000 15816
rect 24117 15811 24183 15814
rect 3913 15808 4229 15809
rect 3913 15744 3919 15808
rect 3983 15744 3999 15808
rect 4063 15744 4079 15808
rect 4143 15744 4159 15808
rect 4223 15744 4229 15808
rect 3913 15743 4229 15744
rect 9847 15808 10163 15809
rect 9847 15744 9853 15808
rect 9917 15744 9933 15808
rect 9997 15744 10013 15808
rect 10077 15744 10093 15808
rect 10157 15744 10163 15808
rect 9847 15743 10163 15744
rect 15781 15808 16097 15809
rect 15781 15744 15787 15808
rect 15851 15744 15867 15808
rect 15931 15744 15947 15808
rect 16011 15744 16027 15808
rect 16091 15744 16097 15808
rect 15781 15743 16097 15744
rect 21715 15808 22031 15809
rect 21715 15744 21721 15808
rect 21785 15744 21801 15808
rect 21865 15744 21881 15808
rect 21945 15744 21961 15808
rect 22025 15744 22031 15808
rect 25840 15784 26000 15814
rect 21715 15743 22031 15744
rect 3969 15602 4035 15605
rect 3374 15600 4035 15602
rect 3374 15544 3974 15600
rect 4030 15544 4035 15600
rect 3374 15542 4035 15544
rect 0 15512 160 15542
rect 3049 15539 3115 15542
rect 3969 15539 4035 15542
rect 4153 15602 4219 15605
rect 4654 15602 4660 15604
rect 4153 15600 4660 15602
rect 4153 15544 4158 15600
rect 4214 15544 4660 15600
rect 4153 15542 4660 15544
rect 4153 15539 4219 15542
rect 4654 15540 4660 15542
rect 4724 15540 4730 15604
rect 8334 15540 8340 15604
rect 8404 15602 8410 15604
rect 9397 15602 9463 15605
rect 16573 15602 16639 15605
rect 8404 15600 16639 15602
rect 8404 15544 9402 15600
rect 9458 15544 16578 15600
rect 16634 15544 16639 15600
rect 8404 15542 16639 15544
rect 8404 15540 8410 15542
rect 9397 15539 9463 15542
rect 16573 15539 16639 15542
rect 12341 15466 12407 15469
rect 13302 15466 13308 15468
rect 12341 15464 13308 15466
rect 12341 15408 12346 15464
rect 12402 15408 13308 15464
rect 12341 15406 13308 15408
rect 12341 15403 12407 15406
rect 13302 15404 13308 15406
rect 13372 15404 13378 15468
rect 17350 15404 17356 15468
rect 17420 15466 17426 15468
rect 22686 15466 22692 15468
rect 17420 15406 22692 15466
rect 17420 15404 17426 15406
rect 22686 15404 22692 15406
rect 22756 15404 22762 15468
rect 0 15330 160 15360
rect 1393 15330 1459 15333
rect 0 15328 1459 15330
rect 0 15272 1398 15328
rect 1454 15272 1459 15328
rect 0 15270 1459 15272
rect 0 15240 160 15270
rect 1393 15267 1459 15270
rect 25313 15330 25379 15333
rect 25840 15330 26000 15360
rect 25313 15328 26000 15330
rect 25313 15272 25318 15328
rect 25374 15272 26000 15328
rect 25313 15270 26000 15272
rect 25313 15267 25379 15270
rect 6880 15264 7196 15265
rect 6880 15200 6886 15264
rect 6950 15200 6966 15264
rect 7030 15200 7046 15264
rect 7110 15200 7126 15264
rect 7190 15200 7196 15264
rect 6880 15199 7196 15200
rect 12814 15264 13130 15265
rect 12814 15200 12820 15264
rect 12884 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13130 15264
rect 12814 15199 13130 15200
rect 18748 15264 19064 15265
rect 18748 15200 18754 15264
rect 18818 15200 18834 15264
rect 18898 15200 18914 15264
rect 18978 15200 18994 15264
rect 19058 15200 19064 15264
rect 18748 15199 19064 15200
rect 24682 15264 24998 15265
rect 24682 15200 24688 15264
rect 24752 15200 24768 15264
rect 24832 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 24998 15264
rect 25840 15240 26000 15270
rect 24682 15199 24998 15200
rect 5073 15194 5139 15197
rect 5206 15194 5212 15196
rect 5073 15192 5212 15194
rect 5073 15136 5078 15192
rect 5134 15136 5212 15192
rect 5073 15134 5212 15136
rect 5073 15131 5139 15134
rect 5206 15132 5212 15134
rect 5276 15132 5282 15196
rect 9949 15194 10015 15197
rect 10358 15194 10364 15196
rect 9949 15192 10364 15194
rect 9949 15136 9954 15192
rect 10010 15136 10364 15192
rect 9949 15134 10364 15136
rect 9949 15131 10015 15134
rect 10358 15132 10364 15134
rect 10428 15194 10434 15196
rect 12065 15194 12131 15197
rect 10428 15192 12131 15194
rect 10428 15136 12070 15192
rect 12126 15136 12131 15192
rect 10428 15134 12131 15136
rect 10428 15132 10434 15134
rect 12065 15131 12131 15134
rect 0 15058 160 15088
rect 2313 15058 2379 15061
rect 0 15056 2379 15058
rect 0 15000 2318 15056
rect 2374 15000 2379 15056
rect 0 14998 2379 15000
rect 0 14968 160 14998
rect 2313 14995 2379 14998
rect 6494 14996 6500 15060
rect 6564 15058 6570 15060
rect 6637 15058 6703 15061
rect 6564 15056 6703 15058
rect 6564 15000 6642 15056
rect 6698 15000 6703 15056
rect 6564 14998 6703 15000
rect 6564 14996 6570 14998
rect 6637 14995 6703 14998
rect 3693 14922 3759 14925
rect 7833 14922 7899 14925
rect 3693 14920 7899 14922
rect 3693 14864 3698 14920
rect 3754 14864 7838 14920
rect 7894 14864 7899 14920
rect 3693 14862 7899 14864
rect 3693 14859 3759 14862
rect 7833 14859 7899 14862
rect 10685 14922 10751 14925
rect 17125 14922 17191 14925
rect 10685 14920 17191 14922
rect 10685 14864 10690 14920
rect 10746 14864 17130 14920
rect 17186 14864 17191 14920
rect 10685 14862 17191 14864
rect 10685 14859 10751 14862
rect 17125 14859 17191 14862
rect 0 14786 160 14816
rect 2773 14786 2839 14789
rect 0 14784 2839 14786
rect 0 14728 2778 14784
rect 2834 14728 2839 14784
rect 0 14726 2839 14728
rect 0 14696 160 14726
rect 2773 14723 2839 14726
rect 24025 14786 24091 14789
rect 25840 14786 26000 14816
rect 24025 14784 26000 14786
rect 24025 14728 24030 14784
rect 24086 14728 26000 14784
rect 24025 14726 26000 14728
rect 24025 14723 24091 14726
rect 3913 14720 4229 14721
rect 3913 14656 3919 14720
rect 3983 14656 3999 14720
rect 4063 14656 4079 14720
rect 4143 14656 4159 14720
rect 4223 14656 4229 14720
rect 3913 14655 4229 14656
rect 9847 14720 10163 14721
rect 9847 14656 9853 14720
rect 9917 14656 9933 14720
rect 9997 14656 10013 14720
rect 10077 14656 10093 14720
rect 10157 14656 10163 14720
rect 9847 14655 10163 14656
rect 15781 14720 16097 14721
rect 15781 14656 15787 14720
rect 15851 14656 15867 14720
rect 15931 14656 15947 14720
rect 16011 14656 16027 14720
rect 16091 14656 16097 14720
rect 15781 14655 16097 14656
rect 21715 14720 22031 14721
rect 21715 14656 21721 14720
rect 21785 14656 21801 14720
rect 21865 14656 21881 14720
rect 21945 14656 21961 14720
rect 22025 14656 22031 14720
rect 25840 14696 26000 14726
rect 21715 14655 22031 14656
rect 16205 14650 16271 14653
rect 16205 14648 17280 14650
rect 16205 14592 16210 14648
rect 16266 14592 17280 14648
rect 16205 14590 17280 14592
rect 16205 14587 16271 14590
rect 0 14514 160 14544
rect 17220 14517 17280 14590
rect 3325 14514 3391 14517
rect 0 14512 3391 14514
rect 0 14456 3330 14512
rect 3386 14456 3391 14512
rect 0 14454 3391 14456
rect 0 14424 160 14454
rect 3325 14451 3391 14454
rect 4245 14514 4311 14517
rect 15285 14514 15351 14517
rect 4245 14512 15351 14514
rect 4245 14456 4250 14512
rect 4306 14456 15290 14512
rect 15346 14456 15351 14512
rect 4245 14454 15351 14456
rect 4245 14451 4311 14454
rect 15285 14451 15351 14454
rect 16021 14514 16087 14517
rect 16297 14514 16363 14517
rect 16021 14512 16363 14514
rect 16021 14456 16026 14512
rect 16082 14456 16302 14512
rect 16358 14456 16363 14512
rect 16021 14454 16363 14456
rect 16021 14451 16087 14454
rect 16297 14451 16363 14454
rect 16757 14512 16823 14517
rect 16757 14456 16762 14512
rect 16818 14456 16823 14512
rect 16757 14451 16823 14456
rect 17217 14512 17283 14517
rect 17217 14456 17222 14512
rect 17278 14456 17283 14512
rect 17217 14451 17283 14456
rect 1853 14378 1919 14381
rect 4797 14378 4863 14381
rect 1853 14376 4863 14378
rect 1853 14320 1858 14376
rect 1914 14320 4802 14376
rect 4858 14320 4863 14376
rect 1853 14318 4863 14320
rect 1853 14315 1919 14318
rect 4797 14315 4863 14318
rect 6453 14378 6519 14381
rect 6913 14378 6979 14381
rect 6453 14376 6979 14378
rect 6453 14320 6458 14376
rect 6514 14320 6918 14376
rect 6974 14320 6979 14376
rect 6453 14318 6979 14320
rect 6453 14315 6519 14318
rect 6913 14315 6979 14318
rect 0 14242 160 14272
rect 16760 14245 16820 14451
rect 10041 14242 10107 14245
rect 10409 14242 10475 14245
rect 0 14182 1962 14242
rect 0 14152 160 14182
rect 0 13970 160 14000
rect 1669 13970 1735 13973
rect 0 13968 1735 13970
rect 0 13912 1674 13968
rect 1730 13912 1735 13968
rect 0 13910 1735 13912
rect 0 13880 160 13910
rect 1669 13907 1735 13910
rect 1761 13834 1827 13837
rect 1902 13834 1962 14182
rect 10041 14240 10475 14242
rect 10041 14184 10046 14240
rect 10102 14184 10414 14240
rect 10470 14184 10475 14240
rect 10041 14182 10475 14184
rect 10041 14179 10107 14182
rect 10409 14179 10475 14182
rect 16757 14240 16823 14245
rect 16757 14184 16762 14240
rect 16818 14184 16823 14240
rect 16757 14179 16823 14184
rect 25129 14242 25195 14245
rect 25840 14242 26000 14272
rect 25129 14240 26000 14242
rect 25129 14184 25134 14240
rect 25190 14184 26000 14240
rect 25129 14182 26000 14184
rect 25129 14179 25195 14182
rect 6880 14176 7196 14177
rect 6880 14112 6886 14176
rect 6950 14112 6966 14176
rect 7030 14112 7046 14176
rect 7110 14112 7126 14176
rect 7190 14112 7196 14176
rect 6880 14111 7196 14112
rect 12814 14176 13130 14177
rect 12814 14112 12820 14176
rect 12884 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13130 14176
rect 12814 14111 13130 14112
rect 18748 14176 19064 14177
rect 18748 14112 18754 14176
rect 18818 14112 18834 14176
rect 18898 14112 18914 14176
rect 18978 14112 18994 14176
rect 19058 14112 19064 14176
rect 18748 14111 19064 14112
rect 24682 14176 24998 14177
rect 24682 14112 24688 14176
rect 24752 14112 24768 14176
rect 24832 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 24998 14176
rect 25840 14152 26000 14182
rect 24682 14111 24998 14112
rect 4337 13970 4403 13973
rect 7373 13970 7439 13973
rect 4337 13968 7439 13970
rect 4337 13912 4342 13968
rect 4398 13912 7378 13968
rect 7434 13912 7439 13968
rect 4337 13910 7439 13912
rect 4337 13907 4403 13910
rect 7373 13907 7439 13910
rect 11145 13970 11211 13973
rect 14273 13970 14339 13973
rect 11145 13968 14339 13970
rect 11145 13912 11150 13968
rect 11206 13912 14278 13968
rect 14334 13912 14339 13968
rect 11145 13910 14339 13912
rect 11145 13907 11211 13910
rect 14273 13907 14339 13910
rect 22093 13970 22159 13973
rect 22921 13970 22987 13973
rect 22093 13968 22987 13970
rect 22093 13912 22098 13968
rect 22154 13912 22926 13968
rect 22982 13912 22987 13968
rect 22093 13910 22987 13912
rect 22093 13907 22159 13910
rect 22921 13907 22987 13910
rect 1761 13832 1962 13834
rect 1761 13776 1766 13832
rect 1822 13776 1962 13832
rect 1761 13774 1962 13776
rect 1761 13771 1827 13774
rect 4838 13772 4844 13836
rect 4908 13834 4914 13836
rect 5073 13834 5139 13837
rect 4908 13832 5139 13834
rect 4908 13776 5078 13832
rect 5134 13776 5139 13832
rect 4908 13774 5139 13776
rect 4908 13772 4914 13774
rect 5073 13771 5139 13774
rect 13169 13834 13235 13837
rect 13445 13834 13511 13837
rect 13169 13832 13554 13834
rect 13169 13776 13174 13832
rect 13230 13776 13450 13832
rect 13506 13776 13554 13832
rect 13169 13774 13554 13776
rect 13169 13771 13235 13774
rect 13445 13771 13554 13774
rect 0 13698 160 13728
rect 1301 13698 1367 13701
rect 0 13696 1367 13698
rect 0 13640 1306 13696
rect 1362 13640 1367 13696
rect 0 13638 1367 13640
rect 0 13608 160 13638
rect 1301 13635 1367 13638
rect 1485 13698 1551 13701
rect 2262 13698 2268 13700
rect 1485 13696 2268 13698
rect 1485 13640 1490 13696
rect 1546 13640 2268 13696
rect 1485 13638 2268 13640
rect 1485 13635 1551 13638
rect 2262 13636 2268 13638
rect 2332 13636 2338 13700
rect 8477 13698 8543 13701
rect 9622 13698 9628 13700
rect 8477 13696 9628 13698
rect 8477 13640 8482 13696
rect 8538 13640 9628 13696
rect 8477 13638 9628 13640
rect 8477 13635 8543 13638
rect 9622 13636 9628 13638
rect 9692 13636 9698 13700
rect 3913 13632 4229 13633
rect 3913 13568 3919 13632
rect 3983 13568 3999 13632
rect 4063 13568 4079 13632
rect 4143 13568 4159 13632
rect 4223 13568 4229 13632
rect 3913 13567 4229 13568
rect 9847 13632 10163 13633
rect 9847 13568 9853 13632
rect 9917 13568 9933 13632
rect 9997 13568 10013 13632
rect 10077 13568 10093 13632
rect 10157 13568 10163 13632
rect 9847 13567 10163 13568
rect 13494 13565 13554 13771
rect 19926 13636 19932 13700
rect 19996 13698 20002 13700
rect 20897 13698 20963 13701
rect 19996 13696 20963 13698
rect 19996 13640 20902 13696
rect 20958 13640 20963 13696
rect 19996 13638 20963 13640
rect 19996 13636 20002 13638
rect 20897 13635 20963 13638
rect 22093 13698 22159 13701
rect 23289 13698 23355 13701
rect 22093 13696 23355 13698
rect 22093 13640 22098 13696
rect 22154 13640 23294 13696
rect 23350 13640 23355 13696
rect 22093 13638 23355 13640
rect 22093 13635 22159 13638
rect 23289 13635 23355 13638
rect 24393 13698 24459 13701
rect 25840 13698 26000 13728
rect 24393 13696 26000 13698
rect 24393 13640 24398 13696
rect 24454 13640 26000 13696
rect 24393 13638 26000 13640
rect 24393 13635 24459 13638
rect 15781 13632 16097 13633
rect 15781 13568 15787 13632
rect 15851 13568 15867 13632
rect 15931 13568 15947 13632
rect 16011 13568 16027 13632
rect 16091 13568 16097 13632
rect 15781 13567 16097 13568
rect 21715 13632 22031 13633
rect 21715 13568 21721 13632
rect 21785 13568 21801 13632
rect 21865 13568 21881 13632
rect 21945 13568 21961 13632
rect 22025 13568 22031 13632
rect 25840 13608 26000 13638
rect 21715 13567 22031 13568
rect 13494 13560 13603 13565
rect 13494 13504 13542 13560
rect 13598 13504 13603 13560
rect 13494 13502 13603 13504
rect 13537 13499 13603 13502
rect 19793 13562 19859 13565
rect 20846 13562 20852 13564
rect 19793 13560 20852 13562
rect 19793 13504 19798 13560
rect 19854 13504 20852 13560
rect 19793 13502 20852 13504
rect 19793 13499 19859 13502
rect 20846 13500 20852 13502
rect 20916 13500 20922 13564
rect 22553 13562 22619 13565
rect 23197 13562 23263 13565
rect 22553 13560 23263 13562
rect 22553 13504 22558 13560
rect 22614 13504 23202 13560
rect 23258 13504 23263 13560
rect 22553 13502 23263 13504
rect 22553 13499 22619 13502
rect 23197 13499 23263 13502
rect 0 13426 160 13456
rect 4061 13426 4127 13429
rect 0 13424 4127 13426
rect 0 13368 4066 13424
rect 4122 13368 4127 13424
rect 0 13366 4127 13368
rect 0 13336 160 13366
rect 4061 13363 4127 13366
rect 9254 13364 9260 13428
rect 9324 13426 9330 13428
rect 15193 13426 15259 13429
rect 9324 13424 15259 13426
rect 9324 13368 15198 13424
rect 15254 13368 15259 13424
rect 9324 13366 15259 13368
rect 9324 13364 9330 13366
rect 15193 13363 15259 13366
rect 3550 13228 3556 13292
rect 3620 13290 3626 13292
rect 3877 13290 3943 13293
rect 3620 13288 3943 13290
rect 3620 13232 3882 13288
rect 3938 13232 3943 13288
rect 3620 13230 3943 13232
rect 3620 13228 3626 13230
rect 3877 13227 3943 13230
rect 10409 13290 10475 13293
rect 10685 13290 10751 13293
rect 10409 13288 10751 13290
rect 10409 13232 10414 13288
rect 10470 13232 10690 13288
rect 10746 13232 10751 13288
rect 10409 13230 10751 13232
rect 10409 13227 10475 13230
rect 10685 13227 10751 13230
rect 19977 13290 20043 13293
rect 20529 13290 20595 13293
rect 19977 13288 20595 13290
rect 19977 13232 19982 13288
rect 20038 13232 20534 13288
rect 20590 13232 20595 13288
rect 19977 13230 20595 13232
rect 19977 13227 20043 13230
rect 20529 13227 20595 13230
rect 0 13154 160 13184
rect 1209 13154 1275 13157
rect 0 13152 1275 13154
rect 0 13096 1214 13152
rect 1270 13096 1275 13152
rect 0 13094 1275 13096
rect 0 13064 160 13094
rect 1209 13091 1275 13094
rect 10133 13154 10199 13157
rect 11605 13154 11671 13157
rect 25840 13154 26000 13184
rect 10133 13152 11671 13154
rect 10133 13096 10138 13152
rect 10194 13096 11610 13152
rect 11666 13096 11671 13152
rect 10133 13094 11671 13096
rect 10133 13091 10199 13094
rect 11605 13091 11671 13094
rect 25454 13094 26000 13154
rect 6880 13088 7196 13089
rect 6880 13024 6886 13088
rect 6950 13024 6966 13088
rect 7030 13024 7046 13088
rect 7110 13024 7126 13088
rect 7190 13024 7196 13088
rect 6880 13023 7196 13024
rect 12814 13088 13130 13089
rect 12814 13024 12820 13088
rect 12884 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13130 13088
rect 12814 13023 13130 13024
rect 18748 13088 19064 13089
rect 18748 13024 18754 13088
rect 18818 13024 18834 13088
rect 18898 13024 18914 13088
rect 18978 13024 18994 13088
rect 19058 13024 19064 13088
rect 18748 13023 19064 13024
rect 24682 13088 24998 13089
rect 24682 13024 24688 13088
rect 24752 13024 24768 13088
rect 24832 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 24998 13088
rect 24682 13023 24998 13024
rect 1853 13018 1919 13021
rect 1853 13016 2790 13018
rect 1853 12960 1858 13016
rect 1914 12960 2790 13016
rect 1853 12958 2790 12960
rect 1853 12955 1919 12958
rect 0 12882 160 12912
rect 2129 12882 2195 12885
rect 0 12880 2195 12882
rect 0 12824 2134 12880
rect 2190 12824 2195 12880
rect 0 12822 2195 12824
rect 0 12792 160 12822
rect 2129 12819 2195 12822
rect 2730 12746 2790 12958
rect 3693 12882 3759 12885
rect 8385 12882 8451 12885
rect 3693 12880 8451 12882
rect 3693 12824 3698 12880
rect 3754 12824 8390 12880
rect 8446 12824 8451 12880
rect 3693 12822 8451 12824
rect 3693 12819 3759 12822
rect 8385 12819 8451 12822
rect 7925 12746 7991 12749
rect 2730 12744 7991 12746
rect 2730 12688 7930 12744
rect 7986 12688 7991 12744
rect 2730 12686 7991 12688
rect 7925 12683 7991 12686
rect 25129 12746 25195 12749
rect 25454 12746 25514 13094
rect 25840 13064 26000 13094
rect 25129 12744 25514 12746
rect 25129 12688 25134 12744
rect 25190 12688 25514 12744
rect 25129 12686 25514 12688
rect 25129 12683 25195 12686
rect 0 12610 160 12640
rect 1577 12610 1643 12613
rect 0 12608 1643 12610
rect 0 12552 1582 12608
rect 1638 12552 1643 12608
rect 0 12550 1643 12552
rect 0 12520 160 12550
rect 1577 12547 1643 12550
rect 4797 12610 4863 12613
rect 5441 12610 5507 12613
rect 7373 12610 7439 12613
rect 4797 12608 7439 12610
rect 4797 12552 4802 12608
rect 4858 12552 5446 12608
rect 5502 12552 7378 12608
rect 7434 12552 7439 12608
rect 4797 12550 7439 12552
rect 4797 12547 4863 12550
rect 5441 12547 5507 12550
rect 7373 12547 7439 12550
rect 24209 12610 24275 12613
rect 25840 12610 26000 12640
rect 24209 12608 26000 12610
rect 24209 12552 24214 12608
rect 24270 12552 26000 12608
rect 24209 12550 26000 12552
rect 24209 12547 24275 12550
rect 3913 12544 4229 12545
rect 3913 12480 3919 12544
rect 3983 12480 3999 12544
rect 4063 12480 4079 12544
rect 4143 12480 4159 12544
rect 4223 12480 4229 12544
rect 3913 12479 4229 12480
rect 9847 12544 10163 12545
rect 9847 12480 9853 12544
rect 9917 12480 9933 12544
rect 9997 12480 10013 12544
rect 10077 12480 10093 12544
rect 10157 12480 10163 12544
rect 9847 12479 10163 12480
rect 15781 12544 16097 12545
rect 15781 12480 15787 12544
rect 15851 12480 15867 12544
rect 15931 12480 15947 12544
rect 16011 12480 16027 12544
rect 16091 12480 16097 12544
rect 15781 12479 16097 12480
rect 21715 12544 22031 12545
rect 21715 12480 21721 12544
rect 21785 12480 21801 12544
rect 21865 12480 21881 12544
rect 21945 12480 21961 12544
rect 22025 12480 22031 12544
rect 25840 12520 26000 12550
rect 21715 12479 22031 12480
rect 3233 12476 3299 12477
rect 3182 12412 3188 12476
rect 3252 12474 3299 12476
rect 3252 12472 3344 12474
rect 3294 12416 3344 12472
rect 3252 12414 3344 12416
rect 3252 12412 3299 12414
rect 6494 12412 6500 12476
rect 6564 12474 6570 12476
rect 6821 12474 6887 12477
rect 6564 12472 6887 12474
rect 6564 12416 6826 12472
rect 6882 12416 6887 12472
rect 6564 12414 6887 12416
rect 6564 12412 6570 12414
rect 3233 12411 3299 12412
rect 6821 12411 6887 12414
rect 7097 12474 7163 12477
rect 8477 12474 8543 12477
rect 7097 12472 8543 12474
rect 7097 12416 7102 12472
rect 7158 12416 8482 12472
rect 8538 12416 8543 12472
rect 7097 12414 8543 12416
rect 7097 12411 7163 12414
rect 8477 12411 8543 12414
rect 0 12338 160 12368
rect 3785 12338 3851 12341
rect 0 12336 3851 12338
rect 0 12280 3790 12336
rect 3846 12280 3851 12336
rect 0 12278 3851 12280
rect 0 12248 160 12278
rect 3785 12275 3851 12278
rect 4613 12338 4679 12341
rect 4981 12338 5047 12341
rect 4613 12336 5047 12338
rect 4613 12280 4618 12336
rect 4674 12280 4986 12336
rect 5042 12280 5047 12336
rect 4613 12278 5047 12280
rect 4613 12275 4679 12278
rect 4981 12275 5047 12278
rect 5390 12276 5396 12340
rect 5460 12338 5466 12340
rect 5717 12338 5783 12341
rect 5460 12336 5783 12338
rect 5460 12280 5722 12336
rect 5778 12280 5783 12336
rect 5460 12278 5783 12280
rect 5460 12276 5466 12278
rect 5717 12275 5783 12278
rect 6269 12338 6335 12341
rect 8017 12338 8083 12341
rect 6269 12336 8083 12338
rect 6269 12280 6274 12336
rect 6330 12280 8022 12336
rect 8078 12280 8083 12336
rect 6269 12278 8083 12280
rect 6269 12275 6335 12278
rect 8017 12275 8083 12278
rect 10501 12338 10567 12341
rect 10910 12338 10916 12340
rect 10501 12336 10916 12338
rect 10501 12280 10506 12336
rect 10562 12280 10916 12336
rect 10501 12278 10916 12280
rect 10501 12275 10567 12278
rect 10910 12276 10916 12278
rect 10980 12276 10986 12340
rect 11237 12338 11303 12341
rect 19149 12338 19215 12341
rect 11237 12336 19215 12338
rect 11237 12280 11242 12336
rect 11298 12280 19154 12336
rect 19210 12280 19215 12336
rect 11237 12278 19215 12280
rect 11237 12275 11303 12278
rect 19149 12275 19215 12278
rect 2865 12202 2931 12205
rect 4797 12202 4863 12205
rect 2865 12200 4863 12202
rect 2865 12144 2870 12200
rect 2926 12144 4802 12200
rect 4858 12144 4863 12200
rect 2865 12142 4863 12144
rect 2865 12139 2931 12142
rect 4797 12139 4863 12142
rect 6361 12202 6427 12205
rect 7373 12202 7439 12205
rect 8886 12202 8892 12204
rect 6361 12200 8892 12202
rect 6361 12144 6366 12200
rect 6422 12144 7378 12200
rect 7434 12144 8892 12200
rect 6361 12142 8892 12144
rect 6361 12139 6427 12142
rect 7373 12139 7439 12142
rect 8886 12140 8892 12142
rect 8956 12202 8962 12204
rect 18321 12202 18387 12205
rect 8956 12200 18387 12202
rect 8956 12144 18326 12200
rect 18382 12144 18387 12200
rect 8956 12142 18387 12144
rect 8956 12140 8962 12142
rect 18321 12139 18387 12142
rect 0 12066 160 12096
rect 1393 12066 1459 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 160 12006
rect 1393 12003 1459 12006
rect 3693 12066 3759 12069
rect 3969 12066 4035 12069
rect 4654 12066 4660 12068
rect 3693 12064 4660 12066
rect 3693 12008 3698 12064
rect 3754 12008 3974 12064
rect 4030 12008 4660 12064
rect 3693 12006 4660 12008
rect 3693 12003 3759 12006
rect 3969 12003 4035 12006
rect 4654 12004 4660 12006
rect 4724 12004 4730 12068
rect 14917 12066 14983 12069
rect 15837 12066 15903 12069
rect 14917 12064 15903 12066
rect 14917 12008 14922 12064
rect 14978 12008 15842 12064
rect 15898 12008 15903 12064
rect 14917 12006 15903 12008
rect 14917 12003 14983 12006
rect 15837 12003 15903 12006
rect 25221 12066 25287 12069
rect 25840 12066 26000 12096
rect 25221 12064 26000 12066
rect 25221 12008 25226 12064
rect 25282 12008 26000 12064
rect 25221 12006 26000 12008
rect 25221 12003 25287 12006
rect 6880 12000 7196 12001
rect 6880 11936 6886 12000
rect 6950 11936 6966 12000
rect 7030 11936 7046 12000
rect 7110 11936 7126 12000
rect 7190 11936 7196 12000
rect 6880 11935 7196 11936
rect 12814 12000 13130 12001
rect 12814 11936 12820 12000
rect 12884 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13130 12000
rect 12814 11935 13130 11936
rect 18748 12000 19064 12001
rect 18748 11936 18754 12000
rect 18818 11936 18834 12000
rect 18898 11936 18914 12000
rect 18978 11936 18994 12000
rect 19058 11936 19064 12000
rect 18748 11935 19064 11936
rect 24682 12000 24998 12001
rect 24682 11936 24688 12000
rect 24752 11936 24768 12000
rect 24832 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 24998 12000
rect 25840 11976 26000 12006
rect 24682 11935 24998 11936
rect 13721 11930 13787 11933
rect 15326 11930 15332 11932
rect 13721 11928 15332 11930
rect 13721 11872 13726 11928
rect 13782 11872 15332 11928
rect 13721 11870 15332 11872
rect 13721 11867 13787 11870
rect 15326 11868 15332 11870
rect 15396 11868 15402 11932
rect 0 11794 160 11824
rect 3233 11794 3299 11797
rect 0 11792 3299 11794
rect 0 11736 3238 11792
rect 3294 11736 3299 11792
rect 0 11734 3299 11736
rect 0 11704 160 11734
rect 3233 11731 3299 11734
rect 3417 11794 3483 11797
rect 18229 11794 18295 11797
rect 3417 11792 18295 11794
rect 3417 11736 3422 11792
rect 3478 11736 18234 11792
rect 18290 11736 18295 11792
rect 3417 11734 18295 11736
rect 3417 11731 3483 11734
rect 18229 11731 18295 11734
rect 3049 11658 3115 11661
rect 4889 11658 4955 11661
rect 3049 11656 4955 11658
rect 3049 11600 3054 11656
rect 3110 11600 4894 11656
rect 4950 11600 4955 11656
rect 3049 11598 4955 11600
rect 3049 11595 3115 11598
rect 4889 11595 4955 11598
rect 8017 11658 8083 11661
rect 19701 11658 19767 11661
rect 8017 11656 19767 11658
rect 8017 11600 8022 11656
rect 8078 11600 19706 11656
rect 19762 11600 19767 11656
rect 8017 11598 19767 11600
rect 8017 11595 8083 11598
rect 19701 11595 19767 11598
rect 0 11522 160 11552
rect 1945 11522 2011 11525
rect 0 11520 2011 11522
rect 0 11464 1950 11520
rect 2006 11464 2011 11520
rect 0 11462 2011 11464
rect 0 11432 160 11462
rect 1945 11459 2011 11462
rect 23841 11522 23907 11525
rect 25840 11522 26000 11552
rect 23841 11520 26000 11522
rect 23841 11464 23846 11520
rect 23902 11464 26000 11520
rect 23841 11462 26000 11464
rect 23841 11459 23907 11462
rect 3913 11456 4229 11457
rect 3913 11392 3919 11456
rect 3983 11392 3999 11456
rect 4063 11392 4079 11456
rect 4143 11392 4159 11456
rect 4223 11392 4229 11456
rect 3913 11391 4229 11392
rect 9847 11456 10163 11457
rect 9847 11392 9853 11456
rect 9917 11392 9933 11456
rect 9997 11392 10013 11456
rect 10077 11392 10093 11456
rect 10157 11392 10163 11456
rect 9847 11391 10163 11392
rect 15781 11456 16097 11457
rect 15781 11392 15787 11456
rect 15851 11392 15867 11456
rect 15931 11392 15947 11456
rect 16011 11392 16027 11456
rect 16091 11392 16097 11456
rect 15781 11391 16097 11392
rect 21715 11456 22031 11457
rect 21715 11392 21721 11456
rect 21785 11392 21801 11456
rect 21865 11392 21881 11456
rect 21945 11392 21961 11456
rect 22025 11392 22031 11456
rect 25840 11432 26000 11462
rect 21715 11391 22031 11392
rect 0 11250 160 11280
rect 3877 11250 3943 11253
rect 0 11248 3943 11250
rect 0 11192 3882 11248
rect 3938 11192 3943 11248
rect 0 11190 3943 11192
rect 0 11160 160 11190
rect 3877 11187 3943 11190
rect 5165 11250 5231 11253
rect 8334 11250 8340 11252
rect 5165 11248 8340 11250
rect 5165 11192 5170 11248
rect 5226 11192 8340 11248
rect 5165 11190 8340 11192
rect 5165 11187 5231 11190
rect 8334 11188 8340 11190
rect 8404 11188 8410 11252
rect 17033 11250 17099 11253
rect 12390 11248 17099 11250
rect 12390 11192 17038 11248
rect 17094 11192 17099 11248
rect 12390 11190 17099 11192
rect 3325 11114 3391 11117
rect 12390 11114 12450 11190
rect 17033 11187 17099 11190
rect 3325 11112 12450 11114
rect 3325 11056 3330 11112
rect 3386 11056 12450 11112
rect 3325 11054 12450 11056
rect 3325 11051 3391 11054
rect 0 10978 160 11008
rect 2221 10978 2287 10981
rect 0 10976 2287 10978
rect 0 10920 2226 10976
rect 2282 10920 2287 10976
rect 0 10918 2287 10920
rect 0 10888 160 10918
rect 2221 10915 2287 10918
rect 4337 10978 4403 10981
rect 4470 10978 4476 10980
rect 4337 10976 4476 10978
rect 4337 10920 4342 10976
rect 4398 10920 4476 10976
rect 4337 10918 4476 10920
rect 4337 10915 4403 10918
rect 4470 10916 4476 10918
rect 4540 10916 4546 10980
rect 25221 10978 25287 10981
rect 25840 10978 26000 11008
rect 25221 10976 26000 10978
rect 25221 10920 25226 10976
rect 25282 10920 26000 10976
rect 25221 10918 26000 10920
rect 25221 10915 25287 10918
rect 6880 10912 7196 10913
rect 6880 10848 6886 10912
rect 6950 10848 6966 10912
rect 7030 10848 7046 10912
rect 7110 10848 7126 10912
rect 7190 10848 7196 10912
rect 6880 10847 7196 10848
rect 12814 10912 13130 10913
rect 12814 10848 12820 10912
rect 12884 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13130 10912
rect 12814 10847 13130 10848
rect 18748 10912 19064 10913
rect 18748 10848 18754 10912
rect 18818 10848 18834 10912
rect 18898 10848 18914 10912
rect 18978 10848 18994 10912
rect 19058 10848 19064 10912
rect 18748 10847 19064 10848
rect 24682 10912 24998 10913
rect 24682 10848 24688 10912
rect 24752 10848 24768 10912
rect 24832 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 24998 10912
rect 25840 10888 26000 10918
rect 24682 10847 24998 10848
rect 0 10706 160 10736
rect 3969 10706 4035 10709
rect 0 10704 4035 10706
rect 0 10648 3974 10704
rect 4030 10648 4035 10704
rect 0 10646 4035 10648
rect 0 10616 160 10646
rect 3969 10643 4035 10646
rect 4061 10570 4127 10573
rect 11094 10570 11100 10572
rect 4061 10568 4354 10570
rect 4061 10512 4066 10568
rect 4122 10512 4354 10568
rect 4061 10510 4354 10512
rect 4061 10507 4127 10510
rect 0 10434 160 10464
rect 1669 10434 1735 10437
rect 0 10432 1735 10434
rect 0 10376 1674 10432
rect 1730 10376 1735 10432
rect 0 10374 1735 10376
rect 0 10344 160 10374
rect 1669 10371 1735 10374
rect 3913 10368 4229 10369
rect 3913 10304 3919 10368
rect 3983 10304 3999 10368
rect 4063 10304 4079 10368
rect 4143 10304 4159 10368
rect 4223 10304 4229 10368
rect 3913 10303 4229 10304
rect 3049 10300 3115 10301
rect 2998 10298 3004 10300
rect 2958 10238 3004 10298
rect 3068 10296 3115 10300
rect 3110 10240 3115 10296
rect 2998 10236 3004 10238
rect 3068 10236 3115 10240
rect 3049 10235 3115 10236
rect 0 10162 160 10192
rect 933 10162 999 10165
rect 2129 10164 2195 10165
rect 2078 10162 2084 10164
rect 0 10160 999 10162
rect 0 10104 938 10160
rect 994 10104 999 10160
rect 0 10102 999 10104
rect 2038 10102 2084 10162
rect 2148 10162 2195 10164
rect 3969 10162 4035 10165
rect 2148 10160 4035 10162
rect 2190 10104 3974 10160
rect 4030 10104 4035 10160
rect 0 10072 160 10102
rect 933 10099 999 10102
rect 2078 10100 2084 10102
rect 2148 10102 4035 10104
rect 2148 10100 2195 10102
rect 2129 10099 2195 10100
rect 3969 10099 4035 10102
rect 4153 10162 4219 10165
rect 4294 10162 4354 10510
rect 4153 10160 4354 10162
rect 4153 10104 4158 10160
rect 4214 10104 4354 10160
rect 4153 10102 4354 10104
rect 5398 10510 11100 10570
rect 4153 10099 4219 10102
rect 2865 10026 2931 10029
rect 4061 10026 4127 10029
rect 2865 10024 4127 10026
rect 2865 9968 2870 10024
rect 2926 9968 4066 10024
rect 4122 9968 4127 10024
rect 2865 9966 4127 9968
rect 2865 9963 2931 9966
rect 4061 9963 4127 9966
rect 0 9890 160 9920
rect 1393 9890 1459 9893
rect 0 9888 1459 9890
rect 0 9832 1398 9888
rect 1454 9832 1459 9888
rect 0 9830 1459 9832
rect 0 9800 160 9830
rect 1393 9827 1459 9830
rect 1894 9828 1900 9892
rect 1964 9890 1970 9892
rect 5073 9890 5139 9893
rect 1964 9888 5139 9890
rect 1964 9832 5078 9888
rect 5134 9832 5139 9888
rect 1964 9830 5139 9832
rect 1964 9828 1970 9830
rect 5073 9827 5139 9830
rect 2313 9754 2379 9757
rect 2681 9754 2747 9757
rect 2957 9756 3023 9757
rect 3141 9756 3207 9757
rect 2957 9754 3004 9756
rect 2313 9752 2747 9754
rect 2313 9696 2318 9752
rect 2374 9696 2686 9752
rect 2742 9696 2747 9752
rect 2313 9694 2747 9696
rect 2912 9752 3004 9754
rect 2912 9696 2962 9752
rect 2912 9694 3004 9696
rect 2313 9691 2379 9694
rect 2681 9691 2747 9694
rect 2957 9692 3004 9694
rect 3068 9692 3074 9756
rect 3141 9752 3188 9756
rect 3252 9754 3258 9756
rect 3601 9754 3667 9757
rect 5398 9754 5458 10510
rect 11094 10508 11100 10510
rect 11164 10508 11170 10572
rect 23289 10434 23355 10437
rect 25840 10434 26000 10464
rect 23289 10432 26000 10434
rect 23289 10376 23294 10432
rect 23350 10376 26000 10432
rect 23289 10374 26000 10376
rect 23289 10371 23355 10374
rect 9847 10368 10163 10369
rect 9847 10304 9853 10368
rect 9917 10304 9933 10368
rect 9997 10304 10013 10368
rect 10077 10304 10093 10368
rect 10157 10304 10163 10368
rect 9847 10303 10163 10304
rect 15781 10368 16097 10369
rect 15781 10304 15787 10368
rect 15851 10304 15867 10368
rect 15931 10304 15947 10368
rect 16011 10304 16027 10368
rect 16091 10304 16097 10368
rect 15781 10303 16097 10304
rect 21715 10368 22031 10369
rect 21715 10304 21721 10368
rect 21785 10304 21801 10368
rect 21865 10304 21881 10368
rect 21945 10304 21961 10368
rect 22025 10304 22031 10368
rect 25840 10344 26000 10374
rect 21715 10303 22031 10304
rect 10777 10298 10843 10301
rect 15193 10298 15259 10301
rect 10777 10296 15259 10298
rect 10777 10240 10782 10296
rect 10838 10240 15198 10296
rect 15254 10240 15259 10296
rect 10777 10238 15259 10240
rect 10777 10235 10843 10238
rect 15193 10235 15259 10238
rect 9765 10162 9831 10165
rect 10358 10162 10364 10164
rect 6134 10102 9322 10162
rect 5993 10026 6059 10029
rect 6134 10026 6194 10102
rect 5993 10024 6194 10026
rect 5993 9968 5998 10024
rect 6054 9968 6194 10024
rect 5993 9966 6194 9968
rect 6453 10026 6519 10029
rect 9070 10026 9076 10028
rect 6453 10024 9076 10026
rect 6453 9968 6458 10024
rect 6514 9968 9076 10024
rect 6453 9966 9076 9968
rect 5993 9963 6059 9966
rect 6453 9963 6519 9966
rect 9070 9964 9076 9966
rect 9140 9964 9146 10028
rect 9262 10026 9322 10102
rect 9765 10160 10364 10162
rect 9765 10104 9770 10160
rect 9826 10104 10364 10160
rect 9765 10102 10364 10104
rect 9765 10099 9831 10102
rect 10358 10100 10364 10102
rect 10428 10100 10434 10164
rect 10961 10162 11027 10165
rect 17309 10162 17375 10165
rect 10961 10160 17375 10162
rect 10961 10104 10966 10160
rect 11022 10104 17314 10160
rect 17370 10104 17375 10160
rect 10961 10102 17375 10104
rect 10961 10099 11027 10102
rect 17309 10099 17375 10102
rect 21582 10100 21588 10164
rect 21652 10162 21658 10164
rect 23197 10162 23263 10165
rect 21652 10160 23263 10162
rect 21652 10104 23202 10160
rect 23258 10104 23263 10160
rect 21652 10102 23263 10104
rect 21652 10100 21658 10102
rect 23197 10099 23263 10102
rect 11462 10026 11468 10028
rect 9262 9966 11468 10026
rect 11462 9964 11468 9966
rect 11532 9964 11538 10028
rect 13261 10026 13327 10029
rect 17585 10026 17651 10029
rect 13261 10024 17651 10026
rect 13261 9968 13266 10024
rect 13322 9968 17590 10024
rect 17646 9968 17651 10024
rect 13261 9966 17651 9968
rect 13261 9963 13327 9966
rect 17585 9963 17651 9966
rect 13629 9890 13695 9893
rect 14590 9890 14596 9892
rect 13629 9888 14596 9890
rect 13629 9832 13634 9888
rect 13690 9832 14596 9888
rect 13629 9830 14596 9832
rect 13629 9827 13695 9830
rect 14590 9828 14596 9830
rect 14660 9828 14666 9892
rect 25129 9890 25195 9893
rect 25840 9890 26000 9920
rect 25129 9888 26000 9890
rect 25129 9832 25134 9888
rect 25190 9832 26000 9888
rect 25129 9830 26000 9832
rect 25129 9827 25195 9830
rect 6880 9824 7196 9825
rect 6880 9760 6886 9824
rect 6950 9760 6966 9824
rect 7030 9760 7046 9824
rect 7110 9760 7126 9824
rect 7190 9760 7196 9824
rect 6880 9759 7196 9760
rect 12814 9824 13130 9825
rect 12814 9760 12820 9824
rect 12884 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13130 9824
rect 12814 9759 13130 9760
rect 18748 9824 19064 9825
rect 18748 9760 18754 9824
rect 18818 9760 18834 9824
rect 18898 9760 18914 9824
rect 18978 9760 18994 9824
rect 19058 9760 19064 9824
rect 18748 9759 19064 9760
rect 24682 9824 24998 9825
rect 24682 9760 24688 9824
rect 24752 9760 24768 9824
rect 24832 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 24998 9824
rect 25840 9800 26000 9830
rect 24682 9759 24998 9760
rect 3141 9696 3146 9752
rect 3141 9692 3188 9696
rect 3252 9694 3298 9754
rect 3601 9752 5458 9754
rect 3601 9696 3606 9752
rect 3662 9696 5458 9752
rect 3601 9694 5458 9696
rect 3252 9692 3258 9694
rect 2957 9691 3023 9692
rect 3141 9691 3207 9692
rect 3601 9691 3667 9694
rect 12198 9692 12204 9756
rect 12268 9754 12274 9756
rect 12341 9754 12407 9757
rect 12268 9752 12407 9754
rect 12268 9696 12346 9752
rect 12402 9696 12407 9752
rect 12268 9694 12407 9696
rect 12268 9692 12274 9694
rect 12341 9691 12407 9694
rect 13813 9754 13879 9757
rect 16798 9754 16804 9756
rect 13813 9752 16804 9754
rect 13813 9696 13818 9752
rect 13874 9696 16804 9752
rect 13813 9694 16804 9696
rect 13813 9691 13879 9694
rect 16798 9692 16804 9694
rect 16868 9692 16874 9756
rect 0 9618 160 9648
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 160 9558
rect 933 9555 999 9558
rect 1577 9618 1643 9621
rect 9305 9618 9371 9621
rect 1577 9616 9371 9618
rect 1577 9560 1582 9616
rect 1638 9560 9310 9616
rect 9366 9560 9371 9616
rect 1577 9558 9371 9560
rect 1577 9555 1643 9558
rect 9305 9555 9371 9558
rect 9673 9618 9739 9621
rect 15653 9618 15719 9621
rect 9673 9616 15719 9618
rect 9673 9560 9678 9616
rect 9734 9560 15658 9616
rect 15714 9560 15719 9616
rect 9673 9558 15719 9560
rect 9673 9555 9739 9558
rect 15653 9555 15719 9558
rect 2773 9482 2839 9485
rect 4337 9482 4403 9485
rect 2773 9480 4403 9482
rect 2773 9424 2778 9480
rect 2834 9424 4342 9480
rect 4398 9424 4403 9480
rect 2773 9422 4403 9424
rect 2773 9419 2839 9422
rect 4337 9419 4403 9422
rect 7833 9482 7899 9485
rect 9581 9482 9647 9485
rect 7833 9480 9647 9482
rect 7833 9424 7838 9480
rect 7894 9424 9586 9480
rect 9642 9424 9647 9480
rect 7833 9422 9647 9424
rect 7833 9419 7899 9422
rect 9581 9419 9647 9422
rect 11053 9482 11119 9485
rect 19742 9482 19748 9484
rect 11053 9480 19748 9482
rect 11053 9424 11058 9480
rect 11114 9424 19748 9480
rect 11053 9422 19748 9424
rect 11053 9419 11119 9422
rect 19742 9420 19748 9422
rect 19812 9420 19818 9484
rect 0 9346 160 9376
rect 2313 9346 2379 9349
rect 0 9344 2379 9346
rect 0 9288 2318 9344
rect 2374 9288 2379 9344
rect 0 9286 2379 9288
rect 0 9256 160 9286
rect 2313 9283 2379 9286
rect 24025 9346 24091 9349
rect 25840 9346 26000 9376
rect 24025 9344 26000 9346
rect 24025 9288 24030 9344
rect 24086 9288 26000 9344
rect 24025 9286 26000 9288
rect 24025 9283 24091 9286
rect 3913 9280 4229 9281
rect 3913 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4229 9280
rect 3913 9215 4229 9216
rect 9847 9280 10163 9281
rect 9847 9216 9853 9280
rect 9917 9216 9933 9280
rect 9997 9216 10013 9280
rect 10077 9216 10093 9280
rect 10157 9216 10163 9280
rect 9847 9215 10163 9216
rect 15781 9280 16097 9281
rect 15781 9216 15787 9280
rect 15851 9216 15867 9280
rect 15931 9216 15947 9280
rect 16011 9216 16027 9280
rect 16091 9216 16097 9280
rect 15781 9215 16097 9216
rect 21715 9280 22031 9281
rect 21715 9216 21721 9280
rect 21785 9216 21801 9280
rect 21865 9216 21881 9280
rect 21945 9216 21961 9280
rect 22025 9216 22031 9280
rect 25840 9256 26000 9286
rect 21715 9215 22031 9216
rect 0 9074 160 9104
rect 1209 9074 1275 9077
rect 0 9072 1275 9074
rect 0 9016 1214 9072
rect 1270 9016 1275 9072
rect 0 9014 1275 9016
rect 0 8984 160 9014
rect 1209 9011 1275 9014
rect 14917 9074 14983 9077
rect 15326 9074 15332 9076
rect 14917 9072 15332 9074
rect 14917 9016 14922 9072
rect 14978 9016 15332 9072
rect 14917 9014 15332 9016
rect 14917 9011 14983 9014
rect 15326 9012 15332 9014
rect 15396 9074 15402 9076
rect 15745 9074 15811 9077
rect 15396 9072 15811 9074
rect 15396 9016 15750 9072
rect 15806 9016 15811 9072
rect 15396 9014 15811 9016
rect 15396 9012 15402 9014
rect 15745 9011 15811 9014
rect 1485 8938 1551 8941
rect 3049 8938 3115 8941
rect 1485 8936 3115 8938
rect 1485 8880 1490 8936
rect 1546 8880 3054 8936
rect 3110 8880 3115 8936
rect 1485 8878 3115 8880
rect 1485 8875 1551 8878
rect 3049 8875 3115 8878
rect 8937 8938 9003 8941
rect 9397 8938 9463 8941
rect 14365 8938 14431 8941
rect 8937 8936 14431 8938
rect 8937 8880 8942 8936
rect 8998 8880 9402 8936
rect 9458 8880 14370 8936
rect 14426 8880 14431 8936
rect 8937 8878 14431 8880
rect 8937 8875 9003 8878
rect 9397 8875 9463 8878
rect 14365 8875 14431 8878
rect 23565 8938 23631 8941
rect 23565 8936 25146 8938
rect 23565 8880 23570 8936
rect 23626 8880 25146 8936
rect 23565 8878 25146 8880
rect 23565 8875 23631 8878
rect 0 8802 160 8832
rect 1761 8802 1827 8805
rect 0 8800 1827 8802
rect 0 8744 1766 8800
rect 1822 8744 1827 8800
rect 0 8742 1827 8744
rect 25086 8802 25146 8878
rect 25840 8802 26000 8832
rect 25086 8742 26000 8802
rect 0 8712 160 8742
rect 1761 8739 1827 8742
rect 6880 8736 7196 8737
rect 6880 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7196 8736
rect 6880 8671 7196 8672
rect 12814 8736 13130 8737
rect 12814 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13130 8736
rect 12814 8671 13130 8672
rect 18748 8736 19064 8737
rect 18748 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19064 8736
rect 18748 8671 19064 8672
rect 24682 8736 24998 8737
rect 24682 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 24998 8736
rect 25840 8712 26000 8742
rect 24682 8671 24998 8672
rect 0 8530 160 8560
rect 1301 8530 1367 8533
rect 0 8528 1367 8530
rect 0 8472 1306 8528
rect 1362 8472 1367 8528
rect 0 8470 1367 8472
rect 0 8440 160 8470
rect 1301 8467 1367 8470
rect 3734 8468 3740 8532
rect 3804 8530 3810 8532
rect 9438 8530 9444 8532
rect 3804 8470 9444 8530
rect 3804 8468 3810 8470
rect 9438 8468 9444 8470
rect 9508 8468 9514 8532
rect 10961 8530 11027 8533
rect 18321 8530 18387 8533
rect 10961 8528 18387 8530
rect 10961 8472 10966 8528
rect 11022 8472 18326 8528
rect 18382 8472 18387 8528
rect 10961 8470 18387 8472
rect 10961 8467 11027 8470
rect 18321 8467 18387 8470
rect 8753 8394 8819 8397
rect 9070 8394 9076 8396
rect 8753 8392 9076 8394
rect 8753 8336 8758 8392
rect 8814 8336 9076 8392
rect 8753 8334 9076 8336
rect 8753 8331 8819 8334
rect 9070 8332 9076 8334
rect 9140 8332 9146 8396
rect 11973 8394 12039 8397
rect 19558 8394 19564 8396
rect 11973 8392 19564 8394
rect 11973 8336 11978 8392
rect 12034 8336 19564 8392
rect 11973 8334 19564 8336
rect 11973 8331 12039 8334
rect 19558 8332 19564 8334
rect 19628 8332 19634 8396
rect 19885 8394 19951 8397
rect 20478 8394 20484 8396
rect 19885 8392 20484 8394
rect 19885 8336 19890 8392
rect 19946 8336 20484 8392
rect 19885 8334 20484 8336
rect 19885 8331 19951 8334
rect 20478 8332 20484 8334
rect 20548 8332 20554 8396
rect 0 8258 160 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 160 8198
rect 1577 8195 1643 8198
rect 24485 8258 24551 8261
rect 25840 8258 26000 8288
rect 24485 8256 26000 8258
rect 24485 8200 24490 8256
rect 24546 8200 26000 8256
rect 24485 8198 26000 8200
rect 24485 8195 24551 8198
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 9847 8192 10163 8193
rect 9847 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10163 8192
rect 9847 8127 10163 8128
rect 15781 8192 16097 8193
rect 15781 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16097 8192
rect 15781 8127 16097 8128
rect 21715 8192 22031 8193
rect 21715 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22031 8192
rect 25840 8168 26000 8198
rect 21715 8127 22031 8128
rect 0 7986 160 8016
rect 3325 7986 3391 7989
rect 0 7984 3391 7986
rect 0 7928 3330 7984
rect 3386 7928 3391 7984
rect 0 7926 3391 7928
rect 0 7896 160 7926
rect 3325 7923 3391 7926
rect 7189 7986 7255 7989
rect 8109 7986 8175 7989
rect 7189 7984 8175 7986
rect 7189 7928 7194 7984
rect 7250 7928 8114 7984
rect 8170 7928 8175 7984
rect 7189 7926 8175 7928
rect 7189 7923 7255 7926
rect 8109 7923 8175 7926
rect 9765 7986 9831 7989
rect 16205 7986 16271 7989
rect 9765 7984 16271 7986
rect 9765 7928 9770 7984
rect 9826 7928 16210 7984
rect 16266 7928 16271 7984
rect 9765 7926 16271 7928
rect 9765 7923 9831 7926
rect 16205 7923 16271 7926
rect 2221 7850 2287 7853
rect 9029 7850 9095 7853
rect 2221 7848 9095 7850
rect 2221 7792 2226 7848
rect 2282 7792 9034 7848
rect 9090 7792 9095 7848
rect 2221 7790 9095 7792
rect 2221 7787 2287 7790
rect 9029 7787 9095 7790
rect 21541 7850 21607 7853
rect 21541 7848 25146 7850
rect 21541 7792 21546 7848
rect 21602 7792 25146 7848
rect 21541 7790 25146 7792
rect 21541 7787 21607 7790
rect 0 7714 160 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 160 7654
rect 1393 7651 1459 7654
rect 2630 7652 2636 7716
rect 2700 7714 2706 7716
rect 5717 7714 5783 7717
rect 2700 7712 5783 7714
rect 2700 7656 5722 7712
rect 5778 7656 5783 7712
rect 2700 7654 5783 7656
rect 2700 7652 2706 7654
rect 5717 7651 5783 7654
rect 15510 7652 15516 7716
rect 15580 7714 15586 7716
rect 15653 7714 15719 7717
rect 15580 7712 15719 7714
rect 15580 7656 15658 7712
rect 15714 7656 15719 7712
rect 15580 7654 15719 7656
rect 25086 7714 25146 7790
rect 25840 7714 26000 7744
rect 25086 7654 26000 7714
rect 15580 7652 15586 7654
rect 15653 7651 15719 7654
rect 6880 7648 7196 7649
rect 6880 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7196 7648
rect 6880 7583 7196 7584
rect 12814 7648 13130 7649
rect 12814 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13130 7648
rect 12814 7583 13130 7584
rect 18748 7648 19064 7649
rect 18748 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19064 7648
rect 18748 7583 19064 7584
rect 24682 7648 24998 7649
rect 24682 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 24998 7648
rect 25840 7624 26000 7654
rect 24682 7583 24998 7584
rect 20437 7578 20503 7581
rect 20437 7576 20546 7578
rect 20437 7520 20442 7576
rect 20498 7520 20546 7576
rect 20437 7515 20546 7520
rect 0 7442 160 7472
rect 1761 7442 1827 7445
rect 0 7440 1827 7442
rect 0 7384 1766 7440
rect 1822 7384 1827 7440
rect 0 7382 1827 7384
rect 20486 7442 20546 7515
rect 20621 7442 20687 7445
rect 20486 7440 20687 7442
rect 20486 7384 20626 7440
rect 20682 7384 20687 7440
rect 20486 7382 20687 7384
rect 0 7352 160 7382
rect 1761 7379 1827 7382
rect 20621 7379 20687 7382
rect 4337 7306 4403 7309
rect 6085 7306 6151 7309
rect 4337 7304 6151 7306
rect 4337 7248 4342 7304
rect 4398 7248 6090 7304
rect 6146 7248 6151 7304
rect 4337 7246 6151 7248
rect 4337 7243 4403 7246
rect 6085 7243 6151 7246
rect 0 7170 160 7200
rect 2129 7170 2195 7173
rect 0 7168 2195 7170
rect 0 7112 2134 7168
rect 2190 7112 2195 7168
rect 0 7110 2195 7112
rect 0 7080 160 7110
rect 2129 7107 2195 7110
rect 23749 7170 23815 7173
rect 25840 7170 26000 7200
rect 23749 7168 26000 7170
rect 23749 7112 23754 7168
rect 23810 7112 26000 7168
rect 23749 7110 26000 7112
rect 23749 7107 23815 7110
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 9847 7104 10163 7105
rect 9847 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10163 7104
rect 9847 7039 10163 7040
rect 15781 7104 16097 7105
rect 15781 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16097 7104
rect 15781 7039 16097 7040
rect 21715 7104 22031 7105
rect 21715 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22031 7104
rect 25840 7080 26000 7110
rect 21715 7039 22031 7040
rect 11237 7034 11303 7037
rect 15285 7034 15351 7037
rect 11237 7032 15351 7034
rect 11237 6976 11242 7032
rect 11298 6976 15290 7032
rect 15346 6976 15351 7032
rect 11237 6974 15351 6976
rect 11237 6971 11303 6974
rect 15285 6971 15351 6974
rect 0 6898 160 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 160 6838
rect 1209 6835 1275 6838
rect 3601 6898 3667 6901
rect 8569 6898 8635 6901
rect 3601 6896 8635 6898
rect 3601 6840 3606 6896
rect 3662 6840 8574 6896
rect 8630 6840 8635 6896
rect 3601 6838 8635 6840
rect 3601 6835 3667 6838
rect 8569 6835 8635 6838
rect 16665 6898 16731 6901
rect 21265 6898 21331 6901
rect 16665 6896 21331 6898
rect 16665 6840 16670 6896
rect 16726 6840 21270 6896
rect 21326 6840 21331 6896
rect 16665 6838 21331 6840
rect 16665 6835 16731 6838
rect 21265 6835 21331 6838
rect 21725 6898 21791 6901
rect 25497 6898 25563 6901
rect 21725 6896 25563 6898
rect 21725 6840 21730 6896
rect 21786 6840 25502 6896
rect 25558 6840 25563 6896
rect 21725 6838 25563 6840
rect 21725 6835 21791 6838
rect 25497 6835 25563 6838
rect 23197 6762 23263 6765
rect 12390 6760 23263 6762
rect 12390 6704 23202 6760
rect 23258 6704 23263 6760
rect 12390 6702 23263 6704
rect 0 6626 160 6656
rect 1025 6626 1091 6629
rect 0 6624 1091 6626
rect 0 6568 1030 6624
rect 1086 6568 1091 6624
rect 0 6566 1091 6568
rect 0 6536 160 6566
rect 1025 6563 1091 6566
rect 2589 6626 2655 6629
rect 2957 6626 3023 6629
rect 2589 6624 3023 6626
rect 2589 6568 2594 6624
rect 2650 6568 2962 6624
rect 3018 6568 3023 6624
rect 2589 6566 3023 6568
rect 2589 6563 2655 6566
rect 0 6354 160 6384
rect 1301 6354 1367 6357
rect 0 6352 1367 6354
rect 0 6296 1306 6352
rect 1362 6296 1367 6352
rect 0 6294 1367 6296
rect 2730 6354 2790 6566
rect 2957 6563 3023 6566
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 2957 6490 3023 6493
rect 5717 6490 5783 6493
rect 12390 6490 12450 6702
rect 23197 6699 23263 6702
rect 24534 6702 25146 6762
rect 20713 6626 20779 6629
rect 24534 6626 24594 6702
rect 20713 6624 24594 6626
rect 20713 6568 20718 6624
rect 20774 6568 24594 6624
rect 20713 6566 24594 6568
rect 25086 6626 25146 6702
rect 25840 6626 26000 6656
rect 25086 6566 26000 6626
rect 20713 6563 20779 6566
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 25840 6536 26000 6566
rect 24682 6495 24998 6496
rect 2957 6488 5783 6490
rect 2957 6432 2962 6488
rect 3018 6432 5722 6488
rect 5778 6432 5783 6488
rect 2957 6430 5783 6432
rect 2957 6427 3023 6430
rect 5717 6427 5783 6430
rect 7284 6430 12450 6490
rect 19425 6490 19491 6493
rect 19425 6488 21972 6490
rect 19425 6432 19430 6488
rect 19486 6432 21972 6488
rect 19425 6430 21972 6432
rect 7284 6354 7344 6430
rect 19425 6427 19491 6430
rect 2730 6294 7344 6354
rect 0 6264 160 6294
rect 1301 6291 1367 6294
rect 10910 6292 10916 6356
rect 10980 6354 10986 6356
rect 13721 6354 13787 6357
rect 10980 6352 13787 6354
rect 10980 6296 13726 6352
rect 13782 6296 13787 6352
rect 10980 6294 13787 6296
rect 10980 6292 10986 6294
rect 13721 6291 13787 6294
rect 15561 6354 15627 6357
rect 21725 6354 21791 6357
rect 15561 6352 21791 6354
rect 15561 6296 15566 6352
rect 15622 6296 21730 6352
rect 21786 6296 21791 6352
rect 15561 6294 21791 6296
rect 21912 6354 21972 6430
rect 22318 6354 22324 6356
rect 21912 6294 22324 6354
rect 15561 6291 15627 6294
rect 21725 6291 21791 6294
rect 22318 6292 22324 6294
rect 22388 6292 22394 6356
rect 2957 6218 3023 6221
rect 3550 6218 3556 6220
rect 2957 6216 3556 6218
rect 2957 6160 2962 6216
rect 3018 6160 3556 6216
rect 2957 6158 3556 6160
rect 2957 6155 3023 6158
rect 3550 6156 3556 6158
rect 3620 6218 3626 6220
rect 5165 6218 5231 6221
rect 13353 6218 13419 6221
rect 19425 6218 19491 6221
rect 3620 6158 4354 6218
rect 3620 6156 3626 6158
rect 0 6082 160 6112
rect 4294 6082 4354 6158
rect 5165 6216 13419 6218
rect 5165 6160 5170 6216
rect 5226 6160 13358 6216
rect 13414 6160 13419 6216
rect 5165 6158 13419 6160
rect 5165 6155 5231 6158
rect 13353 6155 13419 6158
rect 13494 6216 19491 6218
rect 13494 6160 19430 6216
rect 19486 6160 19491 6216
rect 13494 6158 19491 6160
rect 13494 6085 13554 6158
rect 19425 6155 19491 6158
rect 20253 6218 20319 6221
rect 20253 6216 24042 6218
rect 20253 6160 20258 6216
rect 20314 6160 24042 6216
rect 20253 6158 24042 6160
rect 20253 6155 20319 6158
rect 9305 6082 9371 6085
rect 0 6022 1640 6082
rect 4294 6080 9371 6082
rect 4294 6024 9310 6080
rect 9366 6024 9371 6080
rect 4294 6022 9371 6024
rect 0 5992 160 6022
rect 0 5810 160 5840
rect 1301 5810 1367 5813
rect 0 5808 1367 5810
rect 0 5752 1306 5808
rect 1362 5752 1367 5808
rect 0 5750 1367 5752
rect 0 5720 160 5750
rect 1301 5747 1367 5750
rect 1580 5677 1640 6022
rect 9305 6019 9371 6022
rect 13445 6080 13554 6085
rect 13445 6024 13450 6080
rect 13506 6024 13554 6080
rect 13445 6022 13554 6024
rect 20621 6082 20687 6085
rect 21541 6082 21607 6085
rect 20621 6080 21607 6082
rect 20621 6024 20626 6080
rect 20682 6024 21546 6080
rect 21602 6024 21607 6080
rect 20621 6022 21607 6024
rect 23982 6082 24042 6158
rect 25840 6082 26000 6112
rect 23982 6022 26000 6082
rect 13445 6019 13511 6022
rect 20621 6019 20687 6022
rect 21541 6019 21607 6022
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 25840 5992 26000 6022
rect 21715 5951 22031 5952
rect 10961 5946 11027 5949
rect 14733 5946 14799 5949
rect 10961 5944 14799 5946
rect 10961 5888 10966 5944
rect 11022 5888 14738 5944
rect 14794 5888 14799 5944
rect 10961 5886 14799 5888
rect 10961 5883 11027 5886
rect 14733 5883 14799 5886
rect 3417 5810 3483 5813
rect 10501 5810 10567 5813
rect 17493 5810 17559 5813
rect 3417 5808 10567 5810
rect 3417 5752 3422 5808
rect 3478 5752 10506 5808
rect 10562 5752 10567 5808
rect 3417 5750 10567 5752
rect 3417 5747 3483 5750
rect 10501 5747 10567 5750
rect 12390 5808 17559 5810
rect 12390 5752 17498 5808
rect 17554 5752 17559 5808
rect 12390 5750 17559 5752
rect 1577 5672 1643 5677
rect 1577 5616 1582 5672
rect 1638 5616 1643 5672
rect 1577 5611 1643 5616
rect 5441 5674 5507 5677
rect 9673 5674 9739 5677
rect 12390 5674 12450 5750
rect 17493 5747 17559 5750
rect 21173 5810 21239 5813
rect 25037 5810 25103 5813
rect 21173 5808 25103 5810
rect 21173 5752 21178 5808
rect 21234 5752 25042 5808
rect 25098 5752 25103 5808
rect 21173 5750 25103 5752
rect 21173 5747 21239 5750
rect 25037 5747 25103 5750
rect 5441 5672 9739 5674
rect 5441 5616 5446 5672
rect 5502 5616 9678 5672
rect 9734 5616 9739 5672
rect 5441 5614 9739 5616
rect 5441 5611 5507 5614
rect 9673 5611 9739 5614
rect 9814 5614 12450 5674
rect 16389 5674 16455 5677
rect 23013 5674 23079 5677
rect 16389 5672 23079 5674
rect 16389 5616 16394 5672
rect 16450 5616 23018 5672
rect 23074 5616 23079 5672
rect 16389 5614 23079 5616
rect 0 5538 160 5568
rect 4797 5540 4863 5541
rect 0 5478 1042 5538
rect 0 5448 160 5478
rect 982 5402 1042 5478
rect 4797 5536 4844 5540
rect 4908 5538 4914 5540
rect 9305 5538 9371 5541
rect 9814 5538 9874 5614
rect 16389 5611 16455 5614
rect 23013 5611 23079 5614
rect 4797 5480 4802 5536
rect 4797 5476 4844 5480
rect 4908 5478 4954 5538
rect 9305 5536 9874 5538
rect 9305 5480 9310 5536
rect 9366 5480 9874 5536
rect 9305 5478 9874 5480
rect 13721 5538 13787 5541
rect 17401 5538 17467 5541
rect 13721 5536 17467 5538
rect 13721 5480 13726 5536
rect 13782 5480 17406 5536
rect 17462 5480 17467 5536
rect 13721 5478 17467 5480
rect 4908 5476 4914 5478
rect 4797 5475 4863 5476
rect 9305 5475 9371 5478
rect 13721 5475 13787 5478
rect 17401 5475 17467 5478
rect 20345 5538 20411 5541
rect 22553 5538 22619 5541
rect 25840 5538 26000 5568
rect 20345 5536 22619 5538
rect 20345 5480 20350 5536
rect 20406 5480 22558 5536
rect 22614 5480 22619 5536
rect 20345 5478 22619 5480
rect 20345 5475 20411 5478
rect 22553 5475 22619 5478
rect 25086 5478 26000 5538
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 1945 5402 2011 5405
rect 982 5400 2011 5402
rect 982 5344 1950 5400
rect 2006 5344 2011 5400
rect 982 5342 2011 5344
rect 1945 5339 2011 5342
rect 20529 5400 20595 5405
rect 20529 5344 20534 5400
rect 20590 5344 20595 5400
rect 20529 5339 20595 5344
rect 0 5266 160 5296
rect 2865 5266 2931 5269
rect 0 5264 2931 5266
rect 0 5208 2870 5264
rect 2926 5208 2931 5264
rect 0 5206 2931 5208
rect 0 5176 160 5206
rect 2865 5203 2931 5206
rect 4613 5266 4679 5269
rect 13445 5266 13511 5269
rect 13813 5266 13879 5269
rect 4613 5264 13879 5266
rect 4613 5208 4618 5264
rect 4674 5208 13450 5264
rect 13506 5208 13818 5264
rect 13874 5208 13879 5264
rect 4613 5206 13879 5208
rect 4613 5203 4679 5206
rect 13445 5203 13511 5206
rect 13813 5203 13879 5206
rect 17217 5266 17283 5269
rect 18689 5266 18755 5269
rect 17217 5264 18755 5266
rect 17217 5208 17222 5264
rect 17278 5208 18694 5264
rect 18750 5208 18755 5264
rect 17217 5206 18755 5208
rect 20532 5266 20592 5339
rect 25086 5266 25146 5478
rect 25840 5448 26000 5478
rect 20532 5206 25146 5266
rect 17217 5203 17283 5206
rect 18689 5203 18755 5206
rect 4245 5130 4311 5133
rect 15193 5130 15259 5133
rect 4245 5128 15259 5130
rect 4245 5072 4250 5128
rect 4306 5072 15198 5128
rect 15254 5072 15259 5128
rect 4245 5070 15259 5072
rect 4245 5067 4311 5070
rect 15193 5067 15259 5070
rect 20713 5130 20779 5133
rect 20713 5128 24042 5130
rect 20713 5072 20718 5128
rect 20774 5072 24042 5128
rect 20713 5070 24042 5072
rect 20713 5067 20779 5070
rect 0 4994 160 5024
rect 2129 4994 2195 4997
rect 0 4992 2195 4994
rect 0 4936 2134 4992
rect 2190 4936 2195 4992
rect 0 4934 2195 4936
rect 0 4904 160 4934
rect 2129 4931 2195 4934
rect 13077 4994 13143 4997
rect 14917 4994 14983 4997
rect 13077 4992 14983 4994
rect 13077 4936 13082 4992
rect 13138 4936 14922 4992
rect 14978 4936 14983 4992
rect 13077 4934 14983 4936
rect 23982 4994 24042 5070
rect 25840 4994 26000 5024
rect 23982 4934 26000 4994
rect 13077 4931 13143 4934
rect 14917 4931 14983 4934
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 25840 4904 26000 4934
rect 21715 4863 22031 4864
rect 17033 4860 17099 4861
rect 16982 4796 16988 4860
rect 17052 4858 17099 4860
rect 19333 4858 19399 4861
rect 21449 4858 21515 4861
rect 17052 4856 17144 4858
rect 17094 4800 17144 4856
rect 17052 4798 17144 4800
rect 19333 4856 21515 4858
rect 19333 4800 19338 4856
rect 19394 4800 21454 4856
rect 21510 4800 21515 4856
rect 19333 4798 21515 4800
rect 17052 4796 17099 4798
rect 17033 4795 17099 4796
rect 19333 4795 19399 4798
rect 21449 4795 21515 4798
rect 790 4660 796 4724
rect 860 4722 866 4724
rect 4521 4722 4587 4725
rect 860 4720 4587 4722
rect 860 4664 4526 4720
rect 4582 4664 4587 4720
rect 860 4662 4587 4664
rect 860 4660 866 4662
rect 4521 4659 4587 4662
rect 9213 4722 9279 4725
rect 14365 4722 14431 4725
rect 9213 4720 14431 4722
rect 9213 4664 9218 4720
rect 9274 4664 14370 4720
rect 14426 4664 14431 4720
rect 9213 4662 14431 4664
rect 9213 4659 9279 4662
rect 14365 4659 14431 4662
rect 19885 4722 19951 4725
rect 22001 4722 22067 4725
rect 19885 4720 22067 4722
rect 19885 4664 19890 4720
rect 19946 4664 22006 4720
rect 22062 4664 22067 4720
rect 19885 4662 22067 4664
rect 19885 4659 19951 4662
rect 22001 4659 22067 4662
rect 3969 4586 4035 4589
rect 8017 4586 8083 4589
rect 3969 4584 8083 4586
rect 3969 4528 3974 4584
rect 4030 4528 8022 4584
rect 8078 4528 8083 4584
rect 3969 4526 8083 4528
rect 3969 4523 4035 4526
rect 8017 4523 8083 4526
rect 11421 4586 11487 4589
rect 14917 4586 14983 4589
rect 11421 4584 14983 4586
rect 11421 4528 11426 4584
rect 11482 4528 14922 4584
rect 14978 4528 14983 4584
rect 11421 4526 14983 4528
rect 11421 4523 11487 4526
rect 14917 4523 14983 4526
rect 21265 4586 21331 4589
rect 21265 4584 25146 4586
rect 21265 4528 21270 4584
rect 21326 4528 25146 4584
rect 21265 4526 25146 4528
rect 21265 4523 21331 4526
rect 606 4388 612 4452
rect 676 4450 682 4452
rect 4889 4450 4955 4453
rect 676 4448 4955 4450
rect 676 4392 4894 4448
rect 4950 4392 4955 4448
rect 676 4390 4955 4392
rect 25086 4450 25146 4526
rect 25840 4450 26000 4480
rect 25086 4390 26000 4450
rect 676 4388 682 4390
rect 4889 4387 4955 4390
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 25840 4360 26000 4390
rect 24682 4319 24998 4320
rect 2313 4178 2379 4181
rect 3141 4178 3207 4181
rect 13169 4178 13235 4181
rect 2313 4176 9690 4178
rect 2313 4120 2318 4176
rect 2374 4120 3146 4176
rect 3202 4120 9690 4176
rect 2313 4118 9690 4120
rect 2313 4115 2379 4118
rect 3141 4115 3207 4118
rect 974 3980 980 4044
rect 1044 4042 1050 4044
rect 3325 4042 3391 4045
rect 1044 4040 3391 4042
rect 1044 3984 3330 4040
rect 3386 3984 3391 4040
rect 1044 3982 3391 3984
rect 9630 4042 9690 4118
rect 13169 4176 21282 4178
rect 13169 4120 13174 4176
rect 13230 4120 21282 4176
rect 13169 4118 21282 4120
rect 13169 4115 13235 4118
rect 11513 4042 11579 4045
rect 11789 4044 11855 4045
rect 11646 4042 11652 4044
rect 9630 3982 10426 4042
rect 1044 3980 1050 3982
rect 3325 3979 3391 3982
rect 10366 3906 10426 3982
rect 11513 4040 11652 4042
rect 11513 3984 11518 4040
rect 11574 3984 11652 4040
rect 11513 3982 11652 3984
rect 11513 3979 11579 3982
rect 11646 3980 11652 3982
rect 11716 3980 11722 4044
rect 11789 4040 11836 4044
rect 11900 4042 11906 4044
rect 21081 4042 21147 4045
rect 11789 3984 11794 4040
rect 11789 3980 11836 3984
rect 11900 3982 11946 4042
rect 12022 4040 21147 4042
rect 12022 3984 21086 4040
rect 21142 3984 21147 4040
rect 12022 3982 21147 3984
rect 21222 4042 21282 4118
rect 21633 4044 21699 4045
rect 21582 4042 21588 4044
rect 21222 3982 21588 4042
rect 21652 4040 21699 4044
rect 21694 3984 21699 4040
rect 11900 3980 11906 3982
rect 11789 3979 11855 3980
rect 12022 3906 12082 3982
rect 21081 3979 21147 3982
rect 21582 3980 21588 3982
rect 21652 3980 21699 3984
rect 21633 3979 21699 3980
rect 21817 4042 21883 4045
rect 21817 4040 24042 4042
rect 21817 3984 21822 4040
rect 21878 3984 24042 4040
rect 21817 3982 24042 3984
rect 21817 3979 21883 3982
rect 10366 3846 12082 3906
rect 12198 3844 12204 3908
rect 12268 3906 12274 3908
rect 12341 3906 12407 3909
rect 12268 3904 12407 3906
rect 12268 3848 12346 3904
rect 12402 3848 12407 3904
rect 12268 3846 12407 3848
rect 12268 3844 12274 3846
rect 12341 3843 12407 3846
rect 17217 3906 17283 3909
rect 17677 3908 17743 3909
rect 17350 3906 17356 3908
rect 17217 3904 17356 3906
rect 17217 3848 17222 3904
rect 17278 3848 17356 3904
rect 17217 3846 17356 3848
rect 17217 3843 17283 3846
rect 17350 3844 17356 3846
rect 17420 3844 17426 3908
rect 17677 3904 17724 3908
rect 17788 3906 17794 3908
rect 17953 3906 18019 3909
rect 18505 3908 18571 3909
rect 18086 3906 18092 3908
rect 17677 3848 17682 3904
rect 17677 3844 17724 3848
rect 17788 3846 17834 3906
rect 17953 3904 18092 3906
rect 17953 3848 17958 3904
rect 18014 3848 18092 3904
rect 17953 3846 18092 3848
rect 17788 3844 17794 3846
rect 17677 3843 17743 3844
rect 17953 3843 18019 3846
rect 18086 3844 18092 3846
rect 18156 3844 18162 3908
rect 18454 3906 18460 3908
rect 18414 3846 18460 3906
rect 18524 3904 18571 3908
rect 18566 3848 18571 3904
rect 18454 3844 18460 3846
rect 18524 3844 18571 3848
rect 23982 3906 24042 3982
rect 25840 3906 26000 3936
rect 23982 3846 26000 3906
rect 18505 3843 18571 3844
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 25840 3816 26000 3846
rect 21715 3775 22031 3776
rect 6361 3770 6427 3773
rect 9673 3770 9739 3773
rect 6361 3768 9739 3770
rect 6361 3712 6366 3768
rect 6422 3712 9678 3768
rect 9734 3712 9739 3768
rect 6361 3710 9739 3712
rect 6361 3707 6427 3710
rect 9673 3707 9739 3710
rect 11053 3770 11119 3773
rect 12893 3770 12959 3773
rect 20294 3770 20300 3772
rect 11053 3768 12959 3770
rect 11053 3712 11058 3768
rect 11114 3712 12898 3768
rect 12954 3712 12959 3768
rect 11053 3710 12959 3712
rect 11053 3707 11119 3710
rect 12893 3707 12959 3710
rect 16254 3710 20300 3770
rect 9029 3634 9095 3637
rect 16254 3634 16314 3710
rect 20294 3708 20300 3710
rect 20364 3708 20370 3772
rect 22369 3770 22435 3773
rect 25221 3770 25287 3773
rect 22369 3768 25287 3770
rect 22369 3712 22374 3768
rect 22430 3712 25226 3768
rect 25282 3712 25287 3768
rect 22369 3710 25287 3712
rect 22369 3707 22435 3710
rect 25221 3707 25287 3710
rect 25589 3634 25655 3637
rect 9029 3632 16314 3634
rect 9029 3576 9034 3632
rect 9090 3576 16314 3632
rect 9029 3574 16314 3576
rect 17174 3632 25655 3634
rect 17174 3576 25594 3632
rect 25650 3576 25655 3632
rect 17174 3574 25655 3576
rect 9029 3571 9095 3574
rect 6177 3498 6243 3501
rect 9949 3498 10015 3501
rect 17174 3498 17234 3574
rect 25589 3571 25655 3574
rect 6177 3496 9506 3498
rect 6177 3440 6182 3496
rect 6238 3440 9506 3496
rect 6177 3438 9506 3440
rect 6177 3435 6243 3438
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 9446 3226 9506 3438
rect 9949 3496 17234 3498
rect 9949 3440 9954 3496
rect 10010 3440 17234 3496
rect 9949 3438 17234 3440
rect 21173 3498 21239 3501
rect 23749 3498 23815 3501
rect 21173 3496 23815 3498
rect 21173 3440 21178 3496
rect 21234 3440 23754 3496
rect 23810 3440 23815 3496
rect 21173 3438 23815 3440
rect 9949 3435 10015 3438
rect 21173 3435 21239 3438
rect 23749 3435 23815 3438
rect 24350 3438 25146 3498
rect 9673 3362 9739 3365
rect 10685 3362 10751 3365
rect 9673 3360 10751 3362
rect 9673 3304 9678 3360
rect 9734 3304 10690 3360
rect 10746 3304 10751 3360
rect 9673 3302 10751 3304
rect 9673 3299 9739 3302
rect 10685 3299 10751 3302
rect 20713 3362 20779 3365
rect 24350 3362 24410 3438
rect 20713 3360 24410 3362
rect 20713 3304 20718 3360
rect 20774 3304 24410 3360
rect 20713 3302 24410 3304
rect 25086 3362 25146 3438
rect 25840 3362 26000 3392
rect 25086 3302 26000 3362
rect 20713 3299 20779 3302
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 25840 3272 26000 3302
rect 24682 3231 24998 3232
rect 11421 3226 11487 3229
rect 22502 3226 22508 3228
rect 9446 3224 11487 3226
rect 9446 3168 11426 3224
rect 11482 3168 11487 3224
rect 9446 3166 11487 3168
rect 11421 3163 11487 3166
rect 19198 3166 22508 3226
rect 3141 3090 3207 3093
rect 11053 3090 11119 3093
rect 3141 3088 11119 3090
rect 3141 3032 3146 3088
rect 3202 3032 11058 3088
rect 11114 3032 11119 3088
rect 3141 3030 11119 3032
rect 3141 3027 3207 3030
rect 11053 3027 11119 3030
rect 17585 3090 17651 3093
rect 19198 3090 19258 3166
rect 22502 3164 22508 3166
rect 22572 3164 22578 3228
rect 17585 3088 19258 3090
rect 17585 3032 17590 3088
rect 17646 3032 19258 3088
rect 17585 3030 19258 3032
rect 19977 3090 20043 3093
rect 24025 3090 24091 3093
rect 19977 3088 24091 3090
rect 19977 3032 19982 3088
rect 20038 3032 24030 3088
rect 24086 3032 24091 3088
rect 19977 3030 24091 3032
rect 17585 3027 17651 3030
rect 19977 3027 20043 3030
rect 24025 3027 24091 3030
rect 6545 2954 6611 2957
rect 6821 2954 6887 2957
rect 11881 2954 11947 2957
rect 6545 2952 6887 2954
rect 6545 2896 6550 2952
rect 6606 2896 6826 2952
rect 6882 2896 6887 2952
rect 6545 2894 6887 2896
rect 6545 2891 6611 2894
rect 6821 2891 6887 2894
rect 7054 2952 11947 2954
rect 7054 2896 11886 2952
rect 11942 2896 11947 2952
rect 7054 2894 11947 2896
rect 6269 2818 6335 2821
rect 7054 2818 7114 2894
rect 11881 2891 11947 2894
rect 20713 2954 20779 2957
rect 20713 2952 24042 2954
rect 20713 2896 20718 2952
rect 20774 2896 24042 2952
rect 20713 2894 24042 2896
rect 20713 2891 20779 2894
rect 6269 2816 7114 2818
rect 6269 2760 6274 2816
rect 6330 2760 7114 2816
rect 6269 2758 7114 2760
rect 23982 2818 24042 2894
rect 25840 2818 26000 2848
rect 23982 2758 26000 2818
rect 6269 2755 6335 2758
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 25840 2728 26000 2758
rect 21715 2687 22031 2688
rect 4889 2682 4955 2685
rect 8109 2682 8175 2685
rect 4889 2680 8175 2682
rect 4889 2624 4894 2680
rect 4950 2624 8114 2680
rect 8170 2624 8175 2680
rect 4889 2622 8175 2624
rect 4889 2619 4955 2622
rect 8109 2619 8175 2622
rect 12065 2682 12131 2685
rect 12566 2682 12572 2684
rect 12065 2680 12572 2682
rect 12065 2624 12070 2680
rect 12126 2624 12572 2680
rect 12065 2622 12572 2624
rect 12065 2619 12131 2622
rect 12566 2620 12572 2622
rect 12636 2620 12642 2684
rect 13813 2682 13879 2685
rect 14038 2682 14044 2684
rect 13813 2680 14044 2682
rect 13813 2624 13818 2680
rect 13874 2624 14044 2680
rect 13813 2622 14044 2624
rect 13813 2619 13879 2622
rect 14038 2620 14044 2622
rect 14108 2620 14114 2684
rect 16297 2682 16363 2685
rect 20529 2682 20595 2685
rect 16297 2680 20595 2682
rect 16297 2624 16302 2680
rect 16358 2624 20534 2680
rect 20590 2624 20595 2680
rect 16297 2622 20595 2624
rect 16297 2619 16363 2622
rect 20529 2619 20595 2622
rect 6177 2546 6243 2549
rect 8334 2546 8340 2548
rect 6177 2544 8340 2546
rect 6177 2488 6182 2544
rect 6238 2488 8340 2544
rect 6177 2486 8340 2488
rect 6177 2483 6243 2486
rect 8334 2484 8340 2486
rect 8404 2484 8410 2548
rect 20294 2484 20300 2548
rect 20364 2546 20370 2548
rect 21909 2546 21975 2549
rect 20364 2544 21975 2546
rect 20364 2488 21914 2544
rect 21970 2488 21975 2544
rect 20364 2486 21975 2488
rect 20364 2484 20370 2486
rect 21909 2483 21975 2486
rect 1853 2410 1919 2413
rect 13537 2410 13603 2413
rect 1853 2408 13603 2410
rect 1853 2352 1858 2408
rect 1914 2352 13542 2408
rect 13598 2352 13603 2408
rect 1853 2350 13603 2352
rect 1853 2347 1919 2350
rect 13537 2347 13603 2350
rect 14273 2410 14339 2413
rect 14406 2410 14412 2412
rect 14273 2408 14412 2410
rect 14273 2352 14278 2408
rect 14334 2352 14412 2408
rect 14273 2350 14412 2352
rect 14273 2347 14339 2350
rect 14406 2348 14412 2350
rect 14476 2348 14482 2412
rect 17677 2410 17743 2413
rect 22369 2410 22435 2413
rect 17677 2408 22435 2410
rect 17677 2352 17682 2408
rect 17738 2352 22374 2408
rect 22430 2352 22435 2408
rect 17677 2350 22435 2352
rect 17677 2347 17743 2350
rect 22369 2347 22435 2350
rect 24534 2350 25146 2410
rect 1158 2212 1164 2276
rect 1228 2274 1234 2276
rect 1228 2214 2790 2274
rect 1228 2212 1234 2214
rect 2730 2138 2790 2214
rect 3734 2212 3740 2276
rect 3804 2274 3810 2276
rect 3969 2274 4035 2277
rect 3804 2272 4035 2274
rect 3804 2216 3974 2272
rect 4030 2216 4035 2272
rect 3804 2214 4035 2216
rect 3804 2212 3810 2214
rect 3969 2211 4035 2214
rect 5809 2274 5875 2277
rect 7925 2276 7991 2277
rect 6494 2274 6500 2276
rect 5809 2272 6500 2274
rect 5809 2216 5814 2272
rect 5870 2216 6500 2272
rect 5809 2214 6500 2216
rect 5809 2211 5875 2214
rect 6494 2212 6500 2214
rect 6564 2212 6570 2276
rect 7925 2274 7972 2276
rect 7880 2272 7972 2274
rect 7880 2216 7930 2272
rect 7880 2214 7972 2216
rect 7925 2212 7972 2214
rect 8036 2212 8042 2276
rect 10317 2274 10383 2277
rect 10910 2274 10916 2276
rect 10317 2272 10916 2274
rect 10317 2216 10322 2272
rect 10378 2216 10916 2272
rect 10317 2214 10916 2216
rect 7925 2211 7991 2212
rect 10317 2211 10383 2214
rect 10910 2212 10916 2214
rect 10980 2212 10986 2276
rect 22093 2274 22159 2277
rect 24534 2274 24594 2350
rect 22093 2272 24594 2274
rect 22093 2216 22098 2272
rect 22154 2216 24594 2272
rect 22093 2214 24594 2216
rect 25086 2274 25146 2350
rect 25840 2274 26000 2304
rect 25086 2214 26000 2274
rect 22093 2211 22159 2214
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 25840 2184 26000 2214
rect 24682 2143 24998 2144
rect 4981 2138 5047 2141
rect 2730 2136 5047 2138
rect 2730 2080 4986 2136
rect 5042 2080 5047 2136
rect 2730 2078 5047 2080
rect 4981 2075 5047 2078
rect 8017 2002 8083 2005
rect 14181 2002 14247 2005
rect 8017 2000 14247 2002
rect 8017 1944 8022 2000
rect 8078 1944 14186 2000
rect 14242 1944 14247 2000
rect 8017 1942 14247 1944
rect 8017 1939 8083 1942
rect 14181 1939 14247 1942
rect 657 1866 723 1869
rect 13813 1866 13879 1869
rect 657 1864 13879 1866
rect 657 1808 662 1864
rect 718 1808 13818 1864
rect 13874 1808 13879 1864
rect 657 1806 13879 1808
rect 657 1803 723 1806
rect 13813 1803 13879 1806
rect 20713 1866 20779 1869
rect 20713 1864 24042 1866
rect 20713 1808 20718 1864
rect 20774 1808 24042 1864
rect 20713 1806 24042 1808
rect 20713 1803 20779 1806
rect 5073 1730 5139 1733
rect 8886 1730 8892 1732
rect 5073 1728 8892 1730
rect 5073 1672 5078 1728
rect 5134 1672 8892 1728
rect 5073 1670 8892 1672
rect 5073 1667 5139 1670
rect 8886 1668 8892 1670
rect 8956 1668 8962 1732
rect 23982 1730 24042 1806
rect 25840 1730 26000 1760
rect 23982 1670 26000 1730
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 25840 1640 26000 1670
rect 21715 1599 22031 1600
rect 841 1458 907 1461
rect 11513 1458 11579 1461
rect 841 1456 11579 1458
rect 841 1400 846 1456
rect 902 1400 11518 1456
rect 11574 1400 11579 1456
rect 841 1398 11579 1400
rect 841 1395 907 1398
rect 11513 1395 11579 1398
rect 1853 1324 1919 1325
rect 1853 1322 1900 1324
rect 1808 1320 1900 1322
rect 1808 1264 1858 1320
rect 1808 1262 1900 1264
rect 1853 1260 1900 1262
rect 1964 1260 1970 1324
rect 2497 1322 2563 1325
rect 2630 1322 2636 1324
rect 2497 1320 2636 1322
rect 2497 1264 2502 1320
rect 2558 1264 2636 1320
rect 2497 1262 2636 1264
rect 1853 1259 1919 1260
rect 2497 1259 2563 1262
rect 2630 1260 2636 1262
rect 2700 1260 2706 1324
rect 5022 1260 5028 1324
rect 5092 1322 5098 1324
rect 5533 1322 5599 1325
rect 9029 1324 9095 1325
rect 5092 1320 5599 1322
rect 5092 1264 5538 1320
rect 5594 1264 5599 1320
rect 5092 1262 5599 1264
rect 5092 1260 5098 1262
rect 5533 1259 5599 1262
rect 6126 1260 6132 1324
rect 6196 1260 6202 1324
rect 9029 1322 9076 1324
rect 8984 1320 9076 1322
rect 8984 1264 9034 1320
rect 8984 1262 9076 1264
rect 9029 1260 9076 1262
rect 9140 1260 9146 1324
rect 19057 1322 19123 1325
rect 19374 1322 19380 1324
rect 19057 1320 19380 1322
rect 19057 1264 19062 1320
rect 19118 1264 19380 1320
rect 19057 1262 19380 1264
rect 5073 1186 5139 1189
rect 6134 1186 6194 1260
rect 9029 1259 9095 1260
rect 19057 1259 19123 1262
rect 19374 1260 19380 1262
rect 19444 1260 19450 1324
rect 20478 1260 20484 1324
rect 20548 1322 20554 1324
rect 21633 1322 21699 1325
rect 20548 1320 21699 1322
rect 20548 1264 21638 1320
rect 21694 1264 21699 1320
rect 20548 1262 21699 1264
rect 20548 1260 20554 1262
rect 21633 1259 21699 1262
rect 5073 1184 6194 1186
rect 5073 1128 5078 1184
rect 5134 1128 6194 1184
rect 5073 1126 6194 1128
rect 21357 1186 21423 1189
rect 23238 1186 23244 1188
rect 21357 1184 23244 1186
rect 21357 1128 21362 1184
rect 21418 1128 23244 1184
rect 21357 1126 23244 1128
rect 5073 1123 5139 1126
rect 21357 1123 21423 1126
rect 23238 1124 23244 1126
rect 23308 1124 23314 1188
rect 25497 1186 25563 1189
rect 25840 1186 26000 1216
rect 25497 1184 26000 1186
rect 25497 1128 25502 1184
rect 25558 1128 26000 1184
rect 25497 1126 26000 1128
rect 25497 1123 25563 1126
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 25840 1096 26000 1126
rect 24682 1055 24998 1056
rect 7557 914 7623 917
rect 19926 914 19932 916
rect 7557 912 19932 914
rect 7557 856 7562 912
rect 7618 856 19932 912
rect 7557 854 19932 856
rect 7557 851 7623 854
rect 19926 852 19932 854
rect 19996 852 20002 916
rect 20713 642 20779 645
rect 25840 642 26000 672
rect 20713 640 26000 642
rect 20713 584 20718 640
rect 20774 584 26000 640
rect 20713 582 26000 584
rect 20713 579 20779 582
rect 25840 552 26000 582
<< via3 >>
rect 18460 44508 18524 44572
rect 6886 43548 6950 43552
rect 6886 43492 6890 43548
rect 6890 43492 6946 43548
rect 6946 43492 6950 43548
rect 6886 43488 6950 43492
rect 6966 43548 7030 43552
rect 6966 43492 6970 43548
rect 6970 43492 7026 43548
rect 7026 43492 7030 43548
rect 6966 43488 7030 43492
rect 7046 43548 7110 43552
rect 7046 43492 7050 43548
rect 7050 43492 7106 43548
rect 7106 43492 7110 43548
rect 7046 43488 7110 43492
rect 7126 43548 7190 43552
rect 7126 43492 7130 43548
rect 7130 43492 7186 43548
rect 7186 43492 7190 43548
rect 7126 43488 7190 43492
rect 12820 43548 12884 43552
rect 12820 43492 12824 43548
rect 12824 43492 12880 43548
rect 12880 43492 12884 43548
rect 12820 43488 12884 43492
rect 12900 43548 12964 43552
rect 12900 43492 12904 43548
rect 12904 43492 12960 43548
rect 12960 43492 12964 43548
rect 12900 43488 12964 43492
rect 12980 43548 13044 43552
rect 12980 43492 12984 43548
rect 12984 43492 13040 43548
rect 13040 43492 13044 43548
rect 12980 43488 13044 43492
rect 13060 43548 13124 43552
rect 13060 43492 13064 43548
rect 13064 43492 13120 43548
rect 13120 43492 13124 43548
rect 13060 43488 13124 43492
rect 18754 43548 18818 43552
rect 18754 43492 18758 43548
rect 18758 43492 18814 43548
rect 18814 43492 18818 43548
rect 18754 43488 18818 43492
rect 18834 43548 18898 43552
rect 18834 43492 18838 43548
rect 18838 43492 18894 43548
rect 18894 43492 18898 43548
rect 18834 43488 18898 43492
rect 18914 43548 18978 43552
rect 18914 43492 18918 43548
rect 18918 43492 18974 43548
rect 18974 43492 18978 43548
rect 18914 43488 18978 43492
rect 18994 43548 19058 43552
rect 18994 43492 18998 43548
rect 18998 43492 19054 43548
rect 19054 43492 19058 43548
rect 18994 43488 19058 43492
rect 24688 43548 24752 43552
rect 24688 43492 24692 43548
rect 24692 43492 24748 43548
rect 24748 43492 24752 43548
rect 24688 43488 24752 43492
rect 24768 43548 24832 43552
rect 24768 43492 24772 43548
rect 24772 43492 24828 43548
rect 24828 43492 24832 43548
rect 24768 43488 24832 43492
rect 24848 43548 24912 43552
rect 24848 43492 24852 43548
rect 24852 43492 24908 43548
rect 24908 43492 24912 43548
rect 24848 43488 24912 43492
rect 24928 43548 24992 43552
rect 24928 43492 24932 43548
rect 24932 43492 24988 43548
rect 24988 43492 24992 43548
rect 24928 43488 24992 43492
rect 15516 43284 15580 43348
rect 21588 43148 21652 43212
rect 14596 43012 14660 43076
rect 3919 43004 3983 43008
rect 3919 42948 3923 43004
rect 3923 42948 3979 43004
rect 3979 42948 3983 43004
rect 3919 42944 3983 42948
rect 3999 43004 4063 43008
rect 3999 42948 4003 43004
rect 4003 42948 4059 43004
rect 4059 42948 4063 43004
rect 3999 42944 4063 42948
rect 4079 43004 4143 43008
rect 4079 42948 4083 43004
rect 4083 42948 4139 43004
rect 4139 42948 4143 43004
rect 4079 42944 4143 42948
rect 4159 43004 4223 43008
rect 4159 42948 4163 43004
rect 4163 42948 4219 43004
rect 4219 42948 4223 43004
rect 4159 42944 4223 42948
rect 9853 43004 9917 43008
rect 9853 42948 9857 43004
rect 9857 42948 9913 43004
rect 9913 42948 9917 43004
rect 9853 42944 9917 42948
rect 9933 43004 9997 43008
rect 9933 42948 9937 43004
rect 9937 42948 9993 43004
rect 9993 42948 9997 43004
rect 9933 42944 9997 42948
rect 10013 43004 10077 43008
rect 10013 42948 10017 43004
rect 10017 42948 10073 43004
rect 10073 42948 10077 43004
rect 10013 42944 10077 42948
rect 10093 43004 10157 43008
rect 10093 42948 10097 43004
rect 10097 42948 10153 43004
rect 10153 42948 10157 43004
rect 10093 42944 10157 42948
rect 15787 43004 15851 43008
rect 15787 42948 15791 43004
rect 15791 42948 15847 43004
rect 15847 42948 15851 43004
rect 15787 42944 15851 42948
rect 15867 43004 15931 43008
rect 15867 42948 15871 43004
rect 15871 42948 15927 43004
rect 15927 42948 15931 43004
rect 15867 42944 15931 42948
rect 15947 43004 16011 43008
rect 15947 42948 15951 43004
rect 15951 42948 16007 43004
rect 16007 42948 16011 43004
rect 15947 42944 16011 42948
rect 16027 43004 16091 43008
rect 16027 42948 16031 43004
rect 16031 42948 16087 43004
rect 16087 42948 16091 43004
rect 16027 42944 16091 42948
rect 10364 42876 10428 42940
rect 13308 42876 13372 42940
rect 14964 42936 15028 42940
rect 14964 42880 14978 42936
rect 14978 42880 15028 42936
rect 14964 42876 15028 42880
rect 6886 42460 6950 42464
rect 6886 42404 6890 42460
rect 6890 42404 6946 42460
rect 6946 42404 6950 42460
rect 6886 42400 6950 42404
rect 6966 42460 7030 42464
rect 6966 42404 6970 42460
rect 6970 42404 7026 42460
rect 7026 42404 7030 42460
rect 6966 42400 7030 42404
rect 7046 42460 7110 42464
rect 7046 42404 7050 42460
rect 7050 42404 7106 42460
rect 7106 42404 7110 42460
rect 7046 42400 7110 42404
rect 7126 42460 7190 42464
rect 7126 42404 7130 42460
rect 7130 42404 7186 42460
rect 7186 42404 7190 42460
rect 7126 42400 7190 42404
rect 12820 42460 12884 42464
rect 12820 42404 12824 42460
rect 12824 42404 12880 42460
rect 12880 42404 12884 42460
rect 12820 42400 12884 42404
rect 12900 42460 12964 42464
rect 12900 42404 12904 42460
rect 12904 42404 12960 42460
rect 12960 42404 12964 42460
rect 12900 42400 12964 42404
rect 12980 42460 13044 42464
rect 12980 42404 12984 42460
rect 12984 42404 13040 42460
rect 13040 42404 13044 42460
rect 12980 42400 13044 42404
rect 13060 42460 13124 42464
rect 13060 42404 13064 42460
rect 13064 42404 13120 42460
rect 13120 42404 13124 42460
rect 13060 42400 13124 42404
rect 18754 42460 18818 42464
rect 18754 42404 18758 42460
rect 18758 42404 18814 42460
rect 18814 42404 18818 42460
rect 18754 42400 18818 42404
rect 18834 42460 18898 42464
rect 18834 42404 18838 42460
rect 18838 42404 18894 42460
rect 18894 42404 18898 42460
rect 18834 42400 18898 42404
rect 18914 42460 18978 42464
rect 18914 42404 18918 42460
rect 18918 42404 18974 42460
rect 18974 42404 18978 42460
rect 18914 42400 18978 42404
rect 18994 42460 19058 42464
rect 18994 42404 18998 42460
rect 18998 42404 19054 42460
rect 19054 42404 19058 42460
rect 18994 42400 19058 42404
rect 21721 43004 21785 43008
rect 21721 42948 21725 43004
rect 21725 42948 21781 43004
rect 21781 42948 21785 43004
rect 21721 42944 21785 42948
rect 21801 43004 21865 43008
rect 21801 42948 21805 43004
rect 21805 42948 21861 43004
rect 21861 42948 21865 43004
rect 21801 42944 21865 42948
rect 21881 43004 21945 43008
rect 21881 42948 21885 43004
rect 21885 42948 21941 43004
rect 21941 42948 21945 43004
rect 21881 42944 21945 42948
rect 21961 43004 22025 43008
rect 21961 42948 21965 43004
rect 21965 42948 22021 43004
rect 22021 42948 22025 43004
rect 21961 42944 22025 42948
rect 24688 42460 24752 42464
rect 24688 42404 24692 42460
rect 24692 42404 24748 42460
rect 24748 42404 24752 42460
rect 24688 42400 24752 42404
rect 24768 42460 24832 42464
rect 24768 42404 24772 42460
rect 24772 42404 24828 42460
rect 24828 42404 24832 42460
rect 24768 42400 24832 42404
rect 24848 42460 24912 42464
rect 24848 42404 24852 42460
rect 24852 42404 24908 42460
rect 24908 42404 24912 42460
rect 24848 42400 24912 42404
rect 24928 42460 24992 42464
rect 24928 42404 24932 42460
rect 24932 42404 24988 42460
rect 24988 42404 24992 42460
rect 24928 42400 24992 42404
rect 1164 42196 1228 42260
rect 11652 42060 11716 42124
rect 18460 42196 18524 42260
rect 20668 42060 20732 42124
rect 11836 41984 11900 41988
rect 11836 41928 11850 41984
rect 11850 41928 11900 41984
rect 11836 41924 11900 41928
rect 3919 41916 3983 41920
rect 3919 41860 3923 41916
rect 3923 41860 3979 41916
rect 3979 41860 3983 41916
rect 3919 41856 3983 41860
rect 3999 41916 4063 41920
rect 3999 41860 4003 41916
rect 4003 41860 4059 41916
rect 4059 41860 4063 41916
rect 3999 41856 4063 41860
rect 4079 41916 4143 41920
rect 4079 41860 4083 41916
rect 4083 41860 4139 41916
rect 4139 41860 4143 41916
rect 4079 41856 4143 41860
rect 4159 41916 4223 41920
rect 4159 41860 4163 41916
rect 4163 41860 4219 41916
rect 4219 41860 4223 41916
rect 4159 41856 4223 41860
rect 9853 41916 9917 41920
rect 9853 41860 9857 41916
rect 9857 41860 9913 41916
rect 9913 41860 9917 41916
rect 9853 41856 9917 41860
rect 9933 41916 9997 41920
rect 9933 41860 9937 41916
rect 9937 41860 9993 41916
rect 9993 41860 9997 41916
rect 9933 41856 9997 41860
rect 10013 41916 10077 41920
rect 10013 41860 10017 41916
rect 10017 41860 10073 41916
rect 10073 41860 10077 41916
rect 10013 41856 10077 41860
rect 10093 41916 10157 41920
rect 10093 41860 10097 41916
rect 10097 41860 10153 41916
rect 10153 41860 10157 41916
rect 10093 41856 10157 41860
rect 15787 41916 15851 41920
rect 15787 41860 15791 41916
rect 15791 41860 15847 41916
rect 15847 41860 15851 41916
rect 15787 41856 15851 41860
rect 15867 41916 15931 41920
rect 15867 41860 15871 41916
rect 15871 41860 15927 41916
rect 15927 41860 15931 41916
rect 15867 41856 15931 41860
rect 15947 41916 16011 41920
rect 15947 41860 15951 41916
rect 15951 41860 16007 41916
rect 16007 41860 16011 41916
rect 15947 41856 16011 41860
rect 16027 41916 16091 41920
rect 16027 41860 16031 41916
rect 16031 41860 16087 41916
rect 16087 41860 16091 41916
rect 16027 41856 16091 41860
rect 21721 41916 21785 41920
rect 21721 41860 21725 41916
rect 21725 41860 21781 41916
rect 21781 41860 21785 41916
rect 21721 41856 21785 41860
rect 21801 41916 21865 41920
rect 21801 41860 21805 41916
rect 21805 41860 21861 41916
rect 21861 41860 21865 41916
rect 21801 41856 21865 41860
rect 21881 41916 21945 41920
rect 21881 41860 21885 41916
rect 21885 41860 21941 41916
rect 21941 41860 21945 41916
rect 21881 41856 21945 41860
rect 21961 41916 22025 41920
rect 21961 41860 21965 41916
rect 21965 41860 22021 41916
rect 22021 41860 22025 41916
rect 21961 41856 22025 41860
rect 6316 41848 6380 41852
rect 6316 41792 6330 41848
rect 6330 41792 6380 41848
rect 6316 41788 6380 41792
rect 7604 41788 7668 41852
rect 8156 41848 8220 41852
rect 8156 41792 8206 41848
rect 8206 41792 8220 41848
rect 8156 41788 8220 41792
rect 16988 41712 17052 41716
rect 16988 41656 17002 41712
rect 17002 41656 17052 41712
rect 16988 41652 17052 41656
rect 17724 41712 17788 41716
rect 17724 41656 17738 41712
rect 17738 41656 17788 41712
rect 17724 41652 17788 41656
rect 18276 41712 18340 41716
rect 18276 41656 18326 41712
rect 18326 41656 18340 41712
rect 18276 41652 18340 41656
rect 19564 41712 19628 41716
rect 19564 41656 19578 41712
rect 19578 41656 19628 41712
rect 19564 41652 19628 41656
rect 980 41380 1044 41444
rect 18460 41440 18524 41444
rect 18460 41384 18474 41440
rect 18474 41384 18524 41440
rect 18460 41380 18524 41384
rect 6886 41372 6950 41376
rect 6886 41316 6890 41372
rect 6890 41316 6946 41372
rect 6946 41316 6950 41372
rect 6886 41312 6950 41316
rect 6966 41372 7030 41376
rect 6966 41316 6970 41372
rect 6970 41316 7026 41372
rect 7026 41316 7030 41372
rect 6966 41312 7030 41316
rect 7046 41372 7110 41376
rect 7046 41316 7050 41372
rect 7050 41316 7106 41372
rect 7106 41316 7110 41372
rect 7046 41312 7110 41316
rect 7126 41372 7190 41376
rect 7126 41316 7130 41372
rect 7130 41316 7186 41372
rect 7186 41316 7190 41372
rect 7126 41312 7190 41316
rect 12820 41372 12884 41376
rect 12820 41316 12824 41372
rect 12824 41316 12880 41372
rect 12880 41316 12884 41372
rect 12820 41312 12884 41316
rect 12900 41372 12964 41376
rect 12900 41316 12904 41372
rect 12904 41316 12960 41372
rect 12960 41316 12964 41372
rect 12900 41312 12964 41316
rect 12980 41372 13044 41376
rect 12980 41316 12984 41372
rect 12984 41316 13040 41372
rect 13040 41316 13044 41372
rect 12980 41312 13044 41316
rect 13060 41372 13124 41376
rect 13060 41316 13064 41372
rect 13064 41316 13120 41372
rect 13120 41316 13124 41372
rect 13060 41312 13124 41316
rect 18754 41372 18818 41376
rect 18754 41316 18758 41372
rect 18758 41316 18814 41372
rect 18814 41316 18818 41372
rect 18754 41312 18818 41316
rect 18834 41372 18898 41376
rect 18834 41316 18838 41372
rect 18838 41316 18894 41372
rect 18894 41316 18898 41372
rect 18834 41312 18898 41316
rect 18914 41372 18978 41376
rect 18914 41316 18918 41372
rect 18918 41316 18974 41372
rect 18974 41316 18978 41372
rect 18914 41312 18978 41316
rect 18994 41372 19058 41376
rect 18994 41316 18998 41372
rect 18998 41316 19054 41372
rect 19054 41316 19058 41372
rect 18994 41312 19058 41316
rect 24688 41372 24752 41376
rect 24688 41316 24692 41372
rect 24692 41316 24748 41372
rect 24748 41316 24752 41372
rect 24688 41312 24752 41316
rect 24768 41372 24832 41376
rect 24768 41316 24772 41372
rect 24772 41316 24828 41372
rect 24828 41316 24832 41372
rect 24768 41312 24832 41316
rect 24848 41372 24912 41376
rect 24848 41316 24852 41372
rect 24852 41316 24908 41372
rect 24908 41316 24912 41372
rect 24848 41312 24912 41316
rect 24928 41372 24992 41376
rect 24928 41316 24932 41372
rect 24932 41316 24988 41372
rect 24988 41316 24992 41372
rect 24928 41312 24992 41316
rect 21588 40972 21652 41036
rect 3919 40828 3983 40832
rect 3919 40772 3923 40828
rect 3923 40772 3979 40828
rect 3979 40772 3983 40828
rect 3919 40768 3983 40772
rect 3999 40828 4063 40832
rect 3999 40772 4003 40828
rect 4003 40772 4059 40828
rect 4059 40772 4063 40828
rect 3999 40768 4063 40772
rect 4079 40828 4143 40832
rect 4079 40772 4083 40828
rect 4083 40772 4139 40828
rect 4139 40772 4143 40828
rect 4079 40768 4143 40772
rect 4159 40828 4223 40832
rect 4159 40772 4163 40828
rect 4163 40772 4219 40828
rect 4219 40772 4223 40828
rect 4159 40768 4223 40772
rect 9853 40828 9917 40832
rect 9853 40772 9857 40828
rect 9857 40772 9913 40828
rect 9913 40772 9917 40828
rect 9853 40768 9917 40772
rect 9933 40828 9997 40832
rect 9933 40772 9937 40828
rect 9937 40772 9993 40828
rect 9993 40772 9997 40828
rect 9933 40768 9997 40772
rect 10013 40828 10077 40832
rect 10013 40772 10017 40828
rect 10017 40772 10073 40828
rect 10073 40772 10077 40828
rect 10013 40768 10077 40772
rect 10093 40828 10157 40832
rect 10093 40772 10097 40828
rect 10097 40772 10153 40828
rect 10153 40772 10157 40828
rect 10093 40768 10157 40772
rect 15787 40828 15851 40832
rect 15787 40772 15791 40828
rect 15791 40772 15847 40828
rect 15847 40772 15851 40828
rect 15787 40768 15851 40772
rect 15867 40828 15931 40832
rect 15867 40772 15871 40828
rect 15871 40772 15927 40828
rect 15927 40772 15931 40828
rect 15867 40768 15931 40772
rect 15947 40828 16011 40832
rect 15947 40772 15951 40828
rect 15951 40772 16007 40828
rect 16007 40772 16011 40828
rect 15947 40768 16011 40772
rect 16027 40828 16091 40832
rect 16027 40772 16031 40828
rect 16031 40772 16087 40828
rect 16087 40772 16091 40828
rect 16027 40768 16091 40772
rect 21721 40828 21785 40832
rect 21721 40772 21725 40828
rect 21725 40772 21781 40828
rect 21781 40772 21785 40828
rect 21721 40768 21785 40772
rect 21801 40828 21865 40832
rect 21801 40772 21805 40828
rect 21805 40772 21861 40828
rect 21861 40772 21865 40828
rect 21801 40768 21865 40772
rect 21881 40828 21945 40832
rect 21881 40772 21885 40828
rect 21885 40772 21941 40828
rect 21941 40772 21945 40828
rect 21881 40768 21945 40772
rect 21961 40828 22025 40832
rect 21961 40772 21965 40828
rect 21965 40772 22021 40828
rect 22021 40772 22025 40828
rect 21961 40768 22025 40772
rect 612 40564 676 40628
rect 796 40292 860 40356
rect 6886 40284 6950 40288
rect 6886 40228 6890 40284
rect 6890 40228 6946 40284
rect 6946 40228 6950 40284
rect 6886 40224 6950 40228
rect 6966 40284 7030 40288
rect 6966 40228 6970 40284
rect 6970 40228 7026 40284
rect 7026 40228 7030 40284
rect 6966 40224 7030 40228
rect 7046 40284 7110 40288
rect 7046 40228 7050 40284
rect 7050 40228 7106 40284
rect 7106 40228 7110 40284
rect 7046 40224 7110 40228
rect 7126 40284 7190 40288
rect 7126 40228 7130 40284
rect 7130 40228 7186 40284
rect 7186 40228 7190 40284
rect 7126 40224 7190 40228
rect 12820 40284 12884 40288
rect 12820 40228 12824 40284
rect 12824 40228 12880 40284
rect 12880 40228 12884 40284
rect 12820 40224 12884 40228
rect 12900 40284 12964 40288
rect 12900 40228 12904 40284
rect 12904 40228 12960 40284
rect 12960 40228 12964 40284
rect 12900 40224 12964 40228
rect 12980 40284 13044 40288
rect 12980 40228 12984 40284
rect 12984 40228 13040 40284
rect 13040 40228 13044 40284
rect 12980 40224 13044 40228
rect 13060 40284 13124 40288
rect 13060 40228 13064 40284
rect 13064 40228 13120 40284
rect 13120 40228 13124 40284
rect 13060 40224 13124 40228
rect 18754 40284 18818 40288
rect 18754 40228 18758 40284
rect 18758 40228 18814 40284
rect 18814 40228 18818 40284
rect 18754 40224 18818 40228
rect 18834 40284 18898 40288
rect 18834 40228 18838 40284
rect 18838 40228 18894 40284
rect 18894 40228 18898 40284
rect 18834 40224 18898 40228
rect 18914 40284 18978 40288
rect 18914 40228 18918 40284
rect 18918 40228 18974 40284
rect 18974 40228 18978 40284
rect 18914 40224 18978 40228
rect 18994 40284 19058 40288
rect 18994 40228 18998 40284
rect 18998 40228 19054 40284
rect 19054 40228 19058 40284
rect 18994 40224 19058 40228
rect 24688 40284 24752 40288
rect 24688 40228 24692 40284
rect 24692 40228 24748 40284
rect 24748 40228 24752 40284
rect 24688 40224 24752 40228
rect 24768 40284 24832 40288
rect 24768 40228 24772 40284
rect 24772 40228 24828 40284
rect 24828 40228 24832 40284
rect 24768 40224 24832 40228
rect 24848 40284 24912 40288
rect 24848 40228 24852 40284
rect 24852 40228 24908 40284
rect 24908 40228 24912 40284
rect 24848 40224 24912 40228
rect 24928 40284 24992 40288
rect 24928 40228 24932 40284
rect 24932 40228 24988 40284
rect 24988 40228 24992 40284
rect 24928 40224 24992 40228
rect 2636 40156 2700 40220
rect 3372 40020 3436 40084
rect 9628 40020 9692 40084
rect 3919 39740 3983 39744
rect 3919 39684 3923 39740
rect 3923 39684 3979 39740
rect 3979 39684 3983 39740
rect 3919 39680 3983 39684
rect 3999 39740 4063 39744
rect 3999 39684 4003 39740
rect 4003 39684 4059 39740
rect 4059 39684 4063 39740
rect 3999 39680 4063 39684
rect 4079 39740 4143 39744
rect 4079 39684 4083 39740
rect 4083 39684 4139 39740
rect 4139 39684 4143 39740
rect 4079 39680 4143 39684
rect 4159 39740 4223 39744
rect 4159 39684 4163 39740
rect 4163 39684 4219 39740
rect 4219 39684 4223 39740
rect 4159 39680 4223 39684
rect 9853 39740 9917 39744
rect 9853 39684 9857 39740
rect 9857 39684 9913 39740
rect 9913 39684 9917 39740
rect 9853 39680 9917 39684
rect 9933 39740 9997 39744
rect 9933 39684 9937 39740
rect 9937 39684 9993 39740
rect 9993 39684 9997 39740
rect 9933 39680 9997 39684
rect 10013 39740 10077 39744
rect 10013 39684 10017 39740
rect 10017 39684 10073 39740
rect 10073 39684 10077 39740
rect 10013 39680 10077 39684
rect 10093 39740 10157 39744
rect 10093 39684 10097 39740
rect 10097 39684 10153 39740
rect 10153 39684 10157 39740
rect 10093 39680 10157 39684
rect 15787 39740 15851 39744
rect 15787 39684 15791 39740
rect 15791 39684 15847 39740
rect 15847 39684 15851 39740
rect 15787 39680 15851 39684
rect 15867 39740 15931 39744
rect 15867 39684 15871 39740
rect 15871 39684 15927 39740
rect 15927 39684 15931 39740
rect 15867 39680 15931 39684
rect 15947 39740 16011 39744
rect 15947 39684 15951 39740
rect 15951 39684 16007 39740
rect 16007 39684 16011 39740
rect 15947 39680 16011 39684
rect 16027 39740 16091 39744
rect 16027 39684 16031 39740
rect 16031 39684 16087 39740
rect 16087 39684 16091 39740
rect 16027 39680 16091 39684
rect 21721 39740 21785 39744
rect 21721 39684 21725 39740
rect 21725 39684 21781 39740
rect 21781 39684 21785 39740
rect 21721 39680 21785 39684
rect 21801 39740 21865 39744
rect 21801 39684 21805 39740
rect 21805 39684 21861 39740
rect 21861 39684 21865 39740
rect 21801 39680 21865 39684
rect 21881 39740 21945 39744
rect 21881 39684 21885 39740
rect 21885 39684 21941 39740
rect 21941 39684 21945 39740
rect 21881 39680 21945 39684
rect 21961 39740 22025 39744
rect 21961 39684 21965 39740
rect 21965 39684 22021 39740
rect 22021 39684 22025 39740
rect 21961 39680 22025 39684
rect 2268 39672 2332 39676
rect 2268 39616 2282 39672
rect 2282 39616 2332 39672
rect 2268 39612 2332 39616
rect 16436 39476 16500 39540
rect 12572 39340 12636 39404
rect 6886 39196 6950 39200
rect 6886 39140 6890 39196
rect 6890 39140 6946 39196
rect 6946 39140 6950 39196
rect 6886 39136 6950 39140
rect 6966 39196 7030 39200
rect 6966 39140 6970 39196
rect 6970 39140 7026 39196
rect 7026 39140 7030 39196
rect 6966 39136 7030 39140
rect 7046 39196 7110 39200
rect 7046 39140 7050 39196
rect 7050 39140 7106 39196
rect 7106 39140 7110 39196
rect 7046 39136 7110 39140
rect 7126 39196 7190 39200
rect 7126 39140 7130 39196
rect 7130 39140 7186 39196
rect 7186 39140 7190 39196
rect 7126 39136 7190 39140
rect 12820 39196 12884 39200
rect 12820 39140 12824 39196
rect 12824 39140 12880 39196
rect 12880 39140 12884 39196
rect 12820 39136 12884 39140
rect 12900 39196 12964 39200
rect 12900 39140 12904 39196
rect 12904 39140 12960 39196
rect 12960 39140 12964 39196
rect 12900 39136 12964 39140
rect 12980 39196 13044 39200
rect 12980 39140 12984 39196
rect 12984 39140 13040 39196
rect 13040 39140 13044 39196
rect 12980 39136 13044 39140
rect 13060 39196 13124 39200
rect 13060 39140 13064 39196
rect 13064 39140 13120 39196
rect 13120 39140 13124 39196
rect 13060 39136 13124 39140
rect 18754 39196 18818 39200
rect 18754 39140 18758 39196
rect 18758 39140 18814 39196
rect 18814 39140 18818 39196
rect 18754 39136 18818 39140
rect 18834 39196 18898 39200
rect 18834 39140 18838 39196
rect 18838 39140 18894 39196
rect 18894 39140 18898 39196
rect 18834 39136 18898 39140
rect 18914 39196 18978 39200
rect 18914 39140 18918 39196
rect 18918 39140 18974 39196
rect 18974 39140 18978 39196
rect 18914 39136 18978 39140
rect 18994 39196 19058 39200
rect 18994 39140 18998 39196
rect 18998 39140 19054 39196
rect 19054 39140 19058 39196
rect 18994 39136 19058 39140
rect 24688 39196 24752 39200
rect 24688 39140 24692 39196
rect 24692 39140 24748 39196
rect 24748 39140 24752 39196
rect 24688 39136 24752 39140
rect 24768 39196 24832 39200
rect 24768 39140 24772 39196
rect 24772 39140 24828 39196
rect 24828 39140 24832 39196
rect 24768 39136 24832 39140
rect 24848 39196 24912 39200
rect 24848 39140 24852 39196
rect 24852 39140 24908 39196
rect 24908 39140 24912 39196
rect 24848 39136 24912 39140
rect 24928 39196 24992 39200
rect 24928 39140 24932 39196
rect 24932 39140 24988 39196
rect 24988 39140 24992 39196
rect 24928 39136 24992 39140
rect 4292 38856 4356 38860
rect 4292 38800 4342 38856
rect 4342 38800 4356 38856
rect 4292 38796 4356 38800
rect 19748 38796 19812 38860
rect 20116 38660 20180 38724
rect 3919 38652 3983 38656
rect 3919 38596 3923 38652
rect 3923 38596 3979 38652
rect 3979 38596 3983 38652
rect 3919 38592 3983 38596
rect 3999 38652 4063 38656
rect 3999 38596 4003 38652
rect 4003 38596 4059 38652
rect 4059 38596 4063 38652
rect 3999 38592 4063 38596
rect 4079 38652 4143 38656
rect 4079 38596 4083 38652
rect 4083 38596 4139 38652
rect 4139 38596 4143 38652
rect 4079 38592 4143 38596
rect 4159 38652 4223 38656
rect 4159 38596 4163 38652
rect 4163 38596 4219 38652
rect 4219 38596 4223 38652
rect 4159 38592 4223 38596
rect 9853 38652 9917 38656
rect 9853 38596 9857 38652
rect 9857 38596 9913 38652
rect 9913 38596 9917 38652
rect 9853 38592 9917 38596
rect 9933 38652 9997 38656
rect 9933 38596 9937 38652
rect 9937 38596 9993 38652
rect 9993 38596 9997 38652
rect 9933 38592 9997 38596
rect 10013 38652 10077 38656
rect 10013 38596 10017 38652
rect 10017 38596 10073 38652
rect 10073 38596 10077 38652
rect 10013 38592 10077 38596
rect 10093 38652 10157 38656
rect 10093 38596 10097 38652
rect 10097 38596 10153 38652
rect 10153 38596 10157 38652
rect 10093 38592 10157 38596
rect 15787 38652 15851 38656
rect 15787 38596 15791 38652
rect 15791 38596 15847 38652
rect 15847 38596 15851 38652
rect 15787 38592 15851 38596
rect 15867 38652 15931 38656
rect 15867 38596 15871 38652
rect 15871 38596 15927 38652
rect 15927 38596 15931 38652
rect 15867 38592 15931 38596
rect 15947 38652 16011 38656
rect 15947 38596 15951 38652
rect 15951 38596 16007 38652
rect 16007 38596 16011 38652
rect 15947 38592 16011 38596
rect 16027 38652 16091 38656
rect 16027 38596 16031 38652
rect 16031 38596 16087 38652
rect 16087 38596 16091 38652
rect 16027 38592 16091 38596
rect 21721 38652 21785 38656
rect 21721 38596 21725 38652
rect 21725 38596 21781 38652
rect 21781 38596 21785 38652
rect 21721 38592 21785 38596
rect 21801 38652 21865 38656
rect 21801 38596 21805 38652
rect 21805 38596 21861 38652
rect 21861 38596 21865 38652
rect 21801 38592 21865 38596
rect 21881 38652 21945 38656
rect 21881 38596 21885 38652
rect 21885 38596 21941 38652
rect 21941 38596 21945 38652
rect 21881 38592 21945 38596
rect 21961 38652 22025 38656
rect 21961 38596 21965 38652
rect 21965 38596 22021 38652
rect 22021 38596 22025 38652
rect 21961 38592 22025 38596
rect 2084 38524 2148 38588
rect 13860 38252 13924 38316
rect 6886 38108 6950 38112
rect 6886 38052 6890 38108
rect 6890 38052 6946 38108
rect 6946 38052 6950 38108
rect 6886 38048 6950 38052
rect 6966 38108 7030 38112
rect 6966 38052 6970 38108
rect 6970 38052 7026 38108
rect 7026 38052 7030 38108
rect 6966 38048 7030 38052
rect 7046 38108 7110 38112
rect 7046 38052 7050 38108
rect 7050 38052 7106 38108
rect 7106 38052 7110 38108
rect 7046 38048 7110 38052
rect 7126 38108 7190 38112
rect 7126 38052 7130 38108
rect 7130 38052 7186 38108
rect 7186 38052 7190 38108
rect 7126 38048 7190 38052
rect 12820 38108 12884 38112
rect 12820 38052 12824 38108
rect 12824 38052 12880 38108
rect 12880 38052 12884 38108
rect 12820 38048 12884 38052
rect 12900 38108 12964 38112
rect 12900 38052 12904 38108
rect 12904 38052 12960 38108
rect 12960 38052 12964 38108
rect 12900 38048 12964 38052
rect 12980 38108 13044 38112
rect 12980 38052 12984 38108
rect 12984 38052 13040 38108
rect 13040 38052 13044 38108
rect 12980 38048 13044 38052
rect 13060 38108 13124 38112
rect 13060 38052 13064 38108
rect 13064 38052 13120 38108
rect 13120 38052 13124 38108
rect 13060 38048 13124 38052
rect 18754 38108 18818 38112
rect 18754 38052 18758 38108
rect 18758 38052 18814 38108
rect 18814 38052 18818 38108
rect 18754 38048 18818 38052
rect 18834 38108 18898 38112
rect 18834 38052 18838 38108
rect 18838 38052 18894 38108
rect 18894 38052 18898 38108
rect 18834 38048 18898 38052
rect 18914 38108 18978 38112
rect 18914 38052 18918 38108
rect 18918 38052 18974 38108
rect 18974 38052 18978 38108
rect 18914 38048 18978 38052
rect 18994 38108 19058 38112
rect 18994 38052 18998 38108
rect 18998 38052 19054 38108
rect 19054 38052 19058 38108
rect 18994 38048 19058 38052
rect 24688 38108 24752 38112
rect 24688 38052 24692 38108
rect 24692 38052 24748 38108
rect 24748 38052 24752 38108
rect 24688 38048 24752 38052
rect 24768 38108 24832 38112
rect 24768 38052 24772 38108
rect 24772 38052 24828 38108
rect 24828 38052 24832 38108
rect 24768 38048 24832 38052
rect 24848 38108 24912 38112
rect 24848 38052 24852 38108
rect 24852 38052 24908 38108
rect 24908 38052 24912 38108
rect 24848 38048 24912 38052
rect 24928 38108 24992 38112
rect 24928 38052 24932 38108
rect 24932 38052 24988 38108
rect 24988 38052 24992 38108
rect 24928 38048 24992 38052
rect 3919 37564 3983 37568
rect 3919 37508 3923 37564
rect 3923 37508 3979 37564
rect 3979 37508 3983 37564
rect 3919 37504 3983 37508
rect 3999 37564 4063 37568
rect 3999 37508 4003 37564
rect 4003 37508 4059 37564
rect 4059 37508 4063 37564
rect 3999 37504 4063 37508
rect 4079 37564 4143 37568
rect 4079 37508 4083 37564
rect 4083 37508 4139 37564
rect 4139 37508 4143 37564
rect 4079 37504 4143 37508
rect 4159 37564 4223 37568
rect 4159 37508 4163 37564
rect 4163 37508 4219 37564
rect 4219 37508 4223 37564
rect 4159 37504 4223 37508
rect 9853 37564 9917 37568
rect 9853 37508 9857 37564
rect 9857 37508 9913 37564
rect 9913 37508 9917 37564
rect 9853 37504 9917 37508
rect 9933 37564 9997 37568
rect 9933 37508 9937 37564
rect 9937 37508 9993 37564
rect 9993 37508 9997 37564
rect 9933 37504 9997 37508
rect 10013 37564 10077 37568
rect 10013 37508 10017 37564
rect 10017 37508 10073 37564
rect 10073 37508 10077 37564
rect 10013 37504 10077 37508
rect 10093 37564 10157 37568
rect 10093 37508 10097 37564
rect 10097 37508 10153 37564
rect 10153 37508 10157 37564
rect 10093 37504 10157 37508
rect 15787 37564 15851 37568
rect 15787 37508 15791 37564
rect 15791 37508 15847 37564
rect 15847 37508 15851 37564
rect 15787 37504 15851 37508
rect 15867 37564 15931 37568
rect 15867 37508 15871 37564
rect 15871 37508 15927 37564
rect 15927 37508 15931 37564
rect 15867 37504 15931 37508
rect 15947 37564 16011 37568
rect 15947 37508 15951 37564
rect 15951 37508 16007 37564
rect 16007 37508 16011 37564
rect 15947 37504 16011 37508
rect 16027 37564 16091 37568
rect 16027 37508 16031 37564
rect 16031 37508 16087 37564
rect 16087 37508 16091 37564
rect 16027 37504 16091 37508
rect 21721 37564 21785 37568
rect 21721 37508 21725 37564
rect 21725 37508 21781 37564
rect 21781 37508 21785 37564
rect 21721 37504 21785 37508
rect 21801 37564 21865 37568
rect 21801 37508 21805 37564
rect 21805 37508 21861 37564
rect 21861 37508 21865 37564
rect 21801 37504 21865 37508
rect 21881 37564 21945 37568
rect 21881 37508 21885 37564
rect 21885 37508 21941 37564
rect 21941 37508 21945 37564
rect 21881 37504 21945 37508
rect 21961 37564 22025 37568
rect 21961 37508 21965 37564
rect 21965 37508 22021 37564
rect 22021 37508 22025 37564
rect 21961 37504 22025 37508
rect 3188 37436 3252 37500
rect 5948 37300 6012 37364
rect 5396 37028 5460 37092
rect 6886 37020 6950 37024
rect 6886 36964 6890 37020
rect 6890 36964 6946 37020
rect 6946 36964 6950 37020
rect 6886 36960 6950 36964
rect 6966 37020 7030 37024
rect 6966 36964 6970 37020
rect 6970 36964 7026 37020
rect 7026 36964 7030 37020
rect 6966 36960 7030 36964
rect 7046 37020 7110 37024
rect 7046 36964 7050 37020
rect 7050 36964 7106 37020
rect 7106 36964 7110 37020
rect 7046 36960 7110 36964
rect 7126 37020 7190 37024
rect 7126 36964 7130 37020
rect 7130 36964 7186 37020
rect 7186 36964 7190 37020
rect 7126 36960 7190 36964
rect 12820 37020 12884 37024
rect 12820 36964 12824 37020
rect 12824 36964 12880 37020
rect 12880 36964 12884 37020
rect 12820 36960 12884 36964
rect 12900 37020 12964 37024
rect 12900 36964 12904 37020
rect 12904 36964 12960 37020
rect 12960 36964 12964 37020
rect 12900 36960 12964 36964
rect 12980 37020 13044 37024
rect 12980 36964 12984 37020
rect 12984 36964 13040 37020
rect 13040 36964 13044 37020
rect 12980 36960 13044 36964
rect 13060 37020 13124 37024
rect 13060 36964 13064 37020
rect 13064 36964 13120 37020
rect 13120 36964 13124 37020
rect 13060 36960 13124 36964
rect 18754 37020 18818 37024
rect 18754 36964 18758 37020
rect 18758 36964 18814 37020
rect 18814 36964 18818 37020
rect 18754 36960 18818 36964
rect 18834 37020 18898 37024
rect 18834 36964 18838 37020
rect 18838 36964 18894 37020
rect 18894 36964 18898 37020
rect 18834 36960 18898 36964
rect 18914 37020 18978 37024
rect 18914 36964 18918 37020
rect 18918 36964 18974 37020
rect 18974 36964 18978 37020
rect 18914 36960 18978 36964
rect 18994 37020 19058 37024
rect 18994 36964 18998 37020
rect 18998 36964 19054 37020
rect 19054 36964 19058 37020
rect 18994 36960 19058 36964
rect 24688 37020 24752 37024
rect 24688 36964 24692 37020
rect 24692 36964 24748 37020
rect 24748 36964 24752 37020
rect 24688 36960 24752 36964
rect 24768 37020 24832 37024
rect 24768 36964 24772 37020
rect 24772 36964 24828 37020
rect 24828 36964 24832 37020
rect 24768 36960 24832 36964
rect 24848 37020 24912 37024
rect 24848 36964 24852 37020
rect 24852 36964 24908 37020
rect 24908 36964 24912 37020
rect 24848 36960 24912 36964
rect 24928 37020 24992 37024
rect 24928 36964 24932 37020
rect 24932 36964 24988 37020
rect 24988 36964 24992 37020
rect 24928 36960 24992 36964
rect 8524 36756 8588 36820
rect 8340 36484 8404 36548
rect 3919 36476 3983 36480
rect 3919 36420 3923 36476
rect 3923 36420 3979 36476
rect 3979 36420 3983 36476
rect 3919 36416 3983 36420
rect 3999 36476 4063 36480
rect 3999 36420 4003 36476
rect 4003 36420 4059 36476
rect 4059 36420 4063 36476
rect 3999 36416 4063 36420
rect 4079 36476 4143 36480
rect 4079 36420 4083 36476
rect 4083 36420 4139 36476
rect 4139 36420 4143 36476
rect 4079 36416 4143 36420
rect 4159 36476 4223 36480
rect 4159 36420 4163 36476
rect 4163 36420 4219 36476
rect 4219 36420 4223 36476
rect 4159 36416 4223 36420
rect 9853 36476 9917 36480
rect 9853 36420 9857 36476
rect 9857 36420 9913 36476
rect 9913 36420 9917 36476
rect 9853 36416 9917 36420
rect 9933 36476 9997 36480
rect 9933 36420 9937 36476
rect 9937 36420 9993 36476
rect 9993 36420 9997 36476
rect 9933 36416 9997 36420
rect 10013 36476 10077 36480
rect 10013 36420 10017 36476
rect 10017 36420 10073 36476
rect 10073 36420 10077 36476
rect 10013 36416 10077 36420
rect 10093 36476 10157 36480
rect 10093 36420 10097 36476
rect 10097 36420 10153 36476
rect 10153 36420 10157 36476
rect 10093 36416 10157 36420
rect 15787 36476 15851 36480
rect 15787 36420 15791 36476
rect 15791 36420 15847 36476
rect 15847 36420 15851 36476
rect 15787 36416 15851 36420
rect 15867 36476 15931 36480
rect 15867 36420 15871 36476
rect 15871 36420 15927 36476
rect 15927 36420 15931 36476
rect 15867 36416 15931 36420
rect 15947 36476 16011 36480
rect 15947 36420 15951 36476
rect 15951 36420 16007 36476
rect 16007 36420 16011 36476
rect 15947 36416 16011 36420
rect 16027 36476 16091 36480
rect 16027 36420 16031 36476
rect 16031 36420 16087 36476
rect 16087 36420 16091 36476
rect 16027 36416 16091 36420
rect 21721 36476 21785 36480
rect 21721 36420 21725 36476
rect 21725 36420 21781 36476
rect 21781 36420 21785 36476
rect 21721 36416 21785 36420
rect 21801 36476 21865 36480
rect 21801 36420 21805 36476
rect 21805 36420 21861 36476
rect 21861 36420 21865 36476
rect 21801 36416 21865 36420
rect 21881 36476 21945 36480
rect 21881 36420 21885 36476
rect 21885 36420 21941 36476
rect 21941 36420 21945 36476
rect 21881 36416 21945 36420
rect 21961 36476 22025 36480
rect 21961 36420 21965 36476
rect 21965 36420 22021 36476
rect 22021 36420 22025 36476
rect 21961 36416 22025 36420
rect 5028 36212 5092 36276
rect 11284 36272 11348 36276
rect 11284 36216 11298 36272
rect 11298 36216 11348 36272
rect 11284 36212 11348 36216
rect 22876 35940 22940 36004
rect 6886 35932 6950 35936
rect 6886 35876 6890 35932
rect 6890 35876 6946 35932
rect 6946 35876 6950 35932
rect 6886 35872 6950 35876
rect 6966 35932 7030 35936
rect 6966 35876 6970 35932
rect 6970 35876 7026 35932
rect 7026 35876 7030 35932
rect 6966 35872 7030 35876
rect 7046 35932 7110 35936
rect 7046 35876 7050 35932
rect 7050 35876 7106 35932
rect 7106 35876 7110 35932
rect 7046 35872 7110 35876
rect 7126 35932 7190 35936
rect 7126 35876 7130 35932
rect 7130 35876 7186 35932
rect 7186 35876 7190 35932
rect 7126 35872 7190 35876
rect 12820 35932 12884 35936
rect 12820 35876 12824 35932
rect 12824 35876 12880 35932
rect 12880 35876 12884 35932
rect 12820 35872 12884 35876
rect 12900 35932 12964 35936
rect 12900 35876 12904 35932
rect 12904 35876 12960 35932
rect 12960 35876 12964 35932
rect 12900 35872 12964 35876
rect 12980 35932 13044 35936
rect 12980 35876 12984 35932
rect 12984 35876 13040 35932
rect 13040 35876 13044 35932
rect 12980 35872 13044 35876
rect 13060 35932 13124 35936
rect 13060 35876 13064 35932
rect 13064 35876 13120 35932
rect 13120 35876 13124 35932
rect 13060 35872 13124 35876
rect 18754 35932 18818 35936
rect 18754 35876 18758 35932
rect 18758 35876 18814 35932
rect 18814 35876 18818 35932
rect 18754 35872 18818 35876
rect 18834 35932 18898 35936
rect 18834 35876 18838 35932
rect 18838 35876 18894 35932
rect 18894 35876 18898 35932
rect 18834 35872 18898 35876
rect 18914 35932 18978 35936
rect 18914 35876 18918 35932
rect 18918 35876 18974 35932
rect 18974 35876 18978 35932
rect 18914 35872 18978 35876
rect 18994 35932 19058 35936
rect 18994 35876 18998 35932
rect 18998 35876 19054 35932
rect 19054 35876 19058 35932
rect 18994 35872 19058 35876
rect 24688 35932 24752 35936
rect 24688 35876 24692 35932
rect 24692 35876 24748 35932
rect 24748 35876 24752 35932
rect 24688 35872 24752 35876
rect 24768 35932 24832 35936
rect 24768 35876 24772 35932
rect 24772 35876 24828 35932
rect 24828 35876 24832 35932
rect 24768 35872 24832 35876
rect 24848 35932 24912 35936
rect 24848 35876 24852 35932
rect 24852 35876 24908 35932
rect 24908 35876 24912 35932
rect 24848 35872 24912 35876
rect 24928 35932 24992 35936
rect 24928 35876 24932 35932
rect 24932 35876 24988 35932
rect 24988 35876 24992 35932
rect 24928 35872 24992 35876
rect 4292 35804 4356 35868
rect 18276 35864 18340 35868
rect 18276 35808 18326 35864
rect 18326 35808 18340 35864
rect 18276 35804 18340 35808
rect 5948 35532 6012 35596
rect 22324 35532 22388 35596
rect 13492 35456 13556 35460
rect 13492 35400 13506 35456
rect 13506 35400 13556 35456
rect 13492 35396 13556 35400
rect 3919 35388 3983 35392
rect 3919 35332 3923 35388
rect 3923 35332 3979 35388
rect 3979 35332 3983 35388
rect 3919 35328 3983 35332
rect 3999 35388 4063 35392
rect 3999 35332 4003 35388
rect 4003 35332 4059 35388
rect 4059 35332 4063 35388
rect 3999 35328 4063 35332
rect 4079 35388 4143 35392
rect 4079 35332 4083 35388
rect 4083 35332 4139 35388
rect 4139 35332 4143 35388
rect 4079 35328 4143 35332
rect 4159 35388 4223 35392
rect 4159 35332 4163 35388
rect 4163 35332 4219 35388
rect 4219 35332 4223 35388
rect 4159 35328 4223 35332
rect 9853 35388 9917 35392
rect 9853 35332 9857 35388
rect 9857 35332 9913 35388
rect 9913 35332 9917 35388
rect 9853 35328 9917 35332
rect 9933 35388 9997 35392
rect 9933 35332 9937 35388
rect 9937 35332 9993 35388
rect 9993 35332 9997 35388
rect 9933 35328 9997 35332
rect 10013 35388 10077 35392
rect 10013 35332 10017 35388
rect 10017 35332 10073 35388
rect 10073 35332 10077 35388
rect 10013 35328 10077 35332
rect 10093 35388 10157 35392
rect 10093 35332 10097 35388
rect 10097 35332 10153 35388
rect 10153 35332 10157 35388
rect 10093 35328 10157 35332
rect 15787 35388 15851 35392
rect 15787 35332 15791 35388
rect 15791 35332 15847 35388
rect 15847 35332 15851 35388
rect 15787 35328 15851 35332
rect 15867 35388 15931 35392
rect 15867 35332 15871 35388
rect 15871 35332 15927 35388
rect 15927 35332 15931 35388
rect 15867 35328 15931 35332
rect 15947 35388 16011 35392
rect 15947 35332 15951 35388
rect 15951 35332 16007 35388
rect 16007 35332 16011 35388
rect 15947 35328 16011 35332
rect 16027 35388 16091 35392
rect 16027 35332 16031 35388
rect 16031 35332 16087 35388
rect 16087 35332 16091 35388
rect 16027 35328 16091 35332
rect 21721 35388 21785 35392
rect 21721 35332 21725 35388
rect 21725 35332 21781 35388
rect 21781 35332 21785 35388
rect 21721 35328 21785 35332
rect 21801 35388 21865 35392
rect 21801 35332 21805 35388
rect 21805 35332 21861 35388
rect 21861 35332 21865 35388
rect 21801 35328 21865 35332
rect 21881 35388 21945 35392
rect 21881 35332 21885 35388
rect 21885 35332 21941 35388
rect 21941 35332 21945 35388
rect 21881 35328 21945 35332
rect 21961 35388 22025 35392
rect 21961 35332 21965 35388
rect 21965 35332 22021 35388
rect 22021 35332 22025 35388
rect 21961 35328 22025 35332
rect 12020 35048 12084 35052
rect 12020 34992 12070 35048
rect 12070 34992 12084 35048
rect 12020 34988 12084 34992
rect 6886 34844 6950 34848
rect 6886 34788 6890 34844
rect 6890 34788 6946 34844
rect 6946 34788 6950 34844
rect 6886 34784 6950 34788
rect 6966 34844 7030 34848
rect 6966 34788 6970 34844
rect 6970 34788 7026 34844
rect 7026 34788 7030 34844
rect 6966 34784 7030 34788
rect 7046 34844 7110 34848
rect 7046 34788 7050 34844
rect 7050 34788 7106 34844
rect 7106 34788 7110 34844
rect 7046 34784 7110 34788
rect 7126 34844 7190 34848
rect 7126 34788 7130 34844
rect 7130 34788 7186 34844
rect 7186 34788 7190 34844
rect 7126 34784 7190 34788
rect 12820 34844 12884 34848
rect 12820 34788 12824 34844
rect 12824 34788 12880 34844
rect 12880 34788 12884 34844
rect 12820 34784 12884 34788
rect 12900 34844 12964 34848
rect 12900 34788 12904 34844
rect 12904 34788 12960 34844
rect 12960 34788 12964 34844
rect 12900 34784 12964 34788
rect 12980 34844 13044 34848
rect 12980 34788 12984 34844
rect 12984 34788 13040 34844
rect 13040 34788 13044 34844
rect 12980 34784 13044 34788
rect 13060 34844 13124 34848
rect 13060 34788 13064 34844
rect 13064 34788 13120 34844
rect 13120 34788 13124 34844
rect 13060 34784 13124 34788
rect 18754 34844 18818 34848
rect 18754 34788 18758 34844
rect 18758 34788 18814 34844
rect 18814 34788 18818 34844
rect 18754 34784 18818 34788
rect 18834 34844 18898 34848
rect 18834 34788 18838 34844
rect 18838 34788 18894 34844
rect 18894 34788 18898 34844
rect 18834 34784 18898 34788
rect 18914 34844 18978 34848
rect 18914 34788 18918 34844
rect 18918 34788 18974 34844
rect 18974 34788 18978 34844
rect 18914 34784 18978 34788
rect 18994 34844 19058 34848
rect 18994 34788 18998 34844
rect 18998 34788 19054 34844
rect 19054 34788 19058 34844
rect 18994 34784 19058 34788
rect 24688 34844 24752 34848
rect 24688 34788 24692 34844
rect 24692 34788 24748 34844
rect 24748 34788 24752 34844
rect 24688 34784 24752 34788
rect 24768 34844 24832 34848
rect 24768 34788 24772 34844
rect 24772 34788 24828 34844
rect 24828 34788 24832 34844
rect 24768 34784 24832 34788
rect 24848 34844 24912 34848
rect 24848 34788 24852 34844
rect 24852 34788 24908 34844
rect 24908 34788 24912 34844
rect 24848 34784 24912 34788
rect 24928 34844 24992 34848
rect 24928 34788 24932 34844
rect 24932 34788 24988 34844
rect 24988 34788 24992 34844
rect 24928 34784 24992 34788
rect 12204 34580 12268 34644
rect 3919 34300 3983 34304
rect 3919 34244 3923 34300
rect 3923 34244 3979 34300
rect 3979 34244 3983 34300
rect 3919 34240 3983 34244
rect 3999 34300 4063 34304
rect 3999 34244 4003 34300
rect 4003 34244 4059 34300
rect 4059 34244 4063 34300
rect 3999 34240 4063 34244
rect 4079 34300 4143 34304
rect 4079 34244 4083 34300
rect 4083 34244 4139 34300
rect 4139 34244 4143 34300
rect 4079 34240 4143 34244
rect 4159 34300 4223 34304
rect 4159 34244 4163 34300
rect 4163 34244 4219 34300
rect 4219 34244 4223 34300
rect 4159 34240 4223 34244
rect 9853 34300 9917 34304
rect 9853 34244 9857 34300
rect 9857 34244 9913 34300
rect 9913 34244 9917 34300
rect 9853 34240 9917 34244
rect 9933 34300 9997 34304
rect 9933 34244 9937 34300
rect 9937 34244 9993 34300
rect 9993 34244 9997 34300
rect 9933 34240 9997 34244
rect 10013 34300 10077 34304
rect 10013 34244 10017 34300
rect 10017 34244 10073 34300
rect 10073 34244 10077 34300
rect 10013 34240 10077 34244
rect 10093 34300 10157 34304
rect 10093 34244 10097 34300
rect 10097 34244 10153 34300
rect 10153 34244 10157 34300
rect 10093 34240 10157 34244
rect 15787 34300 15851 34304
rect 15787 34244 15791 34300
rect 15791 34244 15847 34300
rect 15847 34244 15851 34300
rect 15787 34240 15851 34244
rect 15867 34300 15931 34304
rect 15867 34244 15871 34300
rect 15871 34244 15927 34300
rect 15927 34244 15931 34300
rect 15867 34240 15931 34244
rect 15947 34300 16011 34304
rect 15947 34244 15951 34300
rect 15951 34244 16007 34300
rect 16007 34244 16011 34300
rect 15947 34240 16011 34244
rect 16027 34300 16091 34304
rect 16027 34244 16031 34300
rect 16031 34244 16087 34300
rect 16087 34244 16091 34300
rect 16027 34240 16091 34244
rect 21721 34300 21785 34304
rect 21721 34244 21725 34300
rect 21725 34244 21781 34300
rect 21781 34244 21785 34300
rect 21721 34240 21785 34244
rect 21801 34300 21865 34304
rect 21801 34244 21805 34300
rect 21805 34244 21861 34300
rect 21861 34244 21865 34300
rect 21801 34240 21865 34244
rect 21881 34300 21945 34304
rect 21881 34244 21885 34300
rect 21885 34244 21941 34300
rect 21941 34244 21945 34300
rect 21881 34240 21945 34244
rect 21961 34300 22025 34304
rect 21961 34244 21965 34300
rect 21965 34244 22021 34300
rect 22021 34244 22025 34300
rect 21961 34240 22025 34244
rect 10548 34036 10612 34100
rect 6886 33756 6950 33760
rect 6886 33700 6890 33756
rect 6890 33700 6946 33756
rect 6946 33700 6950 33756
rect 6886 33696 6950 33700
rect 6966 33756 7030 33760
rect 6966 33700 6970 33756
rect 6970 33700 7026 33756
rect 7026 33700 7030 33756
rect 6966 33696 7030 33700
rect 7046 33756 7110 33760
rect 7046 33700 7050 33756
rect 7050 33700 7106 33756
rect 7106 33700 7110 33756
rect 7046 33696 7110 33700
rect 7126 33756 7190 33760
rect 7126 33700 7130 33756
rect 7130 33700 7186 33756
rect 7186 33700 7190 33756
rect 7126 33696 7190 33700
rect 12820 33756 12884 33760
rect 12820 33700 12824 33756
rect 12824 33700 12880 33756
rect 12880 33700 12884 33756
rect 12820 33696 12884 33700
rect 12900 33756 12964 33760
rect 12900 33700 12904 33756
rect 12904 33700 12960 33756
rect 12960 33700 12964 33756
rect 12900 33696 12964 33700
rect 12980 33756 13044 33760
rect 12980 33700 12984 33756
rect 12984 33700 13040 33756
rect 13040 33700 13044 33756
rect 12980 33696 13044 33700
rect 13060 33756 13124 33760
rect 13060 33700 13064 33756
rect 13064 33700 13120 33756
rect 13120 33700 13124 33756
rect 13060 33696 13124 33700
rect 18754 33756 18818 33760
rect 18754 33700 18758 33756
rect 18758 33700 18814 33756
rect 18814 33700 18818 33756
rect 18754 33696 18818 33700
rect 18834 33756 18898 33760
rect 18834 33700 18838 33756
rect 18838 33700 18894 33756
rect 18894 33700 18898 33756
rect 18834 33696 18898 33700
rect 18914 33756 18978 33760
rect 18914 33700 18918 33756
rect 18918 33700 18974 33756
rect 18974 33700 18978 33756
rect 18914 33696 18978 33700
rect 18994 33756 19058 33760
rect 18994 33700 18998 33756
rect 18998 33700 19054 33756
rect 19054 33700 19058 33756
rect 18994 33696 19058 33700
rect 24688 33756 24752 33760
rect 24688 33700 24692 33756
rect 24692 33700 24748 33756
rect 24748 33700 24752 33756
rect 24688 33696 24752 33700
rect 24768 33756 24832 33760
rect 24768 33700 24772 33756
rect 24772 33700 24828 33756
rect 24828 33700 24832 33756
rect 24768 33696 24832 33700
rect 24848 33756 24912 33760
rect 24848 33700 24852 33756
rect 24852 33700 24908 33756
rect 24908 33700 24912 33756
rect 24848 33696 24912 33700
rect 24928 33756 24992 33760
rect 24928 33700 24932 33756
rect 24932 33700 24988 33756
rect 24988 33700 24992 33756
rect 24928 33696 24992 33700
rect 22692 33220 22756 33284
rect 3919 33212 3983 33216
rect 3919 33156 3923 33212
rect 3923 33156 3979 33212
rect 3979 33156 3983 33212
rect 3919 33152 3983 33156
rect 3999 33212 4063 33216
rect 3999 33156 4003 33212
rect 4003 33156 4059 33212
rect 4059 33156 4063 33212
rect 3999 33152 4063 33156
rect 4079 33212 4143 33216
rect 4079 33156 4083 33212
rect 4083 33156 4139 33212
rect 4139 33156 4143 33212
rect 4079 33152 4143 33156
rect 4159 33212 4223 33216
rect 4159 33156 4163 33212
rect 4163 33156 4219 33212
rect 4219 33156 4223 33212
rect 4159 33152 4223 33156
rect 9853 33212 9917 33216
rect 9853 33156 9857 33212
rect 9857 33156 9913 33212
rect 9913 33156 9917 33212
rect 9853 33152 9917 33156
rect 9933 33212 9997 33216
rect 9933 33156 9937 33212
rect 9937 33156 9993 33212
rect 9993 33156 9997 33212
rect 9933 33152 9997 33156
rect 10013 33212 10077 33216
rect 10013 33156 10017 33212
rect 10017 33156 10073 33212
rect 10073 33156 10077 33212
rect 10013 33152 10077 33156
rect 10093 33212 10157 33216
rect 10093 33156 10097 33212
rect 10097 33156 10153 33212
rect 10153 33156 10157 33212
rect 10093 33152 10157 33156
rect 15787 33212 15851 33216
rect 15787 33156 15791 33212
rect 15791 33156 15847 33212
rect 15847 33156 15851 33212
rect 15787 33152 15851 33156
rect 15867 33212 15931 33216
rect 15867 33156 15871 33212
rect 15871 33156 15927 33212
rect 15927 33156 15931 33212
rect 15867 33152 15931 33156
rect 15947 33212 16011 33216
rect 15947 33156 15951 33212
rect 15951 33156 16007 33212
rect 16007 33156 16011 33212
rect 15947 33152 16011 33156
rect 16027 33212 16091 33216
rect 16027 33156 16031 33212
rect 16031 33156 16087 33212
rect 16087 33156 16091 33212
rect 16027 33152 16091 33156
rect 21721 33212 21785 33216
rect 21721 33156 21725 33212
rect 21725 33156 21781 33212
rect 21781 33156 21785 33212
rect 21721 33152 21785 33156
rect 21801 33212 21865 33216
rect 21801 33156 21805 33212
rect 21805 33156 21861 33212
rect 21861 33156 21865 33212
rect 21801 33152 21865 33156
rect 21881 33212 21945 33216
rect 21881 33156 21885 33212
rect 21885 33156 21941 33212
rect 21941 33156 21945 33212
rect 21881 33152 21945 33156
rect 21961 33212 22025 33216
rect 21961 33156 21965 33212
rect 21965 33156 22021 33212
rect 22021 33156 22025 33212
rect 21961 33152 22025 33156
rect 18092 33084 18156 33148
rect 11652 32948 11716 33012
rect 4660 32676 4724 32740
rect 11284 32736 11348 32740
rect 11284 32680 11298 32736
rect 11298 32680 11348 32736
rect 11284 32676 11348 32680
rect 6886 32668 6950 32672
rect 6886 32612 6890 32668
rect 6890 32612 6946 32668
rect 6946 32612 6950 32668
rect 6886 32608 6950 32612
rect 6966 32668 7030 32672
rect 6966 32612 6970 32668
rect 6970 32612 7026 32668
rect 7026 32612 7030 32668
rect 6966 32608 7030 32612
rect 7046 32668 7110 32672
rect 7046 32612 7050 32668
rect 7050 32612 7106 32668
rect 7106 32612 7110 32668
rect 7046 32608 7110 32612
rect 7126 32668 7190 32672
rect 7126 32612 7130 32668
rect 7130 32612 7186 32668
rect 7186 32612 7190 32668
rect 7126 32608 7190 32612
rect 12820 32668 12884 32672
rect 12820 32612 12824 32668
rect 12824 32612 12880 32668
rect 12880 32612 12884 32668
rect 12820 32608 12884 32612
rect 12900 32668 12964 32672
rect 12900 32612 12904 32668
rect 12904 32612 12960 32668
rect 12960 32612 12964 32668
rect 12900 32608 12964 32612
rect 12980 32668 13044 32672
rect 12980 32612 12984 32668
rect 12984 32612 13040 32668
rect 13040 32612 13044 32668
rect 12980 32608 13044 32612
rect 13060 32668 13124 32672
rect 13060 32612 13064 32668
rect 13064 32612 13120 32668
rect 13120 32612 13124 32668
rect 13060 32608 13124 32612
rect 18754 32668 18818 32672
rect 18754 32612 18758 32668
rect 18758 32612 18814 32668
rect 18814 32612 18818 32668
rect 18754 32608 18818 32612
rect 18834 32668 18898 32672
rect 18834 32612 18838 32668
rect 18838 32612 18894 32668
rect 18894 32612 18898 32668
rect 18834 32608 18898 32612
rect 18914 32668 18978 32672
rect 18914 32612 18918 32668
rect 18918 32612 18974 32668
rect 18974 32612 18978 32668
rect 18914 32608 18978 32612
rect 18994 32668 19058 32672
rect 18994 32612 18998 32668
rect 18998 32612 19054 32668
rect 19054 32612 19058 32668
rect 18994 32608 19058 32612
rect 24688 32668 24752 32672
rect 24688 32612 24692 32668
rect 24692 32612 24748 32668
rect 24748 32612 24752 32668
rect 24688 32608 24752 32612
rect 24768 32668 24832 32672
rect 24768 32612 24772 32668
rect 24772 32612 24828 32668
rect 24828 32612 24832 32668
rect 24768 32608 24832 32612
rect 24848 32668 24912 32672
rect 24848 32612 24852 32668
rect 24852 32612 24908 32668
rect 24908 32612 24912 32668
rect 24848 32608 24912 32612
rect 24928 32668 24992 32672
rect 24928 32612 24932 32668
rect 24932 32612 24988 32668
rect 24988 32612 24992 32668
rect 24928 32608 24992 32612
rect 2636 32540 2700 32604
rect 3188 32404 3252 32468
rect 3556 32268 3620 32332
rect 11836 32268 11900 32332
rect 3919 32124 3983 32128
rect 3919 32068 3923 32124
rect 3923 32068 3979 32124
rect 3979 32068 3983 32124
rect 3919 32064 3983 32068
rect 3999 32124 4063 32128
rect 3999 32068 4003 32124
rect 4003 32068 4059 32124
rect 4059 32068 4063 32124
rect 3999 32064 4063 32068
rect 4079 32124 4143 32128
rect 4079 32068 4083 32124
rect 4083 32068 4139 32124
rect 4139 32068 4143 32124
rect 4079 32064 4143 32068
rect 4159 32124 4223 32128
rect 4159 32068 4163 32124
rect 4163 32068 4219 32124
rect 4219 32068 4223 32124
rect 4159 32064 4223 32068
rect 9853 32124 9917 32128
rect 9853 32068 9857 32124
rect 9857 32068 9913 32124
rect 9913 32068 9917 32124
rect 9853 32064 9917 32068
rect 9933 32124 9997 32128
rect 9933 32068 9937 32124
rect 9937 32068 9993 32124
rect 9993 32068 9997 32124
rect 9933 32064 9997 32068
rect 10013 32124 10077 32128
rect 10013 32068 10017 32124
rect 10017 32068 10073 32124
rect 10073 32068 10077 32124
rect 10013 32064 10077 32068
rect 10093 32124 10157 32128
rect 10093 32068 10097 32124
rect 10097 32068 10153 32124
rect 10153 32068 10157 32124
rect 10093 32064 10157 32068
rect 15787 32124 15851 32128
rect 15787 32068 15791 32124
rect 15791 32068 15847 32124
rect 15847 32068 15851 32124
rect 15787 32064 15851 32068
rect 15867 32124 15931 32128
rect 15867 32068 15871 32124
rect 15871 32068 15927 32124
rect 15927 32068 15931 32124
rect 15867 32064 15931 32068
rect 15947 32124 16011 32128
rect 15947 32068 15951 32124
rect 15951 32068 16007 32124
rect 16007 32068 16011 32124
rect 15947 32064 16011 32068
rect 16027 32124 16091 32128
rect 16027 32068 16031 32124
rect 16031 32068 16087 32124
rect 16087 32068 16091 32124
rect 16027 32064 16091 32068
rect 21721 32124 21785 32128
rect 21721 32068 21725 32124
rect 21725 32068 21781 32124
rect 21781 32068 21785 32124
rect 21721 32064 21785 32068
rect 21801 32124 21865 32128
rect 21801 32068 21805 32124
rect 21805 32068 21861 32124
rect 21861 32068 21865 32124
rect 21801 32064 21865 32068
rect 21881 32124 21945 32128
rect 21881 32068 21885 32124
rect 21885 32068 21941 32124
rect 21941 32068 21945 32124
rect 21881 32064 21945 32068
rect 21961 32124 22025 32128
rect 21961 32068 21965 32124
rect 21965 32068 22021 32124
rect 22021 32068 22025 32124
rect 21961 32064 22025 32068
rect 4292 31860 4356 31924
rect 5396 31860 5460 31924
rect 23244 31784 23308 31788
rect 23244 31728 23258 31784
rect 23258 31728 23308 31784
rect 23244 31724 23308 31728
rect 8524 31588 8588 31652
rect 6886 31580 6950 31584
rect 6886 31524 6890 31580
rect 6890 31524 6946 31580
rect 6946 31524 6950 31580
rect 6886 31520 6950 31524
rect 6966 31580 7030 31584
rect 6966 31524 6970 31580
rect 6970 31524 7026 31580
rect 7026 31524 7030 31580
rect 6966 31520 7030 31524
rect 7046 31580 7110 31584
rect 7046 31524 7050 31580
rect 7050 31524 7106 31580
rect 7106 31524 7110 31580
rect 7046 31520 7110 31524
rect 7126 31580 7190 31584
rect 7126 31524 7130 31580
rect 7130 31524 7186 31580
rect 7186 31524 7190 31580
rect 7126 31520 7190 31524
rect 12820 31580 12884 31584
rect 12820 31524 12824 31580
rect 12824 31524 12880 31580
rect 12880 31524 12884 31580
rect 12820 31520 12884 31524
rect 12900 31580 12964 31584
rect 12900 31524 12904 31580
rect 12904 31524 12960 31580
rect 12960 31524 12964 31580
rect 12900 31520 12964 31524
rect 12980 31580 13044 31584
rect 12980 31524 12984 31580
rect 12984 31524 13040 31580
rect 13040 31524 13044 31580
rect 12980 31520 13044 31524
rect 13060 31580 13124 31584
rect 13060 31524 13064 31580
rect 13064 31524 13120 31580
rect 13120 31524 13124 31580
rect 13060 31520 13124 31524
rect 18754 31580 18818 31584
rect 18754 31524 18758 31580
rect 18758 31524 18814 31580
rect 18814 31524 18818 31580
rect 18754 31520 18818 31524
rect 18834 31580 18898 31584
rect 18834 31524 18838 31580
rect 18838 31524 18894 31580
rect 18894 31524 18898 31580
rect 18834 31520 18898 31524
rect 18914 31580 18978 31584
rect 18914 31524 18918 31580
rect 18918 31524 18974 31580
rect 18974 31524 18978 31580
rect 18914 31520 18978 31524
rect 18994 31580 19058 31584
rect 18994 31524 18998 31580
rect 18998 31524 19054 31580
rect 19054 31524 19058 31580
rect 18994 31520 19058 31524
rect 24688 31580 24752 31584
rect 24688 31524 24692 31580
rect 24692 31524 24748 31580
rect 24748 31524 24752 31580
rect 24688 31520 24752 31524
rect 24768 31580 24832 31584
rect 24768 31524 24772 31580
rect 24772 31524 24828 31580
rect 24828 31524 24832 31580
rect 24768 31520 24832 31524
rect 24848 31580 24912 31584
rect 24848 31524 24852 31580
rect 24852 31524 24908 31580
rect 24908 31524 24912 31580
rect 24848 31520 24912 31524
rect 24928 31580 24992 31584
rect 24928 31524 24932 31580
rect 24932 31524 24988 31580
rect 24988 31524 24992 31580
rect 24928 31520 24992 31524
rect 3919 31036 3983 31040
rect 3919 30980 3923 31036
rect 3923 30980 3979 31036
rect 3979 30980 3983 31036
rect 3919 30976 3983 30980
rect 3999 31036 4063 31040
rect 3999 30980 4003 31036
rect 4003 30980 4059 31036
rect 4059 30980 4063 31036
rect 3999 30976 4063 30980
rect 4079 31036 4143 31040
rect 4079 30980 4083 31036
rect 4083 30980 4139 31036
rect 4139 30980 4143 31036
rect 4079 30976 4143 30980
rect 4159 31036 4223 31040
rect 4159 30980 4163 31036
rect 4163 30980 4219 31036
rect 4219 30980 4223 31036
rect 4159 30976 4223 30980
rect 9853 31036 9917 31040
rect 9853 30980 9857 31036
rect 9857 30980 9913 31036
rect 9913 30980 9917 31036
rect 9853 30976 9917 30980
rect 9933 31036 9997 31040
rect 9933 30980 9937 31036
rect 9937 30980 9993 31036
rect 9993 30980 9997 31036
rect 9933 30976 9997 30980
rect 10013 31036 10077 31040
rect 10013 30980 10017 31036
rect 10017 30980 10073 31036
rect 10073 30980 10077 31036
rect 10013 30976 10077 30980
rect 10093 31036 10157 31040
rect 10093 30980 10097 31036
rect 10097 30980 10153 31036
rect 10153 30980 10157 31036
rect 10093 30976 10157 30980
rect 1900 30772 1964 30836
rect 2636 30696 2700 30700
rect 13492 31044 13556 31108
rect 15787 31036 15851 31040
rect 15787 30980 15791 31036
rect 15791 30980 15847 31036
rect 15847 30980 15851 31036
rect 15787 30976 15851 30980
rect 15867 31036 15931 31040
rect 15867 30980 15871 31036
rect 15871 30980 15927 31036
rect 15927 30980 15931 31036
rect 15867 30976 15931 30980
rect 15947 31036 16011 31040
rect 15947 30980 15951 31036
rect 15951 30980 16007 31036
rect 16007 30980 16011 31036
rect 15947 30976 16011 30980
rect 16027 31036 16091 31040
rect 16027 30980 16031 31036
rect 16031 30980 16087 31036
rect 16087 30980 16091 31036
rect 16027 30976 16091 30980
rect 21721 31036 21785 31040
rect 21721 30980 21725 31036
rect 21725 30980 21781 31036
rect 21781 30980 21785 31036
rect 21721 30976 21785 30980
rect 21801 31036 21865 31040
rect 21801 30980 21805 31036
rect 21805 30980 21861 31036
rect 21861 30980 21865 31036
rect 21801 30976 21865 30980
rect 21881 31036 21945 31040
rect 21881 30980 21885 31036
rect 21885 30980 21941 31036
rect 21941 30980 21945 31036
rect 21881 30976 21945 30980
rect 21961 31036 22025 31040
rect 21961 30980 21965 31036
rect 21965 30980 22021 31036
rect 22021 30980 22025 31036
rect 21961 30976 22025 30980
rect 14228 30772 14292 30836
rect 16988 30772 17052 30836
rect 2636 30640 2650 30696
rect 2650 30640 2700 30696
rect 2636 30636 2700 30640
rect 8524 30636 8588 30700
rect 9260 30696 9324 30700
rect 9260 30640 9274 30696
rect 9274 30640 9324 30696
rect 9260 30636 9324 30640
rect 9444 30636 9508 30700
rect 10364 30636 10428 30700
rect 10548 30696 10612 30700
rect 10548 30640 10598 30696
rect 10598 30640 10612 30696
rect 10548 30636 10612 30640
rect 16988 30636 17052 30700
rect 2084 30364 2148 30428
rect 6886 30492 6950 30496
rect 6886 30436 6890 30492
rect 6890 30436 6946 30492
rect 6946 30436 6950 30492
rect 6886 30432 6950 30436
rect 6966 30492 7030 30496
rect 6966 30436 6970 30492
rect 6970 30436 7026 30492
rect 7026 30436 7030 30492
rect 6966 30432 7030 30436
rect 7046 30492 7110 30496
rect 7046 30436 7050 30492
rect 7050 30436 7106 30492
rect 7106 30436 7110 30492
rect 7046 30432 7110 30436
rect 7126 30492 7190 30496
rect 7126 30436 7130 30492
rect 7130 30436 7186 30492
rect 7186 30436 7190 30492
rect 7126 30432 7190 30436
rect 12820 30492 12884 30496
rect 12820 30436 12824 30492
rect 12824 30436 12880 30492
rect 12880 30436 12884 30492
rect 12820 30432 12884 30436
rect 12900 30492 12964 30496
rect 12900 30436 12904 30492
rect 12904 30436 12960 30492
rect 12960 30436 12964 30492
rect 12900 30432 12964 30436
rect 12980 30492 13044 30496
rect 12980 30436 12984 30492
rect 12984 30436 13040 30492
rect 13040 30436 13044 30492
rect 12980 30432 13044 30436
rect 13060 30492 13124 30496
rect 13060 30436 13064 30492
rect 13064 30436 13120 30492
rect 13120 30436 13124 30492
rect 13060 30432 13124 30436
rect 18754 30492 18818 30496
rect 18754 30436 18758 30492
rect 18758 30436 18814 30492
rect 18814 30436 18818 30492
rect 18754 30432 18818 30436
rect 18834 30492 18898 30496
rect 18834 30436 18838 30492
rect 18838 30436 18894 30492
rect 18894 30436 18898 30492
rect 18834 30432 18898 30436
rect 18914 30492 18978 30496
rect 18914 30436 18918 30492
rect 18918 30436 18974 30492
rect 18974 30436 18978 30492
rect 18914 30432 18978 30436
rect 18994 30492 19058 30496
rect 18994 30436 18998 30492
rect 18998 30436 19054 30492
rect 19054 30436 19058 30492
rect 18994 30432 19058 30436
rect 24688 30492 24752 30496
rect 24688 30436 24692 30492
rect 24692 30436 24748 30492
rect 24748 30436 24752 30492
rect 24688 30432 24752 30436
rect 24768 30492 24832 30496
rect 24768 30436 24772 30492
rect 24772 30436 24828 30492
rect 24828 30436 24832 30492
rect 24768 30432 24832 30436
rect 24848 30492 24912 30496
rect 24848 30436 24852 30492
rect 24852 30436 24908 30492
rect 24908 30436 24912 30492
rect 24848 30432 24912 30436
rect 24928 30492 24992 30496
rect 24928 30436 24932 30492
rect 24932 30436 24988 30492
rect 24988 30436 24992 30492
rect 24928 30432 24992 30436
rect 8340 30364 8404 30428
rect 8708 30364 8772 30428
rect 10916 30228 10980 30292
rect 6132 29956 6196 30020
rect 3919 29948 3983 29952
rect 3919 29892 3923 29948
rect 3923 29892 3979 29948
rect 3979 29892 3983 29948
rect 3919 29888 3983 29892
rect 3999 29948 4063 29952
rect 3999 29892 4003 29948
rect 4003 29892 4059 29948
rect 4059 29892 4063 29948
rect 3999 29888 4063 29892
rect 4079 29948 4143 29952
rect 4079 29892 4083 29948
rect 4083 29892 4139 29948
rect 4139 29892 4143 29948
rect 4079 29888 4143 29892
rect 4159 29948 4223 29952
rect 4159 29892 4163 29948
rect 4163 29892 4219 29948
rect 4219 29892 4223 29948
rect 4159 29888 4223 29892
rect 9853 29948 9917 29952
rect 9853 29892 9857 29948
rect 9857 29892 9913 29948
rect 9913 29892 9917 29948
rect 9853 29888 9917 29892
rect 9933 29948 9997 29952
rect 9933 29892 9937 29948
rect 9937 29892 9993 29948
rect 9993 29892 9997 29948
rect 9933 29888 9997 29892
rect 10013 29948 10077 29952
rect 10013 29892 10017 29948
rect 10017 29892 10073 29948
rect 10073 29892 10077 29948
rect 10013 29888 10077 29892
rect 10093 29948 10157 29952
rect 10093 29892 10097 29948
rect 10097 29892 10153 29948
rect 10153 29892 10157 29948
rect 10093 29888 10157 29892
rect 15787 29948 15851 29952
rect 15787 29892 15791 29948
rect 15791 29892 15847 29948
rect 15847 29892 15851 29948
rect 15787 29888 15851 29892
rect 15867 29948 15931 29952
rect 15867 29892 15871 29948
rect 15871 29892 15927 29948
rect 15927 29892 15931 29948
rect 15867 29888 15931 29892
rect 15947 29948 16011 29952
rect 15947 29892 15951 29948
rect 15951 29892 16007 29948
rect 16007 29892 16011 29948
rect 15947 29888 16011 29892
rect 16027 29948 16091 29952
rect 16027 29892 16031 29948
rect 16031 29892 16087 29948
rect 16087 29892 16091 29948
rect 16027 29888 16091 29892
rect 21721 29948 21785 29952
rect 21721 29892 21725 29948
rect 21725 29892 21781 29948
rect 21781 29892 21785 29948
rect 21721 29888 21785 29892
rect 21801 29948 21865 29952
rect 21801 29892 21805 29948
rect 21805 29892 21861 29948
rect 21861 29892 21865 29948
rect 21801 29888 21865 29892
rect 21881 29948 21945 29952
rect 21881 29892 21885 29948
rect 21885 29892 21941 29948
rect 21941 29892 21945 29948
rect 21881 29888 21945 29892
rect 21961 29948 22025 29952
rect 21961 29892 21965 29948
rect 21965 29892 22021 29948
rect 22021 29892 22025 29948
rect 21961 29888 22025 29892
rect 6886 29404 6950 29408
rect 6886 29348 6890 29404
rect 6890 29348 6946 29404
rect 6946 29348 6950 29404
rect 6886 29344 6950 29348
rect 6966 29404 7030 29408
rect 6966 29348 6970 29404
rect 6970 29348 7026 29404
rect 7026 29348 7030 29404
rect 6966 29344 7030 29348
rect 7046 29404 7110 29408
rect 7046 29348 7050 29404
rect 7050 29348 7106 29404
rect 7106 29348 7110 29404
rect 7046 29344 7110 29348
rect 7126 29404 7190 29408
rect 7126 29348 7130 29404
rect 7130 29348 7186 29404
rect 7186 29348 7190 29404
rect 7126 29344 7190 29348
rect 4292 29140 4356 29204
rect 5028 29064 5092 29068
rect 5028 29008 5078 29064
rect 5078 29008 5092 29064
rect 5028 29004 5092 29008
rect 11836 29064 11900 29068
rect 16620 29412 16684 29476
rect 17724 29684 17788 29748
rect 12820 29404 12884 29408
rect 12820 29348 12824 29404
rect 12824 29348 12880 29404
rect 12880 29348 12884 29404
rect 12820 29344 12884 29348
rect 12900 29404 12964 29408
rect 12900 29348 12904 29404
rect 12904 29348 12960 29404
rect 12960 29348 12964 29404
rect 12900 29344 12964 29348
rect 12980 29404 13044 29408
rect 12980 29348 12984 29404
rect 12984 29348 13040 29404
rect 13040 29348 13044 29404
rect 12980 29344 13044 29348
rect 13060 29404 13124 29408
rect 13060 29348 13064 29404
rect 13064 29348 13120 29404
rect 13120 29348 13124 29404
rect 13060 29344 13124 29348
rect 18754 29404 18818 29408
rect 18754 29348 18758 29404
rect 18758 29348 18814 29404
rect 18814 29348 18818 29404
rect 18754 29344 18818 29348
rect 18834 29404 18898 29408
rect 18834 29348 18838 29404
rect 18838 29348 18894 29404
rect 18894 29348 18898 29404
rect 18834 29344 18898 29348
rect 18914 29404 18978 29408
rect 18914 29348 18918 29404
rect 18918 29348 18974 29404
rect 18974 29348 18978 29404
rect 18914 29344 18978 29348
rect 18994 29404 19058 29408
rect 18994 29348 18998 29404
rect 18998 29348 19054 29404
rect 19054 29348 19058 29404
rect 18994 29344 19058 29348
rect 24688 29404 24752 29408
rect 24688 29348 24692 29404
rect 24692 29348 24748 29404
rect 24748 29348 24752 29404
rect 24688 29344 24752 29348
rect 24768 29404 24832 29408
rect 24768 29348 24772 29404
rect 24772 29348 24828 29404
rect 24828 29348 24832 29404
rect 24768 29344 24832 29348
rect 24848 29404 24912 29408
rect 24848 29348 24852 29404
rect 24852 29348 24908 29404
rect 24908 29348 24912 29404
rect 24848 29344 24912 29348
rect 24928 29404 24992 29408
rect 24928 29348 24932 29404
rect 24932 29348 24988 29404
rect 24988 29348 24992 29404
rect 24928 29344 24992 29348
rect 11836 29008 11850 29064
rect 11850 29008 11900 29064
rect 11836 29004 11900 29008
rect 20852 29004 20916 29068
rect 10916 28868 10980 28932
rect 3919 28860 3983 28864
rect 3919 28804 3923 28860
rect 3923 28804 3979 28860
rect 3979 28804 3983 28860
rect 3919 28800 3983 28804
rect 3999 28860 4063 28864
rect 3999 28804 4003 28860
rect 4003 28804 4059 28860
rect 4059 28804 4063 28860
rect 3999 28800 4063 28804
rect 4079 28860 4143 28864
rect 4079 28804 4083 28860
rect 4083 28804 4139 28860
rect 4139 28804 4143 28860
rect 4079 28800 4143 28804
rect 4159 28860 4223 28864
rect 4159 28804 4163 28860
rect 4163 28804 4219 28860
rect 4219 28804 4223 28860
rect 4159 28800 4223 28804
rect 9853 28860 9917 28864
rect 9853 28804 9857 28860
rect 9857 28804 9913 28860
rect 9913 28804 9917 28860
rect 9853 28800 9917 28804
rect 9933 28860 9997 28864
rect 9933 28804 9937 28860
rect 9937 28804 9993 28860
rect 9993 28804 9997 28860
rect 9933 28800 9997 28804
rect 10013 28860 10077 28864
rect 10013 28804 10017 28860
rect 10017 28804 10073 28860
rect 10073 28804 10077 28860
rect 10013 28800 10077 28804
rect 10093 28860 10157 28864
rect 10093 28804 10097 28860
rect 10097 28804 10153 28860
rect 10153 28804 10157 28860
rect 10093 28800 10157 28804
rect 15787 28860 15851 28864
rect 15787 28804 15791 28860
rect 15791 28804 15847 28860
rect 15847 28804 15851 28860
rect 15787 28800 15851 28804
rect 15867 28860 15931 28864
rect 15867 28804 15871 28860
rect 15871 28804 15927 28860
rect 15927 28804 15931 28860
rect 15867 28800 15931 28804
rect 15947 28860 16011 28864
rect 15947 28804 15951 28860
rect 15951 28804 16007 28860
rect 16007 28804 16011 28860
rect 15947 28800 16011 28804
rect 16027 28860 16091 28864
rect 16027 28804 16031 28860
rect 16031 28804 16087 28860
rect 16087 28804 16091 28860
rect 16027 28800 16091 28804
rect 21721 28860 21785 28864
rect 21721 28804 21725 28860
rect 21725 28804 21781 28860
rect 21781 28804 21785 28860
rect 21721 28800 21785 28804
rect 21801 28860 21865 28864
rect 21801 28804 21805 28860
rect 21805 28804 21861 28860
rect 21861 28804 21865 28860
rect 21801 28800 21865 28804
rect 21881 28860 21945 28864
rect 21881 28804 21885 28860
rect 21885 28804 21941 28860
rect 21941 28804 21945 28860
rect 21881 28800 21945 28804
rect 21961 28860 22025 28864
rect 21961 28804 21965 28860
rect 21965 28804 22021 28860
rect 22021 28804 22025 28860
rect 21961 28800 22025 28804
rect 4476 28732 4540 28796
rect 2084 28596 2148 28660
rect 4660 28596 4724 28660
rect 2452 28460 2516 28524
rect 8892 28460 8956 28524
rect 13676 28460 13740 28524
rect 6886 28316 6950 28320
rect 6886 28260 6890 28316
rect 6890 28260 6946 28316
rect 6946 28260 6950 28316
rect 6886 28256 6950 28260
rect 6966 28316 7030 28320
rect 6966 28260 6970 28316
rect 6970 28260 7026 28316
rect 7026 28260 7030 28316
rect 6966 28256 7030 28260
rect 7046 28316 7110 28320
rect 7046 28260 7050 28316
rect 7050 28260 7106 28316
rect 7106 28260 7110 28316
rect 7046 28256 7110 28260
rect 7126 28316 7190 28320
rect 7126 28260 7130 28316
rect 7130 28260 7186 28316
rect 7186 28260 7190 28316
rect 7126 28256 7190 28260
rect 12820 28316 12884 28320
rect 12820 28260 12824 28316
rect 12824 28260 12880 28316
rect 12880 28260 12884 28316
rect 12820 28256 12884 28260
rect 12900 28316 12964 28320
rect 12900 28260 12904 28316
rect 12904 28260 12960 28316
rect 12960 28260 12964 28316
rect 12900 28256 12964 28260
rect 12980 28316 13044 28320
rect 12980 28260 12984 28316
rect 12984 28260 13040 28316
rect 13040 28260 13044 28316
rect 12980 28256 13044 28260
rect 13060 28316 13124 28320
rect 13060 28260 13064 28316
rect 13064 28260 13120 28316
rect 13120 28260 13124 28316
rect 13060 28256 13124 28260
rect 18754 28316 18818 28320
rect 18754 28260 18758 28316
rect 18758 28260 18814 28316
rect 18814 28260 18818 28316
rect 18754 28256 18818 28260
rect 18834 28316 18898 28320
rect 18834 28260 18838 28316
rect 18838 28260 18894 28316
rect 18894 28260 18898 28316
rect 18834 28256 18898 28260
rect 18914 28316 18978 28320
rect 18914 28260 18918 28316
rect 18918 28260 18974 28316
rect 18974 28260 18978 28316
rect 18914 28256 18978 28260
rect 18994 28316 19058 28320
rect 18994 28260 18998 28316
rect 18998 28260 19054 28316
rect 19054 28260 19058 28316
rect 18994 28256 19058 28260
rect 24688 28316 24752 28320
rect 24688 28260 24692 28316
rect 24692 28260 24748 28316
rect 24748 28260 24752 28316
rect 24688 28256 24752 28260
rect 24768 28316 24832 28320
rect 24768 28260 24772 28316
rect 24772 28260 24828 28316
rect 24828 28260 24832 28316
rect 24768 28256 24832 28260
rect 24848 28316 24912 28320
rect 24848 28260 24852 28316
rect 24852 28260 24908 28316
rect 24908 28260 24912 28316
rect 24848 28256 24912 28260
rect 24928 28316 24992 28320
rect 24928 28260 24932 28316
rect 24932 28260 24988 28316
rect 24988 28260 24992 28316
rect 24928 28256 24992 28260
rect 1716 27916 1780 27980
rect 3919 27772 3983 27776
rect 3919 27716 3923 27772
rect 3923 27716 3979 27772
rect 3979 27716 3983 27772
rect 3919 27712 3983 27716
rect 3999 27772 4063 27776
rect 3999 27716 4003 27772
rect 4003 27716 4059 27772
rect 4059 27716 4063 27772
rect 3999 27712 4063 27716
rect 4079 27772 4143 27776
rect 4079 27716 4083 27772
rect 4083 27716 4139 27772
rect 4139 27716 4143 27772
rect 4079 27712 4143 27716
rect 4159 27772 4223 27776
rect 4159 27716 4163 27772
rect 4163 27716 4219 27772
rect 4219 27716 4223 27772
rect 4159 27712 4223 27716
rect 9853 27772 9917 27776
rect 9853 27716 9857 27772
rect 9857 27716 9913 27772
rect 9913 27716 9917 27772
rect 9853 27712 9917 27716
rect 9933 27772 9997 27776
rect 9933 27716 9937 27772
rect 9937 27716 9993 27772
rect 9993 27716 9997 27772
rect 9933 27712 9997 27716
rect 10013 27772 10077 27776
rect 10013 27716 10017 27772
rect 10017 27716 10073 27772
rect 10073 27716 10077 27772
rect 10013 27712 10077 27716
rect 10093 27772 10157 27776
rect 10093 27716 10097 27772
rect 10097 27716 10153 27772
rect 10153 27716 10157 27772
rect 10093 27712 10157 27716
rect 15787 27772 15851 27776
rect 15787 27716 15791 27772
rect 15791 27716 15847 27772
rect 15847 27716 15851 27772
rect 15787 27712 15851 27716
rect 15867 27772 15931 27776
rect 15867 27716 15871 27772
rect 15871 27716 15927 27772
rect 15927 27716 15931 27772
rect 15867 27712 15931 27716
rect 15947 27772 16011 27776
rect 15947 27716 15951 27772
rect 15951 27716 16007 27772
rect 16007 27716 16011 27772
rect 15947 27712 16011 27716
rect 16027 27772 16091 27776
rect 16027 27716 16031 27772
rect 16031 27716 16087 27772
rect 16087 27716 16091 27772
rect 16027 27712 16091 27716
rect 21721 27772 21785 27776
rect 21721 27716 21725 27772
rect 21725 27716 21781 27772
rect 21781 27716 21785 27772
rect 21721 27712 21785 27716
rect 21801 27772 21865 27776
rect 21801 27716 21805 27772
rect 21805 27716 21861 27772
rect 21861 27716 21865 27772
rect 21801 27712 21865 27716
rect 21881 27772 21945 27776
rect 21881 27716 21885 27772
rect 21885 27716 21941 27772
rect 21941 27716 21945 27772
rect 21881 27712 21945 27716
rect 21961 27772 22025 27776
rect 21961 27716 21965 27772
rect 21965 27716 22021 27772
rect 22021 27716 22025 27772
rect 21961 27712 22025 27716
rect 17540 27644 17604 27708
rect 7420 27236 7484 27300
rect 15332 27372 15396 27436
rect 16436 27296 16500 27300
rect 16436 27240 16486 27296
rect 16486 27240 16500 27296
rect 16436 27236 16500 27240
rect 6886 27228 6950 27232
rect 6886 27172 6890 27228
rect 6890 27172 6946 27228
rect 6946 27172 6950 27228
rect 6886 27168 6950 27172
rect 6966 27228 7030 27232
rect 6966 27172 6970 27228
rect 6970 27172 7026 27228
rect 7026 27172 7030 27228
rect 6966 27168 7030 27172
rect 7046 27228 7110 27232
rect 7046 27172 7050 27228
rect 7050 27172 7106 27228
rect 7106 27172 7110 27228
rect 7046 27168 7110 27172
rect 7126 27228 7190 27232
rect 7126 27172 7130 27228
rect 7130 27172 7186 27228
rect 7186 27172 7190 27228
rect 7126 27168 7190 27172
rect 12820 27228 12884 27232
rect 12820 27172 12824 27228
rect 12824 27172 12880 27228
rect 12880 27172 12884 27228
rect 12820 27168 12884 27172
rect 12900 27228 12964 27232
rect 12900 27172 12904 27228
rect 12904 27172 12960 27228
rect 12960 27172 12964 27228
rect 12900 27168 12964 27172
rect 12980 27228 13044 27232
rect 12980 27172 12984 27228
rect 12984 27172 13040 27228
rect 13040 27172 13044 27228
rect 12980 27168 13044 27172
rect 13060 27228 13124 27232
rect 13060 27172 13064 27228
rect 13064 27172 13120 27228
rect 13120 27172 13124 27228
rect 13060 27168 13124 27172
rect 18754 27228 18818 27232
rect 18754 27172 18758 27228
rect 18758 27172 18814 27228
rect 18814 27172 18818 27228
rect 18754 27168 18818 27172
rect 18834 27228 18898 27232
rect 18834 27172 18838 27228
rect 18838 27172 18894 27228
rect 18894 27172 18898 27228
rect 18834 27168 18898 27172
rect 18914 27228 18978 27232
rect 18914 27172 18918 27228
rect 18918 27172 18974 27228
rect 18974 27172 18978 27228
rect 18914 27168 18978 27172
rect 18994 27228 19058 27232
rect 18994 27172 18998 27228
rect 18998 27172 19054 27228
rect 19054 27172 19058 27228
rect 18994 27168 19058 27172
rect 24688 27228 24752 27232
rect 24688 27172 24692 27228
rect 24692 27172 24748 27228
rect 24748 27172 24752 27228
rect 24688 27168 24752 27172
rect 24768 27228 24832 27232
rect 24768 27172 24772 27228
rect 24772 27172 24828 27228
rect 24828 27172 24832 27228
rect 24768 27168 24832 27172
rect 24848 27228 24912 27232
rect 24848 27172 24852 27228
rect 24852 27172 24908 27228
rect 24908 27172 24912 27228
rect 24848 27168 24912 27172
rect 24928 27228 24992 27232
rect 24928 27172 24932 27228
rect 24932 27172 24988 27228
rect 24988 27172 24992 27228
rect 24928 27168 24992 27172
rect 6132 26964 6196 27028
rect 11100 26964 11164 27028
rect 21220 27024 21284 27028
rect 21220 26968 21270 27024
rect 21270 26968 21284 27024
rect 21220 26964 21284 26968
rect 15516 26828 15580 26892
rect 20300 26828 20364 26892
rect 17356 26752 17420 26756
rect 17356 26696 17370 26752
rect 17370 26696 17420 26752
rect 17356 26692 17420 26696
rect 3919 26684 3983 26688
rect 3919 26628 3923 26684
rect 3923 26628 3979 26684
rect 3979 26628 3983 26684
rect 3919 26624 3983 26628
rect 3999 26684 4063 26688
rect 3999 26628 4003 26684
rect 4003 26628 4059 26684
rect 4059 26628 4063 26684
rect 3999 26624 4063 26628
rect 4079 26684 4143 26688
rect 4079 26628 4083 26684
rect 4083 26628 4139 26684
rect 4139 26628 4143 26684
rect 4079 26624 4143 26628
rect 4159 26684 4223 26688
rect 4159 26628 4163 26684
rect 4163 26628 4219 26684
rect 4219 26628 4223 26684
rect 4159 26624 4223 26628
rect 9853 26684 9917 26688
rect 9853 26628 9857 26684
rect 9857 26628 9913 26684
rect 9913 26628 9917 26684
rect 9853 26624 9917 26628
rect 9933 26684 9997 26688
rect 9933 26628 9937 26684
rect 9937 26628 9993 26684
rect 9993 26628 9997 26684
rect 9933 26624 9997 26628
rect 10013 26684 10077 26688
rect 10013 26628 10017 26684
rect 10017 26628 10073 26684
rect 10073 26628 10077 26684
rect 10013 26624 10077 26628
rect 10093 26684 10157 26688
rect 10093 26628 10097 26684
rect 10097 26628 10153 26684
rect 10153 26628 10157 26684
rect 10093 26624 10157 26628
rect 15787 26684 15851 26688
rect 15787 26628 15791 26684
rect 15791 26628 15847 26684
rect 15847 26628 15851 26684
rect 15787 26624 15851 26628
rect 15867 26684 15931 26688
rect 15867 26628 15871 26684
rect 15871 26628 15927 26684
rect 15927 26628 15931 26684
rect 15867 26624 15931 26628
rect 15947 26684 16011 26688
rect 15947 26628 15951 26684
rect 15951 26628 16007 26684
rect 16007 26628 16011 26684
rect 15947 26624 16011 26628
rect 16027 26684 16091 26688
rect 16027 26628 16031 26684
rect 16031 26628 16087 26684
rect 16087 26628 16091 26684
rect 16027 26624 16091 26628
rect 21721 26684 21785 26688
rect 21721 26628 21725 26684
rect 21725 26628 21781 26684
rect 21781 26628 21785 26684
rect 21721 26624 21785 26628
rect 21801 26684 21865 26688
rect 21801 26628 21805 26684
rect 21805 26628 21861 26684
rect 21861 26628 21865 26684
rect 21801 26624 21865 26628
rect 21881 26684 21945 26688
rect 21881 26628 21885 26684
rect 21885 26628 21941 26684
rect 21941 26628 21945 26684
rect 21881 26624 21945 26628
rect 21961 26684 22025 26688
rect 21961 26628 21965 26684
rect 21965 26628 22021 26684
rect 22021 26628 22025 26684
rect 21961 26624 22025 26628
rect 1900 26284 1964 26348
rect 11652 26208 11716 26212
rect 11652 26152 11702 26208
rect 11702 26152 11716 26208
rect 11652 26148 11716 26152
rect 6886 26140 6950 26144
rect 6886 26084 6890 26140
rect 6890 26084 6946 26140
rect 6946 26084 6950 26140
rect 6886 26080 6950 26084
rect 6966 26140 7030 26144
rect 6966 26084 6970 26140
rect 6970 26084 7026 26140
rect 7026 26084 7030 26140
rect 6966 26080 7030 26084
rect 7046 26140 7110 26144
rect 7046 26084 7050 26140
rect 7050 26084 7106 26140
rect 7106 26084 7110 26140
rect 7046 26080 7110 26084
rect 7126 26140 7190 26144
rect 7126 26084 7130 26140
rect 7130 26084 7186 26140
rect 7186 26084 7190 26140
rect 7126 26080 7190 26084
rect 12820 26140 12884 26144
rect 12820 26084 12824 26140
rect 12824 26084 12880 26140
rect 12880 26084 12884 26140
rect 12820 26080 12884 26084
rect 12900 26140 12964 26144
rect 12900 26084 12904 26140
rect 12904 26084 12960 26140
rect 12960 26084 12964 26140
rect 12900 26080 12964 26084
rect 12980 26140 13044 26144
rect 12980 26084 12984 26140
rect 12984 26084 13040 26140
rect 13040 26084 13044 26140
rect 12980 26080 13044 26084
rect 13060 26140 13124 26144
rect 13060 26084 13064 26140
rect 13064 26084 13120 26140
rect 13120 26084 13124 26140
rect 13060 26080 13124 26084
rect 18754 26140 18818 26144
rect 18754 26084 18758 26140
rect 18758 26084 18814 26140
rect 18814 26084 18818 26140
rect 18754 26080 18818 26084
rect 18834 26140 18898 26144
rect 18834 26084 18838 26140
rect 18838 26084 18894 26140
rect 18894 26084 18898 26140
rect 18834 26080 18898 26084
rect 18914 26140 18978 26144
rect 18914 26084 18918 26140
rect 18918 26084 18974 26140
rect 18974 26084 18978 26140
rect 18914 26080 18978 26084
rect 18994 26140 19058 26144
rect 18994 26084 18998 26140
rect 18998 26084 19054 26140
rect 19054 26084 19058 26140
rect 18994 26080 19058 26084
rect 24688 26140 24752 26144
rect 24688 26084 24692 26140
rect 24692 26084 24748 26140
rect 24748 26084 24752 26140
rect 24688 26080 24752 26084
rect 24768 26140 24832 26144
rect 24768 26084 24772 26140
rect 24772 26084 24828 26140
rect 24828 26084 24832 26140
rect 24768 26080 24832 26084
rect 24848 26140 24912 26144
rect 24848 26084 24852 26140
rect 24852 26084 24908 26140
rect 24908 26084 24912 26140
rect 24848 26080 24912 26084
rect 24928 26140 24992 26144
rect 24928 26084 24932 26140
rect 24932 26084 24988 26140
rect 24988 26084 24992 26140
rect 24928 26080 24992 26084
rect 2268 26012 2332 26076
rect 12020 26012 12084 26076
rect 16252 25876 16316 25940
rect 8340 25740 8404 25804
rect 17172 25604 17236 25668
rect 3919 25596 3983 25600
rect 3919 25540 3923 25596
rect 3923 25540 3979 25596
rect 3979 25540 3983 25596
rect 3919 25536 3983 25540
rect 3999 25596 4063 25600
rect 3999 25540 4003 25596
rect 4003 25540 4059 25596
rect 4059 25540 4063 25596
rect 3999 25536 4063 25540
rect 4079 25596 4143 25600
rect 4079 25540 4083 25596
rect 4083 25540 4139 25596
rect 4139 25540 4143 25596
rect 4079 25536 4143 25540
rect 4159 25596 4223 25600
rect 4159 25540 4163 25596
rect 4163 25540 4219 25596
rect 4219 25540 4223 25596
rect 4159 25536 4223 25540
rect 9853 25596 9917 25600
rect 9853 25540 9857 25596
rect 9857 25540 9913 25596
rect 9913 25540 9917 25596
rect 9853 25536 9917 25540
rect 9933 25596 9997 25600
rect 9933 25540 9937 25596
rect 9937 25540 9993 25596
rect 9993 25540 9997 25596
rect 9933 25536 9997 25540
rect 10013 25596 10077 25600
rect 10013 25540 10017 25596
rect 10017 25540 10073 25596
rect 10073 25540 10077 25596
rect 10013 25536 10077 25540
rect 10093 25596 10157 25600
rect 10093 25540 10097 25596
rect 10097 25540 10153 25596
rect 10153 25540 10157 25596
rect 10093 25536 10157 25540
rect 15787 25596 15851 25600
rect 15787 25540 15791 25596
rect 15791 25540 15847 25596
rect 15847 25540 15851 25596
rect 15787 25536 15851 25540
rect 15867 25596 15931 25600
rect 15867 25540 15871 25596
rect 15871 25540 15927 25596
rect 15927 25540 15931 25596
rect 15867 25536 15931 25540
rect 15947 25596 16011 25600
rect 15947 25540 15951 25596
rect 15951 25540 16007 25596
rect 16007 25540 16011 25596
rect 15947 25536 16011 25540
rect 16027 25596 16091 25600
rect 16027 25540 16031 25596
rect 16031 25540 16087 25596
rect 16087 25540 16091 25596
rect 16027 25536 16091 25540
rect 21721 25596 21785 25600
rect 21721 25540 21725 25596
rect 21725 25540 21781 25596
rect 21781 25540 21785 25596
rect 21721 25536 21785 25540
rect 21801 25596 21865 25600
rect 21801 25540 21805 25596
rect 21805 25540 21861 25596
rect 21861 25540 21865 25596
rect 21801 25536 21865 25540
rect 21881 25596 21945 25600
rect 21881 25540 21885 25596
rect 21885 25540 21941 25596
rect 21941 25540 21945 25596
rect 21881 25536 21945 25540
rect 21961 25596 22025 25600
rect 21961 25540 21965 25596
rect 21965 25540 22021 25596
rect 22021 25540 22025 25596
rect 21961 25536 22025 25540
rect 2636 25528 2700 25532
rect 2636 25472 2686 25528
rect 2686 25472 2700 25528
rect 2636 25468 2700 25472
rect 17540 25256 17604 25260
rect 17540 25200 17590 25256
rect 17590 25200 17604 25256
rect 17540 25196 17604 25200
rect 12204 25060 12268 25124
rect 14228 25060 14292 25124
rect 6886 25052 6950 25056
rect 6886 24996 6890 25052
rect 6890 24996 6946 25052
rect 6946 24996 6950 25052
rect 6886 24992 6950 24996
rect 6966 25052 7030 25056
rect 6966 24996 6970 25052
rect 6970 24996 7026 25052
rect 7026 24996 7030 25052
rect 6966 24992 7030 24996
rect 7046 25052 7110 25056
rect 7046 24996 7050 25052
rect 7050 24996 7106 25052
rect 7106 24996 7110 25052
rect 7046 24992 7110 24996
rect 7126 25052 7190 25056
rect 7126 24996 7130 25052
rect 7130 24996 7186 25052
rect 7186 24996 7190 25052
rect 7126 24992 7190 24996
rect 12820 25052 12884 25056
rect 12820 24996 12824 25052
rect 12824 24996 12880 25052
rect 12880 24996 12884 25052
rect 12820 24992 12884 24996
rect 12900 25052 12964 25056
rect 12900 24996 12904 25052
rect 12904 24996 12960 25052
rect 12960 24996 12964 25052
rect 12900 24992 12964 24996
rect 12980 25052 13044 25056
rect 12980 24996 12984 25052
rect 12984 24996 13040 25052
rect 13040 24996 13044 25052
rect 12980 24992 13044 24996
rect 13060 25052 13124 25056
rect 13060 24996 13064 25052
rect 13064 24996 13120 25052
rect 13120 24996 13124 25052
rect 13060 24992 13124 24996
rect 3740 24924 3804 24988
rect 18754 25052 18818 25056
rect 18754 24996 18758 25052
rect 18758 24996 18814 25052
rect 18814 24996 18818 25052
rect 18754 24992 18818 24996
rect 18834 25052 18898 25056
rect 18834 24996 18838 25052
rect 18838 24996 18894 25052
rect 18894 24996 18898 25052
rect 18834 24992 18898 24996
rect 18914 25052 18978 25056
rect 18914 24996 18918 25052
rect 18918 24996 18974 25052
rect 18974 24996 18978 25052
rect 18914 24992 18978 24996
rect 18994 25052 19058 25056
rect 18994 24996 18998 25052
rect 18998 24996 19054 25052
rect 19054 24996 19058 25052
rect 18994 24992 19058 24996
rect 24688 25052 24752 25056
rect 24688 24996 24692 25052
rect 24692 24996 24748 25052
rect 24748 24996 24752 25052
rect 24688 24992 24752 24996
rect 24768 25052 24832 25056
rect 24768 24996 24772 25052
rect 24772 24996 24828 25052
rect 24828 24996 24832 25052
rect 24768 24992 24832 24996
rect 24848 25052 24912 25056
rect 24848 24996 24852 25052
rect 24852 24996 24908 25052
rect 24908 24996 24912 25052
rect 24848 24992 24912 24996
rect 24928 25052 24992 25056
rect 24928 24996 24932 25052
rect 24932 24996 24988 25052
rect 24988 24996 24992 25052
rect 24928 24992 24992 24996
rect 16620 24924 16684 24988
rect 2636 24788 2700 24852
rect 22508 24788 22572 24852
rect 4292 24652 4356 24716
rect 15332 24516 15396 24580
rect 19932 24516 19996 24580
rect 3919 24508 3983 24512
rect 3919 24452 3923 24508
rect 3923 24452 3979 24508
rect 3979 24452 3983 24508
rect 3919 24448 3983 24452
rect 3999 24508 4063 24512
rect 3999 24452 4003 24508
rect 4003 24452 4059 24508
rect 4059 24452 4063 24508
rect 3999 24448 4063 24452
rect 4079 24508 4143 24512
rect 4079 24452 4083 24508
rect 4083 24452 4139 24508
rect 4139 24452 4143 24508
rect 4079 24448 4143 24452
rect 4159 24508 4223 24512
rect 4159 24452 4163 24508
rect 4163 24452 4219 24508
rect 4219 24452 4223 24508
rect 4159 24448 4223 24452
rect 9853 24508 9917 24512
rect 9853 24452 9857 24508
rect 9857 24452 9913 24508
rect 9913 24452 9917 24508
rect 9853 24448 9917 24452
rect 9933 24508 9997 24512
rect 9933 24452 9937 24508
rect 9937 24452 9993 24508
rect 9993 24452 9997 24508
rect 9933 24448 9997 24452
rect 10013 24508 10077 24512
rect 10013 24452 10017 24508
rect 10017 24452 10073 24508
rect 10073 24452 10077 24508
rect 10013 24448 10077 24452
rect 10093 24508 10157 24512
rect 10093 24452 10097 24508
rect 10097 24452 10153 24508
rect 10153 24452 10157 24508
rect 10093 24448 10157 24452
rect 15787 24508 15851 24512
rect 15787 24452 15791 24508
rect 15791 24452 15847 24508
rect 15847 24452 15851 24508
rect 15787 24448 15851 24452
rect 15867 24508 15931 24512
rect 15867 24452 15871 24508
rect 15871 24452 15927 24508
rect 15927 24452 15931 24508
rect 15867 24448 15931 24452
rect 15947 24508 16011 24512
rect 15947 24452 15951 24508
rect 15951 24452 16007 24508
rect 16007 24452 16011 24508
rect 15947 24448 16011 24452
rect 16027 24508 16091 24512
rect 16027 24452 16031 24508
rect 16031 24452 16087 24508
rect 16087 24452 16091 24508
rect 16027 24448 16091 24452
rect 21721 24508 21785 24512
rect 21721 24452 21725 24508
rect 21725 24452 21781 24508
rect 21781 24452 21785 24508
rect 21721 24448 21785 24452
rect 21801 24508 21865 24512
rect 21801 24452 21805 24508
rect 21805 24452 21861 24508
rect 21861 24452 21865 24508
rect 21801 24448 21865 24452
rect 21881 24508 21945 24512
rect 21881 24452 21885 24508
rect 21885 24452 21941 24508
rect 21941 24452 21945 24508
rect 21881 24448 21945 24452
rect 21961 24508 22025 24512
rect 21961 24452 21965 24508
rect 21965 24452 22021 24508
rect 22021 24452 22025 24508
rect 21961 24448 22025 24452
rect 4476 24244 4540 24308
rect 6132 23972 6196 24036
rect 16436 24244 16500 24308
rect 22876 24244 22940 24308
rect 17724 24108 17788 24172
rect 6886 23964 6950 23968
rect 6886 23908 6890 23964
rect 6890 23908 6946 23964
rect 6946 23908 6950 23964
rect 6886 23904 6950 23908
rect 6966 23964 7030 23968
rect 6966 23908 6970 23964
rect 6970 23908 7026 23964
rect 7026 23908 7030 23964
rect 6966 23904 7030 23908
rect 7046 23964 7110 23968
rect 7046 23908 7050 23964
rect 7050 23908 7106 23964
rect 7106 23908 7110 23964
rect 7046 23904 7110 23908
rect 7126 23964 7190 23968
rect 7126 23908 7130 23964
rect 7130 23908 7186 23964
rect 7186 23908 7190 23964
rect 7126 23904 7190 23908
rect 12820 23964 12884 23968
rect 12820 23908 12824 23964
rect 12824 23908 12880 23964
rect 12880 23908 12884 23964
rect 12820 23904 12884 23908
rect 12900 23964 12964 23968
rect 12900 23908 12904 23964
rect 12904 23908 12960 23964
rect 12960 23908 12964 23964
rect 12900 23904 12964 23908
rect 12980 23964 13044 23968
rect 12980 23908 12984 23964
rect 12984 23908 13040 23964
rect 13040 23908 13044 23964
rect 12980 23904 13044 23908
rect 13060 23964 13124 23968
rect 13060 23908 13064 23964
rect 13064 23908 13120 23964
rect 13120 23908 13124 23964
rect 13060 23904 13124 23908
rect 18754 23964 18818 23968
rect 18754 23908 18758 23964
rect 18758 23908 18814 23964
rect 18814 23908 18818 23964
rect 18754 23904 18818 23908
rect 18834 23964 18898 23968
rect 18834 23908 18838 23964
rect 18838 23908 18894 23964
rect 18894 23908 18898 23964
rect 18834 23904 18898 23908
rect 18914 23964 18978 23968
rect 18914 23908 18918 23964
rect 18918 23908 18974 23964
rect 18974 23908 18978 23964
rect 18914 23904 18978 23908
rect 18994 23964 19058 23968
rect 18994 23908 18998 23964
rect 18998 23908 19054 23964
rect 19054 23908 19058 23964
rect 18994 23904 19058 23908
rect 24688 23964 24752 23968
rect 24688 23908 24692 23964
rect 24692 23908 24748 23964
rect 24748 23908 24752 23964
rect 24688 23904 24752 23908
rect 24768 23964 24832 23968
rect 24768 23908 24772 23964
rect 24772 23908 24828 23964
rect 24828 23908 24832 23964
rect 24768 23904 24832 23908
rect 24848 23964 24912 23968
rect 24848 23908 24852 23964
rect 24852 23908 24908 23964
rect 24908 23908 24912 23964
rect 24848 23904 24912 23908
rect 24928 23964 24992 23968
rect 24928 23908 24932 23964
rect 24932 23908 24988 23964
rect 24988 23908 24992 23964
rect 24928 23904 24992 23908
rect 10732 23836 10796 23900
rect 7420 23564 7484 23628
rect 22692 23564 22756 23628
rect 22692 23428 22756 23492
rect 3919 23420 3983 23424
rect 3919 23364 3923 23420
rect 3923 23364 3979 23420
rect 3979 23364 3983 23420
rect 3919 23360 3983 23364
rect 3999 23420 4063 23424
rect 3999 23364 4003 23420
rect 4003 23364 4059 23420
rect 4059 23364 4063 23420
rect 3999 23360 4063 23364
rect 4079 23420 4143 23424
rect 4079 23364 4083 23420
rect 4083 23364 4139 23420
rect 4139 23364 4143 23420
rect 4079 23360 4143 23364
rect 4159 23420 4223 23424
rect 4159 23364 4163 23420
rect 4163 23364 4219 23420
rect 4219 23364 4223 23420
rect 4159 23360 4223 23364
rect 9853 23420 9917 23424
rect 9853 23364 9857 23420
rect 9857 23364 9913 23420
rect 9913 23364 9917 23420
rect 9853 23360 9917 23364
rect 9933 23420 9997 23424
rect 9933 23364 9937 23420
rect 9937 23364 9993 23420
rect 9993 23364 9997 23420
rect 9933 23360 9997 23364
rect 10013 23420 10077 23424
rect 10013 23364 10017 23420
rect 10017 23364 10073 23420
rect 10073 23364 10077 23420
rect 10013 23360 10077 23364
rect 10093 23420 10157 23424
rect 10093 23364 10097 23420
rect 10097 23364 10153 23420
rect 10153 23364 10157 23420
rect 10093 23360 10157 23364
rect 15787 23420 15851 23424
rect 15787 23364 15791 23420
rect 15791 23364 15847 23420
rect 15847 23364 15851 23420
rect 15787 23360 15851 23364
rect 15867 23420 15931 23424
rect 15867 23364 15871 23420
rect 15871 23364 15927 23420
rect 15927 23364 15931 23420
rect 15867 23360 15931 23364
rect 15947 23420 16011 23424
rect 15947 23364 15951 23420
rect 15951 23364 16007 23420
rect 16007 23364 16011 23420
rect 15947 23360 16011 23364
rect 16027 23420 16091 23424
rect 16027 23364 16031 23420
rect 16031 23364 16087 23420
rect 16087 23364 16091 23420
rect 16027 23360 16091 23364
rect 21721 23420 21785 23424
rect 21721 23364 21725 23420
rect 21725 23364 21781 23420
rect 21781 23364 21785 23420
rect 21721 23360 21785 23364
rect 21801 23420 21865 23424
rect 21801 23364 21805 23420
rect 21805 23364 21861 23420
rect 21861 23364 21865 23420
rect 21801 23360 21865 23364
rect 21881 23420 21945 23424
rect 21881 23364 21885 23420
rect 21885 23364 21941 23420
rect 21941 23364 21945 23420
rect 21881 23360 21945 23364
rect 21961 23420 22025 23424
rect 21961 23364 21965 23420
rect 21965 23364 22021 23420
rect 22021 23364 22025 23420
rect 21961 23360 22025 23364
rect 3372 23156 3436 23220
rect 5580 23156 5644 23220
rect 2268 22884 2332 22948
rect 6886 22876 6950 22880
rect 6886 22820 6890 22876
rect 6890 22820 6946 22876
rect 6946 22820 6950 22876
rect 6886 22816 6950 22820
rect 6966 22876 7030 22880
rect 6966 22820 6970 22876
rect 6970 22820 7026 22876
rect 7026 22820 7030 22876
rect 6966 22816 7030 22820
rect 7046 22876 7110 22880
rect 7046 22820 7050 22876
rect 7050 22820 7106 22876
rect 7106 22820 7110 22876
rect 7046 22816 7110 22820
rect 7126 22876 7190 22880
rect 7126 22820 7130 22876
rect 7130 22820 7186 22876
rect 7186 22820 7190 22876
rect 7126 22816 7190 22820
rect 12820 22876 12884 22880
rect 12820 22820 12824 22876
rect 12824 22820 12880 22876
rect 12880 22820 12884 22876
rect 12820 22816 12884 22820
rect 12900 22876 12964 22880
rect 12900 22820 12904 22876
rect 12904 22820 12960 22876
rect 12960 22820 12964 22876
rect 12900 22816 12964 22820
rect 12980 22876 13044 22880
rect 12980 22820 12984 22876
rect 12984 22820 13040 22876
rect 13040 22820 13044 22876
rect 12980 22816 13044 22820
rect 13060 22876 13124 22880
rect 13060 22820 13064 22876
rect 13064 22820 13120 22876
rect 13120 22820 13124 22876
rect 13060 22816 13124 22820
rect 18754 22876 18818 22880
rect 18754 22820 18758 22876
rect 18758 22820 18814 22876
rect 18814 22820 18818 22876
rect 18754 22816 18818 22820
rect 18834 22876 18898 22880
rect 18834 22820 18838 22876
rect 18838 22820 18894 22876
rect 18894 22820 18898 22876
rect 18834 22816 18898 22820
rect 18914 22876 18978 22880
rect 18914 22820 18918 22876
rect 18918 22820 18974 22876
rect 18974 22820 18978 22876
rect 18914 22816 18978 22820
rect 18994 22876 19058 22880
rect 18994 22820 18998 22876
rect 18998 22820 19054 22876
rect 19054 22820 19058 22876
rect 18994 22816 19058 22820
rect 24688 22876 24752 22880
rect 24688 22820 24692 22876
rect 24692 22820 24748 22876
rect 24748 22820 24752 22876
rect 24688 22816 24752 22820
rect 24768 22876 24832 22880
rect 24768 22820 24772 22876
rect 24772 22820 24828 22876
rect 24828 22820 24832 22876
rect 24768 22816 24832 22820
rect 24848 22876 24912 22880
rect 24848 22820 24852 22876
rect 24852 22820 24908 22876
rect 24908 22820 24912 22876
rect 24848 22816 24912 22820
rect 24928 22876 24992 22880
rect 24928 22820 24932 22876
rect 24932 22820 24988 22876
rect 24988 22820 24992 22876
rect 24928 22816 24992 22820
rect 5396 22748 5460 22812
rect 11468 22476 11532 22540
rect 3919 22332 3983 22336
rect 3919 22276 3923 22332
rect 3923 22276 3979 22332
rect 3979 22276 3983 22332
rect 3919 22272 3983 22276
rect 3999 22332 4063 22336
rect 3999 22276 4003 22332
rect 4003 22276 4059 22332
rect 4059 22276 4063 22332
rect 3999 22272 4063 22276
rect 4079 22332 4143 22336
rect 4079 22276 4083 22332
rect 4083 22276 4139 22332
rect 4139 22276 4143 22332
rect 4079 22272 4143 22276
rect 4159 22332 4223 22336
rect 4159 22276 4163 22332
rect 4163 22276 4219 22332
rect 4219 22276 4223 22332
rect 4159 22272 4223 22276
rect 9853 22332 9917 22336
rect 9853 22276 9857 22332
rect 9857 22276 9913 22332
rect 9913 22276 9917 22332
rect 9853 22272 9917 22276
rect 9933 22332 9997 22336
rect 9933 22276 9937 22332
rect 9937 22276 9993 22332
rect 9993 22276 9997 22332
rect 9933 22272 9997 22276
rect 10013 22332 10077 22336
rect 10013 22276 10017 22332
rect 10017 22276 10073 22332
rect 10073 22276 10077 22332
rect 10013 22272 10077 22276
rect 10093 22332 10157 22336
rect 10093 22276 10097 22332
rect 10097 22276 10153 22332
rect 10153 22276 10157 22332
rect 10093 22272 10157 22276
rect 15787 22332 15851 22336
rect 15787 22276 15791 22332
rect 15791 22276 15847 22332
rect 15847 22276 15851 22332
rect 15787 22272 15851 22276
rect 15867 22332 15931 22336
rect 15867 22276 15871 22332
rect 15871 22276 15927 22332
rect 15927 22276 15931 22332
rect 15867 22272 15931 22276
rect 15947 22332 16011 22336
rect 15947 22276 15951 22332
rect 15951 22276 16007 22332
rect 16007 22276 16011 22332
rect 15947 22272 16011 22276
rect 16027 22332 16091 22336
rect 16027 22276 16031 22332
rect 16031 22276 16087 22332
rect 16087 22276 16091 22332
rect 16027 22272 16091 22276
rect 21721 22332 21785 22336
rect 21721 22276 21725 22332
rect 21725 22276 21781 22332
rect 21781 22276 21785 22332
rect 21721 22272 21785 22276
rect 21801 22332 21865 22336
rect 21801 22276 21805 22332
rect 21805 22276 21861 22332
rect 21861 22276 21865 22332
rect 21801 22272 21865 22276
rect 21881 22332 21945 22336
rect 21881 22276 21885 22332
rect 21885 22276 21941 22332
rect 21941 22276 21945 22332
rect 21881 22272 21945 22276
rect 21961 22332 22025 22336
rect 21961 22276 21965 22332
rect 21965 22276 22021 22332
rect 22021 22276 22025 22332
rect 21961 22272 22025 22276
rect 13860 21932 13924 21996
rect 17172 21796 17236 21860
rect 6886 21788 6950 21792
rect 6886 21732 6890 21788
rect 6890 21732 6946 21788
rect 6946 21732 6950 21788
rect 6886 21728 6950 21732
rect 6966 21788 7030 21792
rect 6966 21732 6970 21788
rect 6970 21732 7026 21788
rect 7026 21732 7030 21788
rect 6966 21728 7030 21732
rect 7046 21788 7110 21792
rect 7046 21732 7050 21788
rect 7050 21732 7106 21788
rect 7106 21732 7110 21788
rect 7046 21728 7110 21732
rect 7126 21788 7190 21792
rect 7126 21732 7130 21788
rect 7130 21732 7186 21788
rect 7186 21732 7190 21788
rect 7126 21728 7190 21732
rect 12820 21788 12884 21792
rect 12820 21732 12824 21788
rect 12824 21732 12880 21788
rect 12880 21732 12884 21788
rect 12820 21728 12884 21732
rect 12900 21788 12964 21792
rect 12900 21732 12904 21788
rect 12904 21732 12960 21788
rect 12960 21732 12964 21788
rect 12900 21728 12964 21732
rect 12980 21788 13044 21792
rect 12980 21732 12984 21788
rect 12984 21732 13040 21788
rect 13040 21732 13044 21788
rect 12980 21728 13044 21732
rect 13060 21788 13124 21792
rect 13060 21732 13064 21788
rect 13064 21732 13120 21788
rect 13120 21732 13124 21788
rect 13060 21728 13124 21732
rect 18754 21788 18818 21792
rect 18754 21732 18758 21788
rect 18758 21732 18814 21788
rect 18814 21732 18818 21788
rect 18754 21728 18818 21732
rect 18834 21788 18898 21792
rect 18834 21732 18838 21788
rect 18838 21732 18894 21788
rect 18894 21732 18898 21788
rect 18834 21728 18898 21732
rect 18914 21788 18978 21792
rect 18914 21732 18918 21788
rect 18918 21732 18974 21788
rect 18974 21732 18978 21788
rect 18914 21728 18978 21732
rect 18994 21788 19058 21792
rect 18994 21732 18998 21788
rect 18998 21732 19054 21788
rect 19054 21732 19058 21788
rect 18994 21728 19058 21732
rect 24688 21788 24752 21792
rect 24688 21732 24692 21788
rect 24692 21732 24748 21788
rect 24748 21732 24752 21788
rect 24688 21728 24752 21732
rect 24768 21788 24832 21792
rect 24768 21732 24772 21788
rect 24772 21732 24828 21788
rect 24828 21732 24832 21788
rect 24768 21728 24832 21732
rect 24848 21788 24912 21792
rect 24848 21732 24852 21788
rect 24852 21732 24908 21788
rect 24908 21732 24912 21788
rect 24848 21728 24912 21732
rect 24928 21788 24992 21792
rect 24928 21732 24932 21788
rect 24932 21732 24988 21788
rect 24988 21732 24992 21788
rect 24928 21728 24992 21732
rect 5028 21388 5092 21452
rect 17540 21524 17604 21588
rect 9260 21252 9324 21316
rect 16620 21388 16684 21452
rect 3919 21244 3983 21248
rect 3919 21188 3923 21244
rect 3923 21188 3979 21244
rect 3979 21188 3983 21244
rect 3919 21184 3983 21188
rect 3999 21244 4063 21248
rect 3999 21188 4003 21244
rect 4003 21188 4059 21244
rect 4059 21188 4063 21244
rect 3999 21184 4063 21188
rect 4079 21244 4143 21248
rect 4079 21188 4083 21244
rect 4083 21188 4139 21244
rect 4139 21188 4143 21244
rect 4079 21184 4143 21188
rect 4159 21244 4223 21248
rect 4159 21188 4163 21244
rect 4163 21188 4219 21244
rect 4219 21188 4223 21244
rect 4159 21184 4223 21188
rect 9853 21244 9917 21248
rect 9853 21188 9857 21244
rect 9857 21188 9913 21244
rect 9913 21188 9917 21244
rect 9853 21184 9917 21188
rect 9933 21244 9997 21248
rect 9933 21188 9937 21244
rect 9937 21188 9993 21244
rect 9993 21188 9997 21244
rect 9933 21184 9997 21188
rect 10013 21244 10077 21248
rect 10013 21188 10017 21244
rect 10017 21188 10073 21244
rect 10073 21188 10077 21244
rect 10013 21184 10077 21188
rect 10093 21244 10157 21248
rect 10093 21188 10097 21244
rect 10097 21188 10153 21244
rect 10153 21188 10157 21244
rect 10093 21184 10157 21188
rect 16436 21252 16500 21316
rect 15787 21244 15851 21248
rect 15787 21188 15791 21244
rect 15791 21188 15847 21244
rect 15847 21188 15851 21244
rect 15787 21184 15851 21188
rect 15867 21244 15931 21248
rect 15867 21188 15871 21244
rect 15871 21188 15927 21244
rect 15927 21188 15931 21244
rect 15867 21184 15931 21188
rect 15947 21244 16011 21248
rect 15947 21188 15951 21244
rect 15951 21188 16007 21244
rect 16007 21188 16011 21244
rect 15947 21184 16011 21188
rect 16027 21244 16091 21248
rect 16027 21188 16031 21244
rect 16031 21188 16087 21244
rect 16087 21188 16091 21244
rect 16027 21184 16091 21188
rect 21721 21244 21785 21248
rect 21721 21188 21725 21244
rect 21725 21188 21781 21244
rect 21781 21188 21785 21244
rect 21721 21184 21785 21188
rect 21801 21244 21865 21248
rect 21801 21188 21805 21244
rect 21805 21188 21861 21244
rect 21861 21188 21865 21244
rect 21801 21184 21865 21188
rect 21881 21244 21945 21248
rect 21881 21188 21885 21244
rect 21885 21188 21941 21244
rect 21941 21188 21945 21244
rect 21881 21184 21945 21188
rect 21961 21244 22025 21248
rect 21961 21188 21965 21244
rect 21965 21188 22021 21244
rect 22021 21188 22025 21244
rect 21961 21184 22025 21188
rect 17356 21176 17420 21180
rect 17356 21120 17370 21176
rect 17370 21120 17420 21176
rect 17356 21116 17420 21120
rect 19564 21116 19628 21180
rect 19932 21176 19996 21180
rect 19932 21120 19982 21176
rect 19982 21120 19996 21176
rect 19932 21116 19996 21120
rect 6684 20844 6748 20908
rect 9628 20844 9692 20908
rect 12572 20844 12636 20908
rect 2452 20708 2516 20772
rect 3188 20708 3252 20772
rect 6316 20708 6380 20772
rect 7604 20768 7668 20772
rect 7604 20712 7618 20768
rect 7618 20712 7668 20768
rect 7604 20708 7668 20712
rect 19380 20768 19444 20772
rect 19380 20712 19394 20768
rect 19394 20712 19444 20768
rect 19380 20708 19444 20712
rect 6886 20700 6950 20704
rect 6886 20644 6890 20700
rect 6890 20644 6946 20700
rect 6946 20644 6950 20700
rect 6886 20640 6950 20644
rect 6966 20700 7030 20704
rect 6966 20644 6970 20700
rect 6970 20644 7026 20700
rect 7026 20644 7030 20700
rect 6966 20640 7030 20644
rect 7046 20700 7110 20704
rect 7046 20644 7050 20700
rect 7050 20644 7106 20700
rect 7106 20644 7110 20700
rect 7046 20640 7110 20644
rect 7126 20700 7190 20704
rect 7126 20644 7130 20700
rect 7130 20644 7186 20700
rect 7186 20644 7190 20700
rect 7126 20640 7190 20644
rect 12820 20700 12884 20704
rect 12820 20644 12824 20700
rect 12824 20644 12880 20700
rect 12880 20644 12884 20700
rect 12820 20640 12884 20644
rect 12900 20700 12964 20704
rect 12900 20644 12904 20700
rect 12904 20644 12960 20700
rect 12960 20644 12964 20700
rect 12900 20640 12964 20644
rect 12980 20700 13044 20704
rect 12980 20644 12984 20700
rect 12984 20644 13040 20700
rect 13040 20644 13044 20700
rect 12980 20640 13044 20644
rect 13060 20700 13124 20704
rect 13060 20644 13064 20700
rect 13064 20644 13120 20700
rect 13120 20644 13124 20700
rect 13060 20640 13124 20644
rect 18754 20700 18818 20704
rect 18754 20644 18758 20700
rect 18758 20644 18814 20700
rect 18814 20644 18818 20700
rect 18754 20640 18818 20644
rect 18834 20700 18898 20704
rect 18834 20644 18838 20700
rect 18838 20644 18894 20700
rect 18894 20644 18898 20700
rect 18834 20640 18898 20644
rect 18914 20700 18978 20704
rect 18914 20644 18918 20700
rect 18918 20644 18974 20700
rect 18974 20644 18978 20700
rect 18914 20640 18978 20644
rect 18994 20700 19058 20704
rect 18994 20644 18998 20700
rect 18998 20644 19054 20700
rect 19054 20644 19058 20700
rect 18994 20640 19058 20644
rect 24688 20700 24752 20704
rect 24688 20644 24692 20700
rect 24692 20644 24748 20700
rect 24748 20644 24752 20700
rect 24688 20640 24752 20644
rect 24768 20700 24832 20704
rect 24768 20644 24772 20700
rect 24772 20644 24828 20700
rect 24828 20644 24832 20700
rect 24768 20640 24832 20644
rect 24848 20700 24912 20704
rect 24848 20644 24852 20700
rect 24852 20644 24908 20700
rect 24908 20644 24912 20700
rect 24848 20640 24912 20644
rect 24928 20700 24992 20704
rect 24928 20644 24932 20700
rect 24932 20644 24988 20700
rect 24988 20644 24992 20700
rect 24928 20640 24992 20644
rect 3740 20436 3804 20500
rect 3919 20156 3983 20160
rect 3919 20100 3923 20156
rect 3923 20100 3979 20156
rect 3979 20100 3983 20156
rect 3919 20096 3983 20100
rect 3999 20156 4063 20160
rect 3999 20100 4003 20156
rect 4003 20100 4059 20156
rect 4059 20100 4063 20156
rect 3999 20096 4063 20100
rect 4079 20156 4143 20160
rect 4079 20100 4083 20156
rect 4083 20100 4139 20156
rect 4139 20100 4143 20156
rect 4079 20096 4143 20100
rect 4159 20156 4223 20160
rect 4159 20100 4163 20156
rect 4163 20100 4219 20156
rect 4219 20100 4223 20156
rect 4159 20096 4223 20100
rect 9853 20156 9917 20160
rect 9853 20100 9857 20156
rect 9857 20100 9913 20156
rect 9913 20100 9917 20156
rect 9853 20096 9917 20100
rect 9933 20156 9997 20160
rect 9933 20100 9937 20156
rect 9937 20100 9993 20156
rect 9993 20100 9997 20156
rect 9933 20096 9997 20100
rect 10013 20156 10077 20160
rect 10013 20100 10017 20156
rect 10017 20100 10073 20156
rect 10073 20100 10077 20156
rect 10013 20096 10077 20100
rect 10093 20156 10157 20160
rect 10093 20100 10097 20156
rect 10097 20100 10153 20156
rect 10153 20100 10157 20156
rect 10093 20096 10157 20100
rect 15787 20156 15851 20160
rect 15787 20100 15791 20156
rect 15791 20100 15847 20156
rect 15847 20100 15851 20156
rect 15787 20096 15851 20100
rect 15867 20156 15931 20160
rect 15867 20100 15871 20156
rect 15871 20100 15927 20156
rect 15927 20100 15931 20156
rect 15867 20096 15931 20100
rect 15947 20156 16011 20160
rect 15947 20100 15951 20156
rect 15951 20100 16007 20156
rect 16007 20100 16011 20156
rect 15947 20096 16011 20100
rect 16027 20156 16091 20160
rect 16027 20100 16031 20156
rect 16031 20100 16087 20156
rect 16087 20100 16091 20156
rect 16027 20096 16091 20100
rect 21721 20156 21785 20160
rect 21721 20100 21725 20156
rect 21725 20100 21781 20156
rect 21781 20100 21785 20156
rect 21721 20096 21785 20100
rect 21801 20156 21865 20160
rect 21801 20100 21805 20156
rect 21805 20100 21861 20156
rect 21861 20100 21865 20156
rect 21801 20096 21865 20100
rect 21881 20156 21945 20160
rect 21881 20100 21885 20156
rect 21885 20100 21941 20156
rect 21941 20100 21945 20156
rect 21881 20096 21945 20100
rect 21961 20156 22025 20160
rect 21961 20100 21965 20156
rect 21965 20100 22021 20156
rect 22021 20100 22025 20156
rect 21961 20096 22025 20100
rect 2636 19892 2700 19956
rect 14964 19892 15028 19956
rect 8156 19756 8220 19820
rect 10732 19756 10796 19820
rect 13676 19756 13740 19820
rect 21220 19620 21284 19684
rect 6886 19612 6950 19616
rect 6886 19556 6890 19612
rect 6890 19556 6946 19612
rect 6946 19556 6950 19612
rect 6886 19552 6950 19556
rect 6966 19612 7030 19616
rect 6966 19556 6970 19612
rect 6970 19556 7026 19612
rect 7026 19556 7030 19612
rect 6966 19552 7030 19556
rect 7046 19612 7110 19616
rect 7046 19556 7050 19612
rect 7050 19556 7106 19612
rect 7106 19556 7110 19612
rect 7046 19552 7110 19556
rect 7126 19612 7190 19616
rect 7126 19556 7130 19612
rect 7130 19556 7186 19612
rect 7186 19556 7190 19612
rect 7126 19552 7190 19556
rect 12820 19612 12884 19616
rect 12820 19556 12824 19612
rect 12824 19556 12880 19612
rect 12880 19556 12884 19612
rect 12820 19552 12884 19556
rect 12900 19612 12964 19616
rect 12900 19556 12904 19612
rect 12904 19556 12960 19612
rect 12960 19556 12964 19612
rect 12900 19552 12964 19556
rect 12980 19612 13044 19616
rect 12980 19556 12984 19612
rect 12984 19556 13040 19612
rect 13040 19556 13044 19612
rect 12980 19552 13044 19556
rect 13060 19612 13124 19616
rect 13060 19556 13064 19612
rect 13064 19556 13120 19612
rect 13120 19556 13124 19612
rect 13060 19552 13124 19556
rect 18754 19612 18818 19616
rect 18754 19556 18758 19612
rect 18758 19556 18814 19612
rect 18814 19556 18818 19612
rect 18754 19552 18818 19556
rect 18834 19612 18898 19616
rect 18834 19556 18838 19612
rect 18838 19556 18894 19612
rect 18894 19556 18898 19612
rect 18834 19552 18898 19556
rect 18914 19612 18978 19616
rect 18914 19556 18918 19612
rect 18918 19556 18974 19612
rect 18974 19556 18978 19612
rect 18914 19552 18978 19556
rect 18994 19612 19058 19616
rect 18994 19556 18998 19612
rect 18998 19556 19054 19612
rect 19054 19556 19058 19612
rect 18994 19552 19058 19556
rect 15148 19484 15212 19548
rect 9260 19348 9324 19412
rect 16804 19348 16868 19412
rect 24688 19612 24752 19616
rect 24688 19556 24692 19612
rect 24692 19556 24748 19612
rect 24748 19556 24752 19612
rect 24688 19552 24752 19556
rect 24768 19612 24832 19616
rect 24768 19556 24772 19612
rect 24772 19556 24828 19612
rect 24828 19556 24832 19612
rect 24768 19552 24832 19556
rect 24848 19612 24912 19616
rect 24848 19556 24852 19612
rect 24852 19556 24908 19612
rect 24908 19556 24912 19612
rect 24848 19552 24912 19556
rect 24928 19612 24992 19616
rect 24928 19556 24932 19612
rect 24932 19556 24988 19612
rect 24988 19556 24992 19612
rect 24928 19552 24992 19556
rect 4292 19212 4356 19276
rect 9628 19212 9692 19276
rect 16988 19212 17052 19276
rect 3919 19068 3983 19072
rect 3919 19012 3923 19068
rect 3923 19012 3979 19068
rect 3979 19012 3983 19068
rect 3919 19008 3983 19012
rect 3999 19068 4063 19072
rect 3999 19012 4003 19068
rect 4003 19012 4059 19068
rect 4059 19012 4063 19068
rect 3999 19008 4063 19012
rect 4079 19068 4143 19072
rect 4079 19012 4083 19068
rect 4083 19012 4139 19068
rect 4139 19012 4143 19068
rect 4079 19008 4143 19012
rect 4159 19068 4223 19072
rect 4159 19012 4163 19068
rect 4163 19012 4219 19068
rect 4219 19012 4223 19068
rect 4159 19008 4223 19012
rect 9853 19068 9917 19072
rect 9853 19012 9857 19068
rect 9857 19012 9913 19068
rect 9913 19012 9917 19068
rect 9853 19008 9917 19012
rect 9933 19068 9997 19072
rect 9933 19012 9937 19068
rect 9937 19012 9993 19068
rect 9993 19012 9997 19068
rect 9933 19008 9997 19012
rect 10013 19068 10077 19072
rect 10013 19012 10017 19068
rect 10017 19012 10073 19068
rect 10073 19012 10077 19068
rect 10013 19008 10077 19012
rect 10093 19068 10157 19072
rect 10093 19012 10097 19068
rect 10097 19012 10153 19068
rect 10153 19012 10157 19068
rect 10093 19008 10157 19012
rect 15787 19068 15851 19072
rect 15787 19012 15791 19068
rect 15791 19012 15847 19068
rect 15847 19012 15851 19068
rect 15787 19008 15851 19012
rect 15867 19068 15931 19072
rect 15867 19012 15871 19068
rect 15871 19012 15927 19068
rect 15927 19012 15931 19068
rect 15867 19008 15931 19012
rect 15947 19068 16011 19072
rect 15947 19012 15951 19068
rect 15951 19012 16007 19068
rect 16007 19012 16011 19068
rect 15947 19008 16011 19012
rect 16027 19068 16091 19072
rect 16027 19012 16031 19068
rect 16031 19012 16087 19068
rect 16087 19012 16091 19068
rect 16027 19008 16091 19012
rect 21721 19068 21785 19072
rect 21721 19012 21725 19068
rect 21725 19012 21781 19068
rect 21781 19012 21785 19068
rect 21721 19008 21785 19012
rect 21801 19068 21865 19072
rect 21801 19012 21805 19068
rect 21805 19012 21861 19068
rect 21861 19012 21865 19068
rect 21801 19008 21865 19012
rect 21881 19068 21945 19072
rect 21881 19012 21885 19068
rect 21885 19012 21941 19068
rect 21941 19012 21945 19068
rect 21881 19008 21945 19012
rect 21961 19068 22025 19072
rect 21961 19012 21965 19068
rect 21965 19012 22021 19068
rect 22021 19012 22025 19068
rect 21961 19008 22025 19012
rect 2084 18804 2148 18868
rect 17172 18804 17236 18868
rect 14412 18668 14476 18732
rect 15332 18668 15396 18732
rect 16436 18668 16500 18732
rect 6886 18524 6950 18528
rect 6886 18468 6890 18524
rect 6890 18468 6946 18524
rect 6946 18468 6950 18524
rect 6886 18464 6950 18468
rect 6966 18524 7030 18528
rect 6966 18468 6970 18524
rect 6970 18468 7026 18524
rect 7026 18468 7030 18524
rect 6966 18464 7030 18468
rect 7046 18524 7110 18528
rect 7046 18468 7050 18524
rect 7050 18468 7106 18524
rect 7106 18468 7110 18524
rect 7046 18464 7110 18468
rect 7126 18524 7190 18528
rect 7126 18468 7130 18524
rect 7130 18468 7186 18524
rect 7186 18468 7190 18524
rect 7126 18464 7190 18468
rect 12820 18524 12884 18528
rect 12820 18468 12824 18524
rect 12824 18468 12880 18524
rect 12880 18468 12884 18524
rect 12820 18464 12884 18468
rect 12900 18524 12964 18528
rect 12900 18468 12904 18524
rect 12904 18468 12960 18524
rect 12960 18468 12964 18524
rect 12900 18464 12964 18468
rect 12980 18524 13044 18528
rect 12980 18468 12984 18524
rect 12984 18468 13040 18524
rect 13040 18468 13044 18524
rect 12980 18464 13044 18468
rect 13060 18524 13124 18528
rect 13060 18468 13064 18524
rect 13064 18468 13120 18524
rect 13120 18468 13124 18524
rect 13060 18464 13124 18468
rect 18754 18524 18818 18528
rect 18754 18468 18758 18524
rect 18758 18468 18814 18524
rect 18814 18468 18818 18524
rect 18754 18464 18818 18468
rect 18834 18524 18898 18528
rect 18834 18468 18838 18524
rect 18838 18468 18894 18524
rect 18894 18468 18898 18524
rect 18834 18464 18898 18468
rect 18914 18524 18978 18528
rect 18914 18468 18918 18524
rect 18918 18468 18974 18524
rect 18974 18468 18978 18524
rect 18914 18464 18978 18468
rect 18994 18524 19058 18528
rect 18994 18468 18998 18524
rect 18998 18468 19054 18524
rect 19054 18468 19058 18524
rect 18994 18464 19058 18468
rect 24688 18524 24752 18528
rect 24688 18468 24692 18524
rect 24692 18468 24748 18524
rect 24748 18468 24752 18524
rect 24688 18464 24752 18468
rect 24768 18524 24832 18528
rect 24768 18468 24772 18524
rect 24772 18468 24828 18524
rect 24828 18468 24832 18524
rect 24768 18464 24832 18468
rect 24848 18524 24912 18528
rect 24848 18468 24852 18524
rect 24852 18468 24908 18524
rect 24908 18468 24912 18524
rect 24848 18464 24912 18468
rect 24928 18524 24992 18528
rect 24928 18468 24932 18524
rect 24932 18468 24988 18524
rect 24988 18468 24992 18524
rect 24928 18464 24992 18468
rect 1716 18260 1780 18324
rect 4476 17988 4540 18052
rect 10916 17988 10980 18052
rect 15516 18048 15580 18052
rect 15516 17992 15566 18048
rect 15566 17992 15580 18048
rect 15516 17988 15580 17992
rect 3919 17980 3983 17984
rect 3919 17924 3923 17980
rect 3923 17924 3979 17980
rect 3979 17924 3983 17980
rect 3919 17920 3983 17924
rect 3999 17980 4063 17984
rect 3999 17924 4003 17980
rect 4003 17924 4059 17980
rect 4059 17924 4063 17980
rect 3999 17920 4063 17924
rect 4079 17980 4143 17984
rect 4079 17924 4083 17980
rect 4083 17924 4139 17980
rect 4139 17924 4143 17980
rect 4079 17920 4143 17924
rect 4159 17980 4223 17984
rect 4159 17924 4163 17980
rect 4163 17924 4219 17980
rect 4219 17924 4223 17980
rect 4159 17920 4223 17924
rect 9853 17980 9917 17984
rect 9853 17924 9857 17980
rect 9857 17924 9913 17980
rect 9913 17924 9917 17980
rect 9853 17920 9917 17924
rect 9933 17980 9997 17984
rect 9933 17924 9937 17980
rect 9937 17924 9993 17980
rect 9993 17924 9997 17980
rect 9933 17920 9997 17924
rect 10013 17980 10077 17984
rect 10013 17924 10017 17980
rect 10017 17924 10073 17980
rect 10073 17924 10077 17980
rect 10013 17920 10077 17924
rect 10093 17980 10157 17984
rect 10093 17924 10097 17980
rect 10097 17924 10153 17980
rect 10153 17924 10157 17980
rect 10093 17920 10157 17924
rect 15787 17980 15851 17984
rect 15787 17924 15791 17980
rect 15791 17924 15847 17980
rect 15847 17924 15851 17980
rect 15787 17920 15851 17924
rect 15867 17980 15931 17984
rect 15867 17924 15871 17980
rect 15871 17924 15927 17980
rect 15927 17924 15931 17980
rect 15867 17920 15931 17924
rect 15947 17980 16011 17984
rect 15947 17924 15951 17980
rect 15951 17924 16007 17980
rect 16007 17924 16011 17980
rect 15947 17920 16011 17924
rect 16027 17980 16091 17984
rect 16027 17924 16031 17980
rect 16031 17924 16087 17980
rect 16087 17924 16091 17980
rect 16027 17920 16091 17924
rect 21721 17980 21785 17984
rect 21721 17924 21725 17980
rect 21725 17924 21781 17980
rect 21781 17924 21785 17980
rect 21721 17920 21785 17924
rect 21801 17980 21865 17984
rect 21801 17924 21805 17980
rect 21805 17924 21861 17980
rect 21861 17924 21865 17980
rect 21801 17920 21865 17924
rect 21881 17980 21945 17984
rect 21881 17924 21885 17980
rect 21885 17924 21941 17980
rect 21941 17924 21945 17980
rect 21881 17920 21945 17924
rect 21961 17980 22025 17984
rect 21961 17924 21965 17980
rect 21965 17924 22021 17980
rect 22021 17924 22025 17980
rect 21961 17920 22025 17924
rect 16252 17912 16316 17916
rect 16252 17856 16302 17912
rect 16302 17856 16316 17912
rect 16252 17852 16316 17856
rect 12572 17580 12636 17644
rect 6886 17436 6950 17440
rect 6886 17380 6890 17436
rect 6890 17380 6946 17436
rect 6946 17380 6950 17436
rect 6886 17376 6950 17380
rect 6966 17436 7030 17440
rect 6966 17380 6970 17436
rect 6970 17380 7026 17436
rect 7026 17380 7030 17436
rect 6966 17376 7030 17380
rect 7046 17436 7110 17440
rect 7046 17380 7050 17436
rect 7050 17380 7106 17436
rect 7106 17380 7110 17436
rect 7046 17376 7110 17380
rect 7126 17436 7190 17440
rect 7126 17380 7130 17436
rect 7130 17380 7186 17436
rect 7186 17380 7190 17436
rect 7126 17376 7190 17380
rect 12820 17436 12884 17440
rect 12820 17380 12824 17436
rect 12824 17380 12880 17436
rect 12880 17380 12884 17436
rect 12820 17376 12884 17380
rect 12900 17436 12964 17440
rect 12900 17380 12904 17436
rect 12904 17380 12960 17436
rect 12960 17380 12964 17436
rect 12900 17376 12964 17380
rect 12980 17436 13044 17440
rect 12980 17380 12984 17436
rect 12984 17380 13040 17436
rect 13040 17380 13044 17436
rect 12980 17376 13044 17380
rect 13060 17436 13124 17440
rect 13060 17380 13064 17436
rect 13064 17380 13120 17436
rect 13120 17380 13124 17436
rect 13060 17376 13124 17380
rect 18754 17436 18818 17440
rect 18754 17380 18758 17436
rect 18758 17380 18814 17436
rect 18814 17380 18818 17436
rect 18754 17376 18818 17380
rect 18834 17436 18898 17440
rect 18834 17380 18838 17436
rect 18838 17380 18894 17436
rect 18894 17380 18898 17436
rect 18834 17376 18898 17380
rect 18914 17436 18978 17440
rect 18914 17380 18918 17436
rect 18918 17380 18974 17436
rect 18974 17380 18978 17436
rect 18914 17376 18978 17380
rect 18994 17436 19058 17440
rect 18994 17380 18998 17436
rect 18998 17380 19054 17436
rect 19054 17380 19058 17436
rect 18994 17376 19058 17380
rect 24688 17436 24752 17440
rect 24688 17380 24692 17436
rect 24692 17380 24748 17436
rect 24748 17380 24752 17436
rect 24688 17376 24752 17380
rect 24768 17436 24832 17440
rect 24768 17380 24772 17436
rect 24772 17380 24828 17436
rect 24828 17380 24832 17436
rect 24768 17376 24832 17380
rect 24848 17436 24912 17440
rect 24848 17380 24852 17436
rect 24852 17380 24908 17436
rect 24908 17380 24912 17436
rect 24848 17376 24912 17380
rect 24928 17436 24992 17440
rect 24928 17380 24932 17436
rect 24932 17380 24988 17436
rect 24988 17380 24992 17436
rect 24928 17376 24992 17380
rect 16620 17172 16684 17236
rect 16988 17172 17052 17236
rect 20116 17172 20180 17236
rect 20300 17036 20364 17100
rect 2084 16960 2148 16964
rect 2084 16904 2098 16960
rect 2098 16904 2148 16960
rect 2084 16900 2148 16904
rect 8156 16900 8220 16964
rect 9444 16900 9508 16964
rect 3919 16892 3983 16896
rect 3919 16836 3923 16892
rect 3923 16836 3979 16892
rect 3979 16836 3983 16892
rect 3919 16832 3983 16836
rect 3999 16892 4063 16896
rect 3999 16836 4003 16892
rect 4003 16836 4059 16892
rect 4059 16836 4063 16892
rect 3999 16832 4063 16836
rect 4079 16892 4143 16896
rect 4079 16836 4083 16892
rect 4083 16836 4139 16892
rect 4139 16836 4143 16892
rect 4079 16832 4143 16836
rect 4159 16892 4223 16896
rect 4159 16836 4163 16892
rect 4163 16836 4219 16892
rect 4219 16836 4223 16892
rect 4159 16832 4223 16836
rect 9853 16892 9917 16896
rect 9853 16836 9857 16892
rect 9857 16836 9913 16892
rect 9913 16836 9917 16892
rect 9853 16832 9917 16836
rect 9933 16892 9997 16896
rect 9933 16836 9937 16892
rect 9937 16836 9993 16892
rect 9993 16836 9997 16892
rect 9933 16832 9997 16836
rect 10013 16892 10077 16896
rect 10013 16836 10017 16892
rect 10017 16836 10073 16892
rect 10073 16836 10077 16892
rect 10013 16832 10077 16836
rect 10093 16892 10157 16896
rect 10093 16836 10097 16892
rect 10097 16836 10153 16892
rect 10153 16836 10157 16892
rect 10093 16832 10157 16836
rect 15787 16892 15851 16896
rect 15787 16836 15791 16892
rect 15791 16836 15847 16892
rect 15847 16836 15851 16892
rect 15787 16832 15851 16836
rect 15867 16892 15931 16896
rect 15867 16836 15871 16892
rect 15871 16836 15927 16892
rect 15927 16836 15931 16892
rect 15867 16832 15931 16836
rect 15947 16892 16011 16896
rect 15947 16836 15951 16892
rect 15951 16836 16007 16892
rect 16007 16836 16011 16892
rect 15947 16832 16011 16836
rect 16027 16892 16091 16896
rect 16027 16836 16031 16892
rect 16031 16836 16087 16892
rect 16087 16836 16091 16892
rect 16027 16832 16091 16836
rect 21721 16892 21785 16896
rect 21721 16836 21725 16892
rect 21725 16836 21781 16892
rect 21781 16836 21785 16892
rect 21721 16832 21785 16836
rect 21801 16892 21865 16896
rect 21801 16836 21805 16892
rect 21805 16836 21861 16892
rect 21861 16836 21865 16892
rect 21801 16832 21865 16836
rect 21881 16892 21945 16896
rect 21881 16836 21885 16892
rect 21885 16836 21941 16892
rect 21941 16836 21945 16892
rect 21881 16832 21945 16836
rect 21961 16892 22025 16896
rect 21961 16836 21965 16892
rect 21965 16836 22021 16892
rect 22021 16836 22025 16892
rect 21961 16832 22025 16836
rect 12572 16688 12636 16692
rect 12572 16632 12586 16688
rect 12586 16632 12636 16688
rect 12572 16628 12636 16632
rect 15148 16628 15212 16692
rect 20668 16628 20732 16692
rect 2452 16552 2516 16556
rect 2452 16496 2466 16552
rect 2466 16496 2516 16552
rect 2452 16492 2516 16496
rect 5028 16492 5092 16556
rect 8708 16492 8772 16556
rect 19380 16552 19444 16556
rect 19380 16496 19394 16552
rect 19394 16496 19444 16552
rect 19380 16492 19444 16496
rect 6886 16348 6950 16352
rect 6886 16292 6890 16348
rect 6890 16292 6946 16348
rect 6946 16292 6950 16348
rect 6886 16288 6950 16292
rect 6966 16348 7030 16352
rect 6966 16292 6970 16348
rect 6970 16292 7026 16348
rect 7026 16292 7030 16348
rect 6966 16288 7030 16292
rect 7046 16348 7110 16352
rect 7046 16292 7050 16348
rect 7050 16292 7106 16348
rect 7106 16292 7110 16348
rect 7046 16288 7110 16292
rect 7126 16348 7190 16352
rect 7126 16292 7130 16348
rect 7130 16292 7186 16348
rect 7186 16292 7190 16348
rect 7126 16288 7190 16292
rect 12820 16348 12884 16352
rect 12820 16292 12824 16348
rect 12824 16292 12880 16348
rect 12880 16292 12884 16348
rect 12820 16288 12884 16292
rect 12900 16348 12964 16352
rect 12900 16292 12904 16348
rect 12904 16292 12960 16348
rect 12960 16292 12964 16348
rect 12900 16288 12964 16292
rect 12980 16348 13044 16352
rect 12980 16292 12984 16348
rect 12984 16292 13040 16348
rect 13040 16292 13044 16348
rect 12980 16288 13044 16292
rect 13060 16348 13124 16352
rect 13060 16292 13064 16348
rect 13064 16292 13120 16348
rect 13120 16292 13124 16348
rect 13060 16288 13124 16292
rect 18754 16348 18818 16352
rect 18754 16292 18758 16348
rect 18758 16292 18814 16348
rect 18814 16292 18818 16348
rect 18754 16288 18818 16292
rect 18834 16348 18898 16352
rect 18834 16292 18838 16348
rect 18838 16292 18894 16348
rect 18894 16292 18898 16348
rect 18834 16288 18898 16292
rect 18914 16348 18978 16352
rect 18914 16292 18918 16348
rect 18918 16292 18974 16348
rect 18974 16292 18978 16348
rect 18914 16288 18978 16292
rect 18994 16348 19058 16352
rect 18994 16292 18998 16348
rect 18998 16292 19054 16348
rect 19054 16292 19058 16348
rect 18994 16288 19058 16292
rect 24688 16348 24752 16352
rect 24688 16292 24692 16348
rect 24692 16292 24748 16348
rect 24748 16292 24752 16348
rect 24688 16288 24752 16292
rect 24768 16348 24832 16352
rect 24768 16292 24772 16348
rect 24772 16292 24828 16348
rect 24828 16292 24832 16348
rect 24768 16288 24832 16292
rect 24848 16348 24912 16352
rect 24848 16292 24852 16348
rect 24852 16292 24908 16348
rect 24908 16292 24912 16348
rect 24848 16288 24912 16292
rect 24928 16348 24992 16352
rect 24928 16292 24932 16348
rect 24932 16292 24988 16348
rect 24988 16292 24992 16348
rect 24928 16288 24992 16292
rect 3556 16220 3620 16284
rect 10916 16084 10980 16148
rect 17172 16084 17236 16148
rect 14044 15948 14108 16012
rect 3919 15804 3983 15808
rect 3919 15748 3923 15804
rect 3923 15748 3979 15804
rect 3979 15748 3983 15804
rect 3919 15744 3983 15748
rect 3999 15804 4063 15808
rect 3999 15748 4003 15804
rect 4003 15748 4059 15804
rect 4059 15748 4063 15804
rect 3999 15744 4063 15748
rect 4079 15804 4143 15808
rect 4079 15748 4083 15804
rect 4083 15748 4139 15804
rect 4139 15748 4143 15804
rect 4079 15744 4143 15748
rect 4159 15804 4223 15808
rect 4159 15748 4163 15804
rect 4163 15748 4219 15804
rect 4219 15748 4223 15804
rect 4159 15744 4223 15748
rect 9853 15804 9917 15808
rect 9853 15748 9857 15804
rect 9857 15748 9913 15804
rect 9913 15748 9917 15804
rect 9853 15744 9917 15748
rect 9933 15804 9997 15808
rect 9933 15748 9937 15804
rect 9937 15748 9993 15804
rect 9993 15748 9997 15804
rect 9933 15744 9997 15748
rect 10013 15804 10077 15808
rect 10013 15748 10017 15804
rect 10017 15748 10073 15804
rect 10073 15748 10077 15804
rect 10013 15744 10077 15748
rect 10093 15804 10157 15808
rect 10093 15748 10097 15804
rect 10097 15748 10153 15804
rect 10153 15748 10157 15804
rect 10093 15744 10157 15748
rect 15787 15804 15851 15808
rect 15787 15748 15791 15804
rect 15791 15748 15847 15804
rect 15847 15748 15851 15804
rect 15787 15744 15851 15748
rect 15867 15804 15931 15808
rect 15867 15748 15871 15804
rect 15871 15748 15927 15804
rect 15927 15748 15931 15804
rect 15867 15744 15931 15748
rect 15947 15804 16011 15808
rect 15947 15748 15951 15804
rect 15951 15748 16007 15804
rect 16007 15748 16011 15804
rect 15947 15744 16011 15748
rect 16027 15804 16091 15808
rect 16027 15748 16031 15804
rect 16031 15748 16087 15804
rect 16087 15748 16091 15804
rect 16027 15744 16091 15748
rect 21721 15804 21785 15808
rect 21721 15748 21725 15804
rect 21725 15748 21781 15804
rect 21781 15748 21785 15804
rect 21721 15744 21785 15748
rect 21801 15804 21865 15808
rect 21801 15748 21805 15804
rect 21805 15748 21861 15804
rect 21861 15748 21865 15804
rect 21801 15744 21865 15748
rect 21881 15804 21945 15808
rect 21881 15748 21885 15804
rect 21885 15748 21941 15804
rect 21941 15748 21945 15804
rect 21881 15744 21945 15748
rect 21961 15804 22025 15808
rect 21961 15748 21965 15804
rect 21965 15748 22021 15804
rect 22021 15748 22025 15804
rect 21961 15744 22025 15748
rect 4660 15540 4724 15604
rect 8340 15540 8404 15604
rect 13308 15404 13372 15468
rect 17356 15404 17420 15468
rect 22692 15404 22756 15468
rect 6886 15260 6950 15264
rect 6886 15204 6890 15260
rect 6890 15204 6946 15260
rect 6946 15204 6950 15260
rect 6886 15200 6950 15204
rect 6966 15260 7030 15264
rect 6966 15204 6970 15260
rect 6970 15204 7026 15260
rect 7026 15204 7030 15260
rect 6966 15200 7030 15204
rect 7046 15260 7110 15264
rect 7046 15204 7050 15260
rect 7050 15204 7106 15260
rect 7106 15204 7110 15260
rect 7046 15200 7110 15204
rect 7126 15260 7190 15264
rect 7126 15204 7130 15260
rect 7130 15204 7186 15260
rect 7186 15204 7190 15260
rect 7126 15200 7190 15204
rect 12820 15260 12884 15264
rect 12820 15204 12824 15260
rect 12824 15204 12880 15260
rect 12880 15204 12884 15260
rect 12820 15200 12884 15204
rect 12900 15260 12964 15264
rect 12900 15204 12904 15260
rect 12904 15204 12960 15260
rect 12960 15204 12964 15260
rect 12900 15200 12964 15204
rect 12980 15260 13044 15264
rect 12980 15204 12984 15260
rect 12984 15204 13040 15260
rect 13040 15204 13044 15260
rect 12980 15200 13044 15204
rect 13060 15260 13124 15264
rect 13060 15204 13064 15260
rect 13064 15204 13120 15260
rect 13120 15204 13124 15260
rect 13060 15200 13124 15204
rect 18754 15260 18818 15264
rect 18754 15204 18758 15260
rect 18758 15204 18814 15260
rect 18814 15204 18818 15260
rect 18754 15200 18818 15204
rect 18834 15260 18898 15264
rect 18834 15204 18838 15260
rect 18838 15204 18894 15260
rect 18894 15204 18898 15260
rect 18834 15200 18898 15204
rect 18914 15260 18978 15264
rect 18914 15204 18918 15260
rect 18918 15204 18974 15260
rect 18974 15204 18978 15260
rect 18914 15200 18978 15204
rect 18994 15260 19058 15264
rect 18994 15204 18998 15260
rect 18998 15204 19054 15260
rect 19054 15204 19058 15260
rect 18994 15200 19058 15204
rect 24688 15260 24752 15264
rect 24688 15204 24692 15260
rect 24692 15204 24748 15260
rect 24748 15204 24752 15260
rect 24688 15200 24752 15204
rect 24768 15260 24832 15264
rect 24768 15204 24772 15260
rect 24772 15204 24828 15260
rect 24828 15204 24832 15260
rect 24768 15200 24832 15204
rect 24848 15260 24912 15264
rect 24848 15204 24852 15260
rect 24852 15204 24908 15260
rect 24908 15204 24912 15260
rect 24848 15200 24912 15204
rect 24928 15260 24992 15264
rect 24928 15204 24932 15260
rect 24932 15204 24988 15260
rect 24988 15204 24992 15260
rect 24928 15200 24992 15204
rect 5212 15132 5276 15196
rect 10364 15132 10428 15196
rect 6500 14996 6564 15060
rect 3919 14716 3983 14720
rect 3919 14660 3923 14716
rect 3923 14660 3979 14716
rect 3979 14660 3983 14716
rect 3919 14656 3983 14660
rect 3999 14716 4063 14720
rect 3999 14660 4003 14716
rect 4003 14660 4059 14716
rect 4059 14660 4063 14716
rect 3999 14656 4063 14660
rect 4079 14716 4143 14720
rect 4079 14660 4083 14716
rect 4083 14660 4139 14716
rect 4139 14660 4143 14716
rect 4079 14656 4143 14660
rect 4159 14716 4223 14720
rect 4159 14660 4163 14716
rect 4163 14660 4219 14716
rect 4219 14660 4223 14716
rect 4159 14656 4223 14660
rect 9853 14716 9917 14720
rect 9853 14660 9857 14716
rect 9857 14660 9913 14716
rect 9913 14660 9917 14716
rect 9853 14656 9917 14660
rect 9933 14716 9997 14720
rect 9933 14660 9937 14716
rect 9937 14660 9993 14716
rect 9993 14660 9997 14716
rect 9933 14656 9997 14660
rect 10013 14716 10077 14720
rect 10013 14660 10017 14716
rect 10017 14660 10073 14716
rect 10073 14660 10077 14716
rect 10013 14656 10077 14660
rect 10093 14716 10157 14720
rect 10093 14660 10097 14716
rect 10097 14660 10153 14716
rect 10153 14660 10157 14716
rect 10093 14656 10157 14660
rect 15787 14716 15851 14720
rect 15787 14660 15791 14716
rect 15791 14660 15847 14716
rect 15847 14660 15851 14716
rect 15787 14656 15851 14660
rect 15867 14716 15931 14720
rect 15867 14660 15871 14716
rect 15871 14660 15927 14716
rect 15927 14660 15931 14716
rect 15867 14656 15931 14660
rect 15947 14716 16011 14720
rect 15947 14660 15951 14716
rect 15951 14660 16007 14716
rect 16007 14660 16011 14716
rect 15947 14656 16011 14660
rect 16027 14716 16091 14720
rect 16027 14660 16031 14716
rect 16031 14660 16087 14716
rect 16087 14660 16091 14716
rect 16027 14656 16091 14660
rect 21721 14716 21785 14720
rect 21721 14660 21725 14716
rect 21725 14660 21781 14716
rect 21781 14660 21785 14716
rect 21721 14656 21785 14660
rect 21801 14716 21865 14720
rect 21801 14660 21805 14716
rect 21805 14660 21861 14716
rect 21861 14660 21865 14716
rect 21801 14656 21865 14660
rect 21881 14716 21945 14720
rect 21881 14660 21885 14716
rect 21885 14660 21941 14716
rect 21941 14660 21945 14716
rect 21881 14656 21945 14660
rect 21961 14716 22025 14720
rect 21961 14660 21965 14716
rect 21965 14660 22021 14716
rect 22021 14660 22025 14716
rect 21961 14656 22025 14660
rect 6886 14172 6950 14176
rect 6886 14116 6890 14172
rect 6890 14116 6946 14172
rect 6946 14116 6950 14172
rect 6886 14112 6950 14116
rect 6966 14172 7030 14176
rect 6966 14116 6970 14172
rect 6970 14116 7026 14172
rect 7026 14116 7030 14172
rect 6966 14112 7030 14116
rect 7046 14172 7110 14176
rect 7046 14116 7050 14172
rect 7050 14116 7106 14172
rect 7106 14116 7110 14172
rect 7046 14112 7110 14116
rect 7126 14172 7190 14176
rect 7126 14116 7130 14172
rect 7130 14116 7186 14172
rect 7186 14116 7190 14172
rect 7126 14112 7190 14116
rect 12820 14172 12884 14176
rect 12820 14116 12824 14172
rect 12824 14116 12880 14172
rect 12880 14116 12884 14172
rect 12820 14112 12884 14116
rect 12900 14172 12964 14176
rect 12900 14116 12904 14172
rect 12904 14116 12960 14172
rect 12960 14116 12964 14172
rect 12900 14112 12964 14116
rect 12980 14172 13044 14176
rect 12980 14116 12984 14172
rect 12984 14116 13040 14172
rect 13040 14116 13044 14172
rect 12980 14112 13044 14116
rect 13060 14172 13124 14176
rect 13060 14116 13064 14172
rect 13064 14116 13120 14172
rect 13120 14116 13124 14172
rect 13060 14112 13124 14116
rect 18754 14172 18818 14176
rect 18754 14116 18758 14172
rect 18758 14116 18814 14172
rect 18814 14116 18818 14172
rect 18754 14112 18818 14116
rect 18834 14172 18898 14176
rect 18834 14116 18838 14172
rect 18838 14116 18894 14172
rect 18894 14116 18898 14172
rect 18834 14112 18898 14116
rect 18914 14172 18978 14176
rect 18914 14116 18918 14172
rect 18918 14116 18974 14172
rect 18974 14116 18978 14172
rect 18914 14112 18978 14116
rect 18994 14172 19058 14176
rect 18994 14116 18998 14172
rect 18998 14116 19054 14172
rect 19054 14116 19058 14172
rect 18994 14112 19058 14116
rect 24688 14172 24752 14176
rect 24688 14116 24692 14172
rect 24692 14116 24748 14172
rect 24748 14116 24752 14172
rect 24688 14112 24752 14116
rect 24768 14172 24832 14176
rect 24768 14116 24772 14172
rect 24772 14116 24828 14172
rect 24828 14116 24832 14172
rect 24768 14112 24832 14116
rect 24848 14172 24912 14176
rect 24848 14116 24852 14172
rect 24852 14116 24908 14172
rect 24908 14116 24912 14172
rect 24848 14112 24912 14116
rect 24928 14172 24992 14176
rect 24928 14116 24932 14172
rect 24932 14116 24988 14172
rect 24988 14116 24992 14172
rect 24928 14112 24992 14116
rect 4844 13772 4908 13836
rect 2268 13636 2332 13700
rect 9628 13636 9692 13700
rect 3919 13628 3983 13632
rect 3919 13572 3923 13628
rect 3923 13572 3979 13628
rect 3979 13572 3983 13628
rect 3919 13568 3983 13572
rect 3999 13628 4063 13632
rect 3999 13572 4003 13628
rect 4003 13572 4059 13628
rect 4059 13572 4063 13628
rect 3999 13568 4063 13572
rect 4079 13628 4143 13632
rect 4079 13572 4083 13628
rect 4083 13572 4139 13628
rect 4139 13572 4143 13628
rect 4079 13568 4143 13572
rect 4159 13628 4223 13632
rect 4159 13572 4163 13628
rect 4163 13572 4219 13628
rect 4219 13572 4223 13628
rect 4159 13568 4223 13572
rect 9853 13628 9917 13632
rect 9853 13572 9857 13628
rect 9857 13572 9913 13628
rect 9913 13572 9917 13628
rect 9853 13568 9917 13572
rect 9933 13628 9997 13632
rect 9933 13572 9937 13628
rect 9937 13572 9993 13628
rect 9993 13572 9997 13628
rect 9933 13568 9997 13572
rect 10013 13628 10077 13632
rect 10013 13572 10017 13628
rect 10017 13572 10073 13628
rect 10073 13572 10077 13628
rect 10013 13568 10077 13572
rect 10093 13628 10157 13632
rect 10093 13572 10097 13628
rect 10097 13572 10153 13628
rect 10153 13572 10157 13628
rect 10093 13568 10157 13572
rect 19932 13636 19996 13700
rect 15787 13628 15851 13632
rect 15787 13572 15791 13628
rect 15791 13572 15847 13628
rect 15847 13572 15851 13628
rect 15787 13568 15851 13572
rect 15867 13628 15931 13632
rect 15867 13572 15871 13628
rect 15871 13572 15927 13628
rect 15927 13572 15931 13628
rect 15867 13568 15931 13572
rect 15947 13628 16011 13632
rect 15947 13572 15951 13628
rect 15951 13572 16007 13628
rect 16007 13572 16011 13628
rect 15947 13568 16011 13572
rect 16027 13628 16091 13632
rect 16027 13572 16031 13628
rect 16031 13572 16087 13628
rect 16087 13572 16091 13628
rect 16027 13568 16091 13572
rect 21721 13628 21785 13632
rect 21721 13572 21725 13628
rect 21725 13572 21781 13628
rect 21781 13572 21785 13628
rect 21721 13568 21785 13572
rect 21801 13628 21865 13632
rect 21801 13572 21805 13628
rect 21805 13572 21861 13628
rect 21861 13572 21865 13628
rect 21801 13568 21865 13572
rect 21881 13628 21945 13632
rect 21881 13572 21885 13628
rect 21885 13572 21941 13628
rect 21941 13572 21945 13628
rect 21881 13568 21945 13572
rect 21961 13628 22025 13632
rect 21961 13572 21965 13628
rect 21965 13572 22021 13628
rect 22021 13572 22025 13628
rect 21961 13568 22025 13572
rect 20852 13500 20916 13564
rect 9260 13364 9324 13428
rect 3556 13228 3620 13292
rect 6886 13084 6950 13088
rect 6886 13028 6890 13084
rect 6890 13028 6946 13084
rect 6946 13028 6950 13084
rect 6886 13024 6950 13028
rect 6966 13084 7030 13088
rect 6966 13028 6970 13084
rect 6970 13028 7026 13084
rect 7026 13028 7030 13084
rect 6966 13024 7030 13028
rect 7046 13084 7110 13088
rect 7046 13028 7050 13084
rect 7050 13028 7106 13084
rect 7106 13028 7110 13084
rect 7046 13024 7110 13028
rect 7126 13084 7190 13088
rect 7126 13028 7130 13084
rect 7130 13028 7186 13084
rect 7186 13028 7190 13084
rect 7126 13024 7190 13028
rect 12820 13084 12884 13088
rect 12820 13028 12824 13084
rect 12824 13028 12880 13084
rect 12880 13028 12884 13084
rect 12820 13024 12884 13028
rect 12900 13084 12964 13088
rect 12900 13028 12904 13084
rect 12904 13028 12960 13084
rect 12960 13028 12964 13084
rect 12900 13024 12964 13028
rect 12980 13084 13044 13088
rect 12980 13028 12984 13084
rect 12984 13028 13040 13084
rect 13040 13028 13044 13084
rect 12980 13024 13044 13028
rect 13060 13084 13124 13088
rect 13060 13028 13064 13084
rect 13064 13028 13120 13084
rect 13120 13028 13124 13084
rect 13060 13024 13124 13028
rect 18754 13084 18818 13088
rect 18754 13028 18758 13084
rect 18758 13028 18814 13084
rect 18814 13028 18818 13084
rect 18754 13024 18818 13028
rect 18834 13084 18898 13088
rect 18834 13028 18838 13084
rect 18838 13028 18894 13084
rect 18894 13028 18898 13084
rect 18834 13024 18898 13028
rect 18914 13084 18978 13088
rect 18914 13028 18918 13084
rect 18918 13028 18974 13084
rect 18974 13028 18978 13084
rect 18914 13024 18978 13028
rect 18994 13084 19058 13088
rect 18994 13028 18998 13084
rect 18998 13028 19054 13084
rect 19054 13028 19058 13084
rect 18994 13024 19058 13028
rect 24688 13084 24752 13088
rect 24688 13028 24692 13084
rect 24692 13028 24748 13084
rect 24748 13028 24752 13084
rect 24688 13024 24752 13028
rect 24768 13084 24832 13088
rect 24768 13028 24772 13084
rect 24772 13028 24828 13084
rect 24828 13028 24832 13084
rect 24768 13024 24832 13028
rect 24848 13084 24912 13088
rect 24848 13028 24852 13084
rect 24852 13028 24908 13084
rect 24908 13028 24912 13084
rect 24848 13024 24912 13028
rect 24928 13084 24992 13088
rect 24928 13028 24932 13084
rect 24932 13028 24988 13084
rect 24988 13028 24992 13084
rect 24928 13024 24992 13028
rect 3919 12540 3983 12544
rect 3919 12484 3923 12540
rect 3923 12484 3979 12540
rect 3979 12484 3983 12540
rect 3919 12480 3983 12484
rect 3999 12540 4063 12544
rect 3999 12484 4003 12540
rect 4003 12484 4059 12540
rect 4059 12484 4063 12540
rect 3999 12480 4063 12484
rect 4079 12540 4143 12544
rect 4079 12484 4083 12540
rect 4083 12484 4139 12540
rect 4139 12484 4143 12540
rect 4079 12480 4143 12484
rect 4159 12540 4223 12544
rect 4159 12484 4163 12540
rect 4163 12484 4219 12540
rect 4219 12484 4223 12540
rect 4159 12480 4223 12484
rect 9853 12540 9917 12544
rect 9853 12484 9857 12540
rect 9857 12484 9913 12540
rect 9913 12484 9917 12540
rect 9853 12480 9917 12484
rect 9933 12540 9997 12544
rect 9933 12484 9937 12540
rect 9937 12484 9993 12540
rect 9993 12484 9997 12540
rect 9933 12480 9997 12484
rect 10013 12540 10077 12544
rect 10013 12484 10017 12540
rect 10017 12484 10073 12540
rect 10073 12484 10077 12540
rect 10013 12480 10077 12484
rect 10093 12540 10157 12544
rect 10093 12484 10097 12540
rect 10097 12484 10153 12540
rect 10153 12484 10157 12540
rect 10093 12480 10157 12484
rect 15787 12540 15851 12544
rect 15787 12484 15791 12540
rect 15791 12484 15847 12540
rect 15847 12484 15851 12540
rect 15787 12480 15851 12484
rect 15867 12540 15931 12544
rect 15867 12484 15871 12540
rect 15871 12484 15927 12540
rect 15927 12484 15931 12540
rect 15867 12480 15931 12484
rect 15947 12540 16011 12544
rect 15947 12484 15951 12540
rect 15951 12484 16007 12540
rect 16007 12484 16011 12540
rect 15947 12480 16011 12484
rect 16027 12540 16091 12544
rect 16027 12484 16031 12540
rect 16031 12484 16087 12540
rect 16087 12484 16091 12540
rect 16027 12480 16091 12484
rect 21721 12540 21785 12544
rect 21721 12484 21725 12540
rect 21725 12484 21781 12540
rect 21781 12484 21785 12540
rect 21721 12480 21785 12484
rect 21801 12540 21865 12544
rect 21801 12484 21805 12540
rect 21805 12484 21861 12540
rect 21861 12484 21865 12540
rect 21801 12480 21865 12484
rect 21881 12540 21945 12544
rect 21881 12484 21885 12540
rect 21885 12484 21941 12540
rect 21941 12484 21945 12540
rect 21881 12480 21945 12484
rect 21961 12540 22025 12544
rect 21961 12484 21965 12540
rect 21965 12484 22021 12540
rect 22021 12484 22025 12540
rect 21961 12480 22025 12484
rect 3188 12472 3252 12476
rect 3188 12416 3238 12472
rect 3238 12416 3252 12472
rect 3188 12412 3252 12416
rect 6500 12412 6564 12476
rect 5396 12276 5460 12340
rect 10916 12276 10980 12340
rect 8892 12140 8956 12204
rect 4660 12004 4724 12068
rect 6886 11996 6950 12000
rect 6886 11940 6890 11996
rect 6890 11940 6946 11996
rect 6946 11940 6950 11996
rect 6886 11936 6950 11940
rect 6966 11996 7030 12000
rect 6966 11940 6970 11996
rect 6970 11940 7026 11996
rect 7026 11940 7030 11996
rect 6966 11936 7030 11940
rect 7046 11996 7110 12000
rect 7046 11940 7050 11996
rect 7050 11940 7106 11996
rect 7106 11940 7110 11996
rect 7046 11936 7110 11940
rect 7126 11996 7190 12000
rect 7126 11940 7130 11996
rect 7130 11940 7186 11996
rect 7186 11940 7190 11996
rect 7126 11936 7190 11940
rect 12820 11996 12884 12000
rect 12820 11940 12824 11996
rect 12824 11940 12880 11996
rect 12880 11940 12884 11996
rect 12820 11936 12884 11940
rect 12900 11996 12964 12000
rect 12900 11940 12904 11996
rect 12904 11940 12960 11996
rect 12960 11940 12964 11996
rect 12900 11936 12964 11940
rect 12980 11996 13044 12000
rect 12980 11940 12984 11996
rect 12984 11940 13040 11996
rect 13040 11940 13044 11996
rect 12980 11936 13044 11940
rect 13060 11996 13124 12000
rect 13060 11940 13064 11996
rect 13064 11940 13120 11996
rect 13120 11940 13124 11996
rect 13060 11936 13124 11940
rect 18754 11996 18818 12000
rect 18754 11940 18758 11996
rect 18758 11940 18814 11996
rect 18814 11940 18818 11996
rect 18754 11936 18818 11940
rect 18834 11996 18898 12000
rect 18834 11940 18838 11996
rect 18838 11940 18894 11996
rect 18894 11940 18898 11996
rect 18834 11936 18898 11940
rect 18914 11996 18978 12000
rect 18914 11940 18918 11996
rect 18918 11940 18974 11996
rect 18974 11940 18978 11996
rect 18914 11936 18978 11940
rect 18994 11996 19058 12000
rect 18994 11940 18998 11996
rect 18998 11940 19054 11996
rect 19054 11940 19058 11996
rect 18994 11936 19058 11940
rect 24688 11996 24752 12000
rect 24688 11940 24692 11996
rect 24692 11940 24748 11996
rect 24748 11940 24752 11996
rect 24688 11936 24752 11940
rect 24768 11996 24832 12000
rect 24768 11940 24772 11996
rect 24772 11940 24828 11996
rect 24828 11940 24832 11996
rect 24768 11936 24832 11940
rect 24848 11996 24912 12000
rect 24848 11940 24852 11996
rect 24852 11940 24908 11996
rect 24908 11940 24912 11996
rect 24848 11936 24912 11940
rect 24928 11996 24992 12000
rect 24928 11940 24932 11996
rect 24932 11940 24988 11996
rect 24988 11940 24992 11996
rect 24928 11936 24992 11940
rect 15332 11868 15396 11932
rect 3919 11452 3983 11456
rect 3919 11396 3923 11452
rect 3923 11396 3979 11452
rect 3979 11396 3983 11452
rect 3919 11392 3983 11396
rect 3999 11452 4063 11456
rect 3999 11396 4003 11452
rect 4003 11396 4059 11452
rect 4059 11396 4063 11452
rect 3999 11392 4063 11396
rect 4079 11452 4143 11456
rect 4079 11396 4083 11452
rect 4083 11396 4139 11452
rect 4139 11396 4143 11452
rect 4079 11392 4143 11396
rect 4159 11452 4223 11456
rect 4159 11396 4163 11452
rect 4163 11396 4219 11452
rect 4219 11396 4223 11452
rect 4159 11392 4223 11396
rect 9853 11452 9917 11456
rect 9853 11396 9857 11452
rect 9857 11396 9913 11452
rect 9913 11396 9917 11452
rect 9853 11392 9917 11396
rect 9933 11452 9997 11456
rect 9933 11396 9937 11452
rect 9937 11396 9993 11452
rect 9993 11396 9997 11452
rect 9933 11392 9997 11396
rect 10013 11452 10077 11456
rect 10013 11396 10017 11452
rect 10017 11396 10073 11452
rect 10073 11396 10077 11452
rect 10013 11392 10077 11396
rect 10093 11452 10157 11456
rect 10093 11396 10097 11452
rect 10097 11396 10153 11452
rect 10153 11396 10157 11452
rect 10093 11392 10157 11396
rect 15787 11452 15851 11456
rect 15787 11396 15791 11452
rect 15791 11396 15847 11452
rect 15847 11396 15851 11452
rect 15787 11392 15851 11396
rect 15867 11452 15931 11456
rect 15867 11396 15871 11452
rect 15871 11396 15927 11452
rect 15927 11396 15931 11452
rect 15867 11392 15931 11396
rect 15947 11452 16011 11456
rect 15947 11396 15951 11452
rect 15951 11396 16007 11452
rect 16007 11396 16011 11452
rect 15947 11392 16011 11396
rect 16027 11452 16091 11456
rect 16027 11396 16031 11452
rect 16031 11396 16087 11452
rect 16087 11396 16091 11452
rect 16027 11392 16091 11396
rect 21721 11452 21785 11456
rect 21721 11396 21725 11452
rect 21725 11396 21781 11452
rect 21781 11396 21785 11452
rect 21721 11392 21785 11396
rect 21801 11452 21865 11456
rect 21801 11396 21805 11452
rect 21805 11396 21861 11452
rect 21861 11396 21865 11452
rect 21801 11392 21865 11396
rect 21881 11452 21945 11456
rect 21881 11396 21885 11452
rect 21885 11396 21941 11452
rect 21941 11396 21945 11452
rect 21881 11392 21945 11396
rect 21961 11452 22025 11456
rect 21961 11396 21965 11452
rect 21965 11396 22021 11452
rect 22021 11396 22025 11452
rect 21961 11392 22025 11396
rect 8340 11188 8404 11252
rect 4476 10916 4540 10980
rect 6886 10908 6950 10912
rect 6886 10852 6890 10908
rect 6890 10852 6946 10908
rect 6946 10852 6950 10908
rect 6886 10848 6950 10852
rect 6966 10908 7030 10912
rect 6966 10852 6970 10908
rect 6970 10852 7026 10908
rect 7026 10852 7030 10908
rect 6966 10848 7030 10852
rect 7046 10908 7110 10912
rect 7046 10852 7050 10908
rect 7050 10852 7106 10908
rect 7106 10852 7110 10908
rect 7046 10848 7110 10852
rect 7126 10908 7190 10912
rect 7126 10852 7130 10908
rect 7130 10852 7186 10908
rect 7186 10852 7190 10908
rect 7126 10848 7190 10852
rect 12820 10908 12884 10912
rect 12820 10852 12824 10908
rect 12824 10852 12880 10908
rect 12880 10852 12884 10908
rect 12820 10848 12884 10852
rect 12900 10908 12964 10912
rect 12900 10852 12904 10908
rect 12904 10852 12960 10908
rect 12960 10852 12964 10908
rect 12900 10848 12964 10852
rect 12980 10908 13044 10912
rect 12980 10852 12984 10908
rect 12984 10852 13040 10908
rect 13040 10852 13044 10908
rect 12980 10848 13044 10852
rect 13060 10908 13124 10912
rect 13060 10852 13064 10908
rect 13064 10852 13120 10908
rect 13120 10852 13124 10908
rect 13060 10848 13124 10852
rect 18754 10908 18818 10912
rect 18754 10852 18758 10908
rect 18758 10852 18814 10908
rect 18814 10852 18818 10908
rect 18754 10848 18818 10852
rect 18834 10908 18898 10912
rect 18834 10852 18838 10908
rect 18838 10852 18894 10908
rect 18894 10852 18898 10908
rect 18834 10848 18898 10852
rect 18914 10908 18978 10912
rect 18914 10852 18918 10908
rect 18918 10852 18974 10908
rect 18974 10852 18978 10908
rect 18914 10848 18978 10852
rect 18994 10908 19058 10912
rect 18994 10852 18998 10908
rect 18998 10852 19054 10908
rect 19054 10852 19058 10908
rect 18994 10848 19058 10852
rect 24688 10908 24752 10912
rect 24688 10852 24692 10908
rect 24692 10852 24748 10908
rect 24748 10852 24752 10908
rect 24688 10848 24752 10852
rect 24768 10908 24832 10912
rect 24768 10852 24772 10908
rect 24772 10852 24828 10908
rect 24828 10852 24832 10908
rect 24768 10848 24832 10852
rect 24848 10908 24912 10912
rect 24848 10852 24852 10908
rect 24852 10852 24908 10908
rect 24908 10852 24912 10908
rect 24848 10848 24912 10852
rect 24928 10908 24992 10912
rect 24928 10852 24932 10908
rect 24932 10852 24988 10908
rect 24988 10852 24992 10908
rect 24928 10848 24992 10852
rect 3919 10364 3983 10368
rect 3919 10308 3923 10364
rect 3923 10308 3979 10364
rect 3979 10308 3983 10364
rect 3919 10304 3983 10308
rect 3999 10364 4063 10368
rect 3999 10308 4003 10364
rect 4003 10308 4059 10364
rect 4059 10308 4063 10364
rect 3999 10304 4063 10308
rect 4079 10364 4143 10368
rect 4079 10308 4083 10364
rect 4083 10308 4139 10364
rect 4139 10308 4143 10364
rect 4079 10304 4143 10308
rect 4159 10364 4223 10368
rect 4159 10308 4163 10364
rect 4163 10308 4219 10364
rect 4219 10308 4223 10364
rect 4159 10304 4223 10308
rect 3004 10296 3068 10300
rect 3004 10240 3054 10296
rect 3054 10240 3068 10296
rect 3004 10236 3068 10240
rect 2084 10160 2148 10164
rect 2084 10104 2134 10160
rect 2134 10104 2148 10160
rect 2084 10100 2148 10104
rect 1900 9828 1964 9892
rect 3004 9752 3068 9756
rect 3004 9696 3018 9752
rect 3018 9696 3068 9752
rect 3004 9692 3068 9696
rect 3188 9752 3252 9756
rect 11100 10508 11164 10572
rect 9853 10364 9917 10368
rect 9853 10308 9857 10364
rect 9857 10308 9913 10364
rect 9913 10308 9917 10364
rect 9853 10304 9917 10308
rect 9933 10364 9997 10368
rect 9933 10308 9937 10364
rect 9937 10308 9993 10364
rect 9993 10308 9997 10364
rect 9933 10304 9997 10308
rect 10013 10364 10077 10368
rect 10013 10308 10017 10364
rect 10017 10308 10073 10364
rect 10073 10308 10077 10364
rect 10013 10304 10077 10308
rect 10093 10364 10157 10368
rect 10093 10308 10097 10364
rect 10097 10308 10153 10364
rect 10153 10308 10157 10364
rect 10093 10304 10157 10308
rect 15787 10364 15851 10368
rect 15787 10308 15791 10364
rect 15791 10308 15847 10364
rect 15847 10308 15851 10364
rect 15787 10304 15851 10308
rect 15867 10364 15931 10368
rect 15867 10308 15871 10364
rect 15871 10308 15927 10364
rect 15927 10308 15931 10364
rect 15867 10304 15931 10308
rect 15947 10364 16011 10368
rect 15947 10308 15951 10364
rect 15951 10308 16007 10364
rect 16007 10308 16011 10364
rect 15947 10304 16011 10308
rect 16027 10364 16091 10368
rect 16027 10308 16031 10364
rect 16031 10308 16087 10364
rect 16087 10308 16091 10364
rect 16027 10304 16091 10308
rect 21721 10364 21785 10368
rect 21721 10308 21725 10364
rect 21725 10308 21781 10364
rect 21781 10308 21785 10364
rect 21721 10304 21785 10308
rect 21801 10364 21865 10368
rect 21801 10308 21805 10364
rect 21805 10308 21861 10364
rect 21861 10308 21865 10364
rect 21801 10304 21865 10308
rect 21881 10364 21945 10368
rect 21881 10308 21885 10364
rect 21885 10308 21941 10364
rect 21941 10308 21945 10364
rect 21881 10304 21945 10308
rect 21961 10364 22025 10368
rect 21961 10308 21965 10364
rect 21965 10308 22021 10364
rect 22021 10308 22025 10364
rect 21961 10304 22025 10308
rect 9076 9964 9140 10028
rect 10364 10100 10428 10164
rect 21588 10100 21652 10164
rect 11468 9964 11532 10028
rect 14596 9828 14660 9892
rect 6886 9820 6950 9824
rect 6886 9764 6890 9820
rect 6890 9764 6946 9820
rect 6946 9764 6950 9820
rect 6886 9760 6950 9764
rect 6966 9820 7030 9824
rect 6966 9764 6970 9820
rect 6970 9764 7026 9820
rect 7026 9764 7030 9820
rect 6966 9760 7030 9764
rect 7046 9820 7110 9824
rect 7046 9764 7050 9820
rect 7050 9764 7106 9820
rect 7106 9764 7110 9820
rect 7046 9760 7110 9764
rect 7126 9820 7190 9824
rect 7126 9764 7130 9820
rect 7130 9764 7186 9820
rect 7186 9764 7190 9820
rect 7126 9760 7190 9764
rect 12820 9820 12884 9824
rect 12820 9764 12824 9820
rect 12824 9764 12880 9820
rect 12880 9764 12884 9820
rect 12820 9760 12884 9764
rect 12900 9820 12964 9824
rect 12900 9764 12904 9820
rect 12904 9764 12960 9820
rect 12960 9764 12964 9820
rect 12900 9760 12964 9764
rect 12980 9820 13044 9824
rect 12980 9764 12984 9820
rect 12984 9764 13040 9820
rect 13040 9764 13044 9820
rect 12980 9760 13044 9764
rect 13060 9820 13124 9824
rect 13060 9764 13064 9820
rect 13064 9764 13120 9820
rect 13120 9764 13124 9820
rect 13060 9760 13124 9764
rect 18754 9820 18818 9824
rect 18754 9764 18758 9820
rect 18758 9764 18814 9820
rect 18814 9764 18818 9820
rect 18754 9760 18818 9764
rect 18834 9820 18898 9824
rect 18834 9764 18838 9820
rect 18838 9764 18894 9820
rect 18894 9764 18898 9820
rect 18834 9760 18898 9764
rect 18914 9820 18978 9824
rect 18914 9764 18918 9820
rect 18918 9764 18974 9820
rect 18974 9764 18978 9820
rect 18914 9760 18978 9764
rect 18994 9820 19058 9824
rect 18994 9764 18998 9820
rect 18998 9764 19054 9820
rect 19054 9764 19058 9820
rect 18994 9760 19058 9764
rect 24688 9820 24752 9824
rect 24688 9764 24692 9820
rect 24692 9764 24748 9820
rect 24748 9764 24752 9820
rect 24688 9760 24752 9764
rect 24768 9820 24832 9824
rect 24768 9764 24772 9820
rect 24772 9764 24828 9820
rect 24828 9764 24832 9820
rect 24768 9760 24832 9764
rect 24848 9820 24912 9824
rect 24848 9764 24852 9820
rect 24852 9764 24908 9820
rect 24908 9764 24912 9820
rect 24848 9760 24912 9764
rect 24928 9820 24992 9824
rect 24928 9764 24932 9820
rect 24932 9764 24988 9820
rect 24988 9764 24992 9820
rect 24928 9760 24992 9764
rect 3188 9696 3202 9752
rect 3202 9696 3252 9752
rect 3188 9692 3252 9696
rect 12204 9692 12268 9756
rect 16804 9692 16868 9756
rect 19748 9420 19812 9484
rect 3919 9276 3983 9280
rect 3919 9220 3923 9276
rect 3923 9220 3979 9276
rect 3979 9220 3983 9276
rect 3919 9216 3983 9220
rect 3999 9276 4063 9280
rect 3999 9220 4003 9276
rect 4003 9220 4059 9276
rect 4059 9220 4063 9276
rect 3999 9216 4063 9220
rect 4079 9276 4143 9280
rect 4079 9220 4083 9276
rect 4083 9220 4139 9276
rect 4139 9220 4143 9276
rect 4079 9216 4143 9220
rect 4159 9276 4223 9280
rect 4159 9220 4163 9276
rect 4163 9220 4219 9276
rect 4219 9220 4223 9276
rect 4159 9216 4223 9220
rect 9853 9276 9917 9280
rect 9853 9220 9857 9276
rect 9857 9220 9913 9276
rect 9913 9220 9917 9276
rect 9853 9216 9917 9220
rect 9933 9276 9997 9280
rect 9933 9220 9937 9276
rect 9937 9220 9993 9276
rect 9993 9220 9997 9276
rect 9933 9216 9997 9220
rect 10013 9276 10077 9280
rect 10013 9220 10017 9276
rect 10017 9220 10073 9276
rect 10073 9220 10077 9276
rect 10013 9216 10077 9220
rect 10093 9276 10157 9280
rect 10093 9220 10097 9276
rect 10097 9220 10153 9276
rect 10153 9220 10157 9276
rect 10093 9216 10157 9220
rect 15787 9276 15851 9280
rect 15787 9220 15791 9276
rect 15791 9220 15847 9276
rect 15847 9220 15851 9276
rect 15787 9216 15851 9220
rect 15867 9276 15931 9280
rect 15867 9220 15871 9276
rect 15871 9220 15927 9276
rect 15927 9220 15931 9276
rect 15867 9216 15931 9220
rect 15947 9276 16011 9280
rect 15947 9220 15951 9276
rect 15951 9220 16007 9276
rect 16007 9220 16011 9276
rect 15947 9216 16011 9220
rect 16027 9276 16091 9280
rect 16027 9220 16031 9276
rect 16031 9220 16087 9276
rect 16087 9220 16091 9276
rect 16027 9216 16091 9220
rect 21721 9276 21785 9280
rect 21721 9220 21725 9276
rect 21725 9220 21781 9276
rect 21781 9220 21785 9276
rect 21721 9216 21785 9220
rect 21801 9276 21865 9280
rect 21801 9220 21805 9276
rect 21805 9220 21861 9276
rect 21861 9220 21865 9276
rect 21801 9216 21865 9220
rect 21881 9276 21945 9280
rect 21881 9220 21885 9276
rect 21885 9220 21941 9276
rect 21941 9220 21945 9276
rect 21881 9216 21945 9220
rect 21961 9276 22025 9280
rect 21961 9220 21965 9276
rect 21965 9220 22021 9276
rect 22021 9220 22025 9276
rect 21961 9216 22025 9220
rect 15332 9012 15396 9076
rect 6886 8732 6950 8736
rect 6886 8676 6890 8732
rect 6890 8676 6946 8732
rect 6946 8676 6950 8732
rect 6886 8672 6950 8676
rect 6966 8732 7030 8736
rect 6966 8676 6970 8732
rect 6970 8676 7026 8732
rect 7026 8676 7030 8732
rect 6966 8672 7030 8676
rect 7046 8732 7110 8736
rect 7046 8676 7050 8732
rect 7050 8676 7106 8732
rect 7106 8676 7110 8732
rect 7046 8672 7110 8676
rect 7126 8732 7190 8736
rect 7126 8676 7130 8732
rect 7130 8676 7186 8732
rect 7186 8676 7190 8732
rect 7126 8672 7190 8676
rect 12820 8732 12884 8736
rect 12820 8676 12824 8732
rect 12824 8676 12880 8732
rect 12880 8676 12884 8732
rect 12820 8672 12884 8676
rect 12900 8732 12964 8736
rect 12900 8676 12904 8732
rect 12904 8676 12960 8732
rect 12960 8676 12964 8732
rect 12900 8672 12964 8676
rect 12980 8732 13044 8736
rect 12980 8676 12984 8732
rect 12984 8676 13040 8732
rect 13040 8676 13044 8732
rect 12980 8672 13044 8676
rect 13060 8732 13124 8736
rect 13060 8676 13064 8732
rect 13064 8676 13120 8732
rect 13120 8676 13124 8732
rect 13060 8672 13124 8676
rect 18754 8732 18818 8736
rect 18754 8676 18758 8732
rect 18758 8676 18814 8732
rect 18814 8676 18818 8732
rect 18754 8672 18818 8676
rect 18834 8732 18898 8736
rect 18834 8676 18838 8732
rect 18838 8676 18894 8732
rect 18894 8676 18898 8732
rect 18834 8672 18898 8676
rect 18914 8732 18978 8736
rect 18914 8676 18918 8732
rect 18918 8676 18974 8732
rect 18974 8676 18978 8732
rect 18914 8672 18978 8676
rect 18994 8732 19058 8736
rect 18994 8676 18998 8732
rect 18998 8676 19054 8732
rect 19054 8676 19058 8732
rect 18994 8672 19058 8676
rect 24688 8732 24752 8736
rect 24688 8676 24692 8732
rect 24692 8676 24748 8732
rect 24748 8676 24752 8732
rect 24688 8672 24752 8676
rect 24768 8732 24832 8736
rect 24768 8676 24772 8732
rect 24772 8676 24828 8732
rect 24828 8676 24832 8732
rect 24768 8672 24832 8676
rect 24848 8732 24912 8736
rect 24848 8676 24852 8732
rect 24852 8676 24908 8732
rect 24908 8676 24912 8732
rect 24848 8672 24912 8676
rect 24928 8732 24992 8736
rect 24928 8676 24932 8732
rect 24932 8676 24988 8732
rect 24988 8676 24992 8732
rect 24928 8672 24992 8676
rect 3740 8468 3804 8532
rect 9444 8468 9508 8532
rect 9076 8332 9140 8396
rect 19564 8332 19628 8396
rect 20484 8332 20548 8396
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 9853 8188 9917 8192
rect 9853 8132 9857 8188
rect 9857 8132 9913 8188
rect 9913 8132 9917 8188
rect 9853 8128 9917 8132
rect 9933 8188 9997 8192
rect 9933 8132 9937 8188
rect 9937 8132 9993 8188
rect 9993 8132 9997 8188
rect 9933 8128 9997 8132
rect 10013 8188 10077 8192
rect 10013 8132 10017 8188
rect 10017 8132 10073 8188
rect 10073 8132 10077 8188
rect 10013 8128 10077 8132
rect 10093 8188 10157 8192
rect 10093 8132 10097 8188
rect 10097 8132 10153 8188
rect 10153 8132 10157 8188
rect 10093 8128 10157 8132
rect 15787 8188 15851 8192
rect 15787 8132 15791 8188
rect 15791 8132 15847 8188
rect 15847 8132 15851 8188
rect 15787 8128 15851 8132
rect 15867 8188 15931 8192
rect 15867 8132 15871 8188
rect 15871 8132 15927 8188
rect 15927 8132 15931 8188
rect 15867 8128 15931 8132
rect 15947 8188 16011 8192
rect 15947 8132 15951 8188
rect 15951 8132 16007 8188
rect 16007 8132 16011 8188
rect 15947 8128 16011 8132
rect 16027 8188 16091 8192
rect 16027 8132 16031 8188
rect 16031 8132 16087 8188
rect 16087 8132 16091 8188
rect 16027 8128 16091 8132
rect 21721 8188 21785 8192
rect 21721 8132 21725 8188
rect 21725 8132 21781 8188
rect 21781 8132 21785 8188
rect 21721 8128 21785 8132
rect 21801 8188 21865 8192
rect 21801 8132 21805 8188
rect 21805 8132 21861 8188
rect 21861 8132 21865 8188
rect 21801 8128 21865 8132
rect 21881 8188 21945 8192
rect 21881 8132 21885 8188
rect 21885 8132 21941 8188
rect 21941 8132 21945 8188
rect 21881 8128 21945 8132
rect 21961 8188 22025 8192
rect 21961 8132 21965 8188
rect 21965 8132 22021 8188
rect 22021 8132 22025 8188
rect 21961 8128 22025 8132
rect 2636 7652 2700 7716
rect 15516 7652 15580 7716
rect 6886 7644 6950 7648
rect 6886 7588 6890 7644
rect 6890 7588 6946 7644
rect 6946 7588 6950 7644
rect 6886 7584 6950 7588
rect 6966 7644 7030 7648
rect 6966 7588 6970 7644
rect 6970 7588 7026 7644
rect 7026 7588 7030 7644
rect 6966 7584 7030 7588
rect 7046 7644 7110 7648
rect 7046 7588 7050 7644
rect 7050 7588 7106 7644
rect 7106 7588 7110 7644
rect 7046 7584 7110 7588
rect 7126 7644 7190 7648
rect 7126 7588 7130 7644
rect 7130 7588 7186 7644
rect 7186 7588 7190 7644
rect 7126 7584 7190 7588
rect 12820 7644 12884 7648
rect 12820 7588 12824 7644
rect 12824 7588 12880 7644
rect 12880 7588 12884 7644
rect 12820 7584 12884 7588
rect 12900 7644 12964 7648
rect 12900 7588 12904 7644
rect 12904 7588 12960 7644
rect 12960 7588 12964 7644
rect 12900 7584 12964 7588
rect 12980 7644 13044 7648
rect 12980 7588 12984 7644
rect 12984 7588 13040 7644
rect 13040 7588 13044 7644
rect 12980 7584 13044 7588
rect 13060 7644 13124 7648
rect 13060 7588 13064 7644
rect 13064 7588 13120 7644
rect 13120 7588 13124 7644
rect 13060 7584 13124 7588
rect 18754 7644 18818 7648
rect 18754 7588 18758 7644
rect 18758 7588 18814 7644
rect 18814 7588 18818 7644
rect 18754 7584 18818 7588
rect 18834 7644 18898 7648
rect 18834 7588 18838 7644
rect 18838 7588 18894 7644
rect 18894 7588 18898 7644
rect 18834 7584 18898 7588
rect 18914 7644 18978 7648
rect 18914 7588 18918 7644
rect 18918 7588 18974 7644
rect 18974 7588 18978 7644
rect 18914 7584 18978 7588
rect 18994 7644 19058 7648
rect 18994 7588 18998 7644
rect 18998 7588 19054 7644
rect 19054 7588 19058 7644
rect 18994 7584 19058 7588
rect 24688 7644 24752 7648
rect 24688 7588 24692 7644
rect 24692 7588 24748 7644
rect 24748 7588 24752 7644
rect 24688 7584 24752 7588
rect 24768 7644 24832 7648
rect 24768 7588 24772 7644
rect 24772 7588 24828 7644
rect 24828 7588 24832 7644
rect 24768 7584 24832 7588
rect 24848 7644 24912 7648
rect 24848 7588 24852 7644
rect 24852 7588 24908 7644
rect 24908 7588 24912 7644
rect 24848 7584 24912 7588
rect 24928 7644 24992 7648
rect 24928 7588 24932 7644
rect 24932 7588 24988 7644
rect 24988 7588 24992 7644
rect 24928 7584 24992 7588
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 9853 7100 9917 7104
rect 9853 7044 9857 7100
rect 9857 7044 9913 7100
rect 9913 7044 9917 7100
rect 9853 7040 9917 7044
rect 9933 7100 9997 7104
rect 9933 7044 9937 7100
rect 9937 7044 9993 7100
rect 9993 7044 9997 7100
rect 9933 7040 9997 7044
rect 10013 7100 10077 7104
rect 10013 7044 10017 7100
rect 10017 7044 10073 7100
rect 10073 7044 10077 7100
rect 10013 7040 10077 7044
rect 10093 7100 10157 7104
rect 10093 7044 10097 7100
rect 10097 7044 10153 7100
rect 10153 7044 10157 7100
rect 10093 7040 10157 7044
rect 15787 7100 15851 7104
rect 15787 7044 15791 7100
rect 15791 7044 15847 7100
rect 15847 7044 15851 7100
rect 15787 7040 15851 7044
rect 15867 7100 15931 7104
rect 15867 7044 15871 7100
rect 15871 7044 15927 7100
rect 15927 7044 15931 7100
rect 15867 7040 15931 7044
rect 15947 7100 16011 7104
rect 15947 7044 15951 7100
rect 15951 7044 16007 7100
rect 16007 7044 16011 7100
rect 15947 7040 16011 7044
rect 16027 7100 16091 7104
rect 16027 7044 16031 7100
rect 16031 7044 16087 7100
rect 16087 7044 16091 7100
rect 16027 7040 16091 7044
rect 21721 7100 21785 7104
rect 21721 7044 21725 7100
rect 21725 7044 21781 7100
rect 21781 7044 21785 7100
rect 21721 7040 21785 7044
rect 21801 7100 21865 7104
rect 21801 7044 21805 7100
rect 21805 7044 21861 7100
rect 21861 7044 21865 7100
rect 21801 7040 21865 7044
rect 21881 7100 21945 7104
rect 21881 7044 21885 7100
rect 21885 7044 21941 7100
rect 21941 7044 21945 7100
rect 21881 7040 21945 7044
rect 21961 7100 22025 7104
rect 21961 7044 21965 7100
rect 21965 7044 22021 7100
rect 22021 7044 22025 7100
rect 21961 7040 22025 7044
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 10916 6292 10980 6356
rect 22324 6292 22388 6356
rect 3556 6156 3620 6220
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 4844 5536 4908 5540
rect 4844 5480 4858 5536
rect 4858 5480 4908 5536
rect 4844 5476 4908 5480
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 16988 4856 17052 4860
rect 16988 4800 17038 4856
rect 17038 4800 17052 4856
rect 16988 4796 17052 4800
rect 796 4660 860 4724
rect 612 4388 676 4452
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 980 3980 1044 4044
rect 11652 3980 11716 4044
rect 11836 4040 11900 4044
rect 11836 3984 11850 4040
rect 11850 3984 11900 4040
rect 11836 3980 11900 3984
rect 21588 4040 21652 4044
rect 21588 3984 21638 4040
rect 21638 3984 21652 4040
rect 21588 3980 21652 3984
rect 12204 3844 12268 3908
rect 17356 3844 17420 3908
rect 17724 3904 17788 3908
rect 17724 3848 17738 3904
rect 17738 3848 17788 3904
rect 17724 3844 17788 3848
rect 18092 3844 18156 3908
rect 18460 3904 18524 3908
rect 18460 3848 18510 3904
rect 18510 3848 18524 3904
rect 18460 3844 18524 3848
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 20300 3708 20364 3772
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 22508 3164 22572 3228
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 12572 2620 12636 2684
rect 14044 2620 14108 2684
rect 8340 2484 8404 2548
rect 20300 2484 20364 2548
rect 14412 2348 14476 2412
rect 1164 2212 1228 2276
rect 3740 2212 3804 2276
rect 6500 2212 6564 2276
rect 7972 2272 8036 2276
rect 7972 2216 7986 2272
rect 7986 2216 8036 2272
rect 7972 2212 8036 2216
rect 10916 2212 10980 2276
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 8892 1668 8956 1732
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 1900 1320 1964 1324
rect 1900 1264 1914 1320
rect 1914 1264 1964 1320
rect 1900 1260 1964 1264
rect 2636 1260 2700 1324
rect 5028 1260 5092 1324
rect 6132 1260 6196 1324
rect 9076 1320 9140 1324
rect 9076 1264 9090 1320
rect 9090 1264 9140 1320
rect 9076 1260 9140 1264
rect 19380 1260 19444 1324
rect 20484 1260 20548 1324
rect 23244 1124 23308 1188
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
rect 19932 852 19996 916
<< metal4 >>
rect 18459 44572 18525 44573
rect 18459 44508 18460 44572
rect 18524 44508 18525 44572
rect 18459 44507 18525 44508
rect 3911 43008 4231 43568
rect 3911 42944 3919 43008
rect 3983 42944 3999 43008
rect 4063 42944 4079 43008
rect 4143 42944 4159 43008
rect 4223 42944 4231 43008
rect 1163 42260 1229 42261
rect 1163 42196 1164 42260
rect 1228 42196 1229 42260
rect 1163 42195 1229 42196
rect 979 41444 1045 41445
rect 979 41380 980 41444
rect 1044 41380 1045 41444
rect 979 41379 1045 41380
rect 611 40628 677 40629
rect 611 40564 612 40628
rect 676 40564 677 40628
rect 611 40563 677 40564
rect 614 4453 674 40563
rect 795 40356 861 40357
rect 795 40292 796 40356
rect 860 40292 861 40356
rect 795 40291 861 40292
rect 798 4725 858 40291
rect 795 4724 861 4725
rect 795 4660 796 4724
rect 860 4660 861 4724
rect 795 4659 861 4660
rect 611 4452 677 4453
rect 611 4388 612 4452
rect 676 4388 677 4452
rect 611 4387 677 4388
rect 982 4045 1042 41379
rect 979 4044 1045 4045
rect 979 3980 980 4044
rect 1044 3980 1045 4044
rect 979 3979 1045 3980
rect 1166 2277 1226 42195
rect 3911 41920 4231 42944
rect 3911 41856 3919 41920
rect 3983 41856 3999 41920
rect 4063 41856 4079 41920
rect 4143 41856 4159 41920
rect 4223 41856 4231 41920
rect 3911 40832 4231 41856
rect 6878 43552 7198 43568
rect 6878 43488 6886 43552
rect 6950 43488 6966 43552
rect 7030 43488 7046 43552
rect 7110 43488 7126 43552
rect 7190 43488 7198 43552
rect 6878 42464 7198 43488
rect 6878 42400 6886 42464
rect 6950 42400 6966 42464
rect 7030 42400 7046 42464
rect 7110 42400 7126 42464
rect 7190 42400 7198 42464
rect 6315 41852 6381 41853
rect 6315 41788 6316 41852
rect 6380 41788 6381 41852
rect 6315 41787 6381 41788
rect 3911 40768 3919 40832
rect 3983 40768 3999 40832
rect 4063 40768 4079 40832
rect 4143 40768 4159 40832
rect 4223 40768 4231 40832
rect 2635 40220 2701 40221
rect 2635 40156 2636 40220
rect 2700 40156 2701 40220
rect 2635 40155 2701 40156
rect 2267 39676 2333 39677
rect 2267 39612 2268 39676
rect 2332 39612 2333 39676
rect 2267 39611 2333 39612
rect 2083 38588 2149 38589
rect 2083 38524 2084 38588
rect 2148 38524 2149 38588
rect 2083 38523 2149 38524
rect 1899 30836 1965 30837
rect 1899 30772 1900 30836
rect 1964 30772 1965 30836
rect 1899 30771 1965 30772
rect 1715 27980 1781 27981
rect 1715 27916 1716 27980
rect 1780 27916 1781 27980
rect 1715 27915 1781 27916
rect 1718 18325 1778 27915
rect 1902 26349 1962 30771
rect 2086 30429 2146 38523
rect 2083 30428 2149 30429
rect 2083 30364 2084 30428
rect 2148 30364 2149 30428
rect 2083 30363 2149 30364
rect 2083 28660 2149 28661
rect 2083 28596 2084 28660
rect 2148 28596 2149 28660
rect 2083 28595 2149 28596
rect 1899 26348 1965 26349
rect 1899 26284 1900 26348
rect 1964 26284 1965 26348
rect 1899 26283 1965 26284
rect 2086 18869 2146 28595
rect 2270 26077 2330 39611
rect 2638 32605 2698 40155
rect 3371 40084 3437 40085
rect 3371 40020 3372 40084
rect 3436 40020 3437 40084
rect 3371 40019 3437 40020
rect 3187 37500 3253 37501
rect 3187 37436 3188 37500
rect 3252 37436 3253 37500
rect 3187 37435 3253 37436
rect 2635 32604 2701 32605
rect 2635 32540 2636 32604
rect 2700 32540 2701 32604
rect 2635 32539 2701 32540
rect 3190 32469 3250 37435
rect 3187 32468 3253 32469
rect 3187 32404 3188 32468
rect 3252 32404 3253 32468
rect 3187 32403 3253 32404
rect 2635 30700 2701 30701
rect 2635 30636 2636 30700
rect 2700 30636 2701 30700
rect 2635 30635 2701 30636
rect 2451 28524 2517 28525
rect 2451 28460 2452 28524
rect 2516 28460 2517 28524
rect 2451 28459 2517 28460
rect 2267 26076 2333 26077
rect 2267 26012 2268 26076
rect 2332 26012 2333 26076
rect 2267 26011 2333 26012
rect 2270 22949 2330 26011
rect 2267 22948 2333 22949
rect 2267 22884 2268 22948
rect 2332 22884 2333 22948
rect 2267 22883 2333 22884
rect 2454 22110 2514 28459
rect 2638 25533 2698 30635
rect 2635 25532 2701 25533
rect 2635 25468 2636 25532
rect 2700 25468 2701 25532
rect 2635 25467 2701 25468
rect 2635 24852 2701 24853
rect 2635 24788 2636 24852
rect 2700 24788 2701 24852
rect 2635 24787 2701 24788
rect 2270 22050 2514 22110
rect 2083 18868 2149 18869
rect 2083 18804 2084 18868
rect 2148 18804 2149 18868
rect 2083 18803 2149 18804
rect 1715 18324 1781 18325
rect 1715 18260 1716 18324
rect 1780 18260 1781 18324
rect 1715 18259 1781 18260
rect 2083 16964 2149 16965
rect 2083 16900 2084 16964
rect 2148 16900 2149 16964
rect 2083 16899 2149 16900
rect 2086 10165 2146 16899
rect 2270 13701 2330 22050
rect 2451 20772 2517 20773
rect 2451 20708 2452 20772
rect 2516 20708 2517 20772
rect 2451 20707 2517 20708
rect 2454 16557 2514 20707
rect 2638 19957 2698 24787
rect 3374 23221 3434 40019
rect 3911 39744 4231 40768
rect 3911 39680 3919 39744
rect 3983 39680 3999 39744
rect 4063 39680 4079 39744
rect 4143 39680 4159 39744
rect 4223 39680 4231 39744
rect 3911 38656 4231 39680
rect 4291 38860 4357 38861
rect 4291 38796 4292 38860
rect 4356 38796 4357 38860
rect 4291 38795 4357 38796
rect 3911 38592 3919 38656
rect 3983 38592 3999 38656
rect 4063 38592 4079 38656
rect 4143 38592 4159 38656
rect 4223 38592 4231 38656
rect 3911 37568 4231 38592
rect 3911 37504 3919 37568
rect 3983 37504 3999 37568
rect 4063 37504 4079 37568
rect 4143 37504 4159 37568
rect 4223 37504 4231 37568
rect 3911 36480 4231 37504
rect 3911 36416 3919 36480
rect 3983 36416 3999 36480
rect 4063 36416 4079 36480
rect 4143 36416 4159 36480
rect 4223 36416 4231 36480
rect 3911 35392 4231 36416
rect 4294 35869 4354 38795
rect 5947 37364 6013 37365
rect 5947 37300 5948 37364
rect 6012 37300 6013 37364
rect 5947 37299 6013 37300
rect 5395 37092 5461 37093
rect 5395 37028 5396 37092
rect 5460 37028 5461 37092
rect 5395 37027 5461 37028
rect 5027 36276 5093 36277
rect 5027 36212 5028 36276
rect 5092 36212 5093 36276
rect 5027 36211 5093 36212
rect 4291 35868 4357 35869
rect 4291 35804 4292 35868
rect 4356 35804 4357 35868
rect 4291 35803 4357 35804
rect 3911 35328 3919 35392
rect 3983 35328 3999 35392
rect 4063 35328 4079 35392
rect 4143 35328 4159 35392
rect 4223 35328 4231 35392
rect 3911 34304 4231 35328
rect 3911 34240 3919 34304
rect 3983 34240 3999 34304
rect 4063 34240 4079 34304
rect 4143 34240 4159 34304
rect 4223 34240 4231 34304
rect 3911 33216 4231 34240
rect 3911 33152 3919 33216
rect 3983 33152 3999 33216
rect 4063 33152 4079 33216
rect 4143 33152 4159 33216
rect 4223 33152 4231 33216
rect 3555 32332 3621 32333
rect 3555 32268 3556 32332
rect 3620 32268 3621 32332
rect 3555 32267 3621 32268
rect 3371 23220 3437 23221
rect 3371 23156 3372 23220
rect 3436 23156 3437 23220
rect 3371 23155 3437 23156
rect 3190 20773 3250 21982
rect 3187 20772 3253 20773
rect 3187 20708 3188 20772
rect 3252 20708 3253 20772
rect 3187 20707 3253 20708
rect 2635 19956 2701 19957
rect 2635 19892 2636 19956
rect 2700 19892 2701 19956
rect 2635 19891 2701 19892
rect 2451 16556 2517 16557
rect 2451 16492 2452 16556
rect 2516 16492 2517 16556
rect 2451 16491 2517 16492
rect 3558 16285 3618 32267
rect 3911 32128 4231 33152
rect 4659 32740 4725 32741
rect 4659 32676 4660 32740
rect 4724 32676 4725 32740
rect 4659 32675 4725 32676
rect 3911 32064 3919 32128
rect 3983 32064 3999 32128
rect 4063 32064 4079 32128
rect 4143 32064 4159 32128
rect 4223 32064 4231 32128
rect 3911 31040 4231 32064
rect 4291 31924 4357 31925
rect 4291 31860 4292 31924
rect 4356 31860 4357 31924
rect 4291 31859 4357 31860
rect 3911 30976 3919 31040
rect 3983 30976 3999 31040
rect 4063 30976 4079 31040
rect 4143 30976 4159 31040
rect 4223 30976 4231 31040
rect 3911 29952 4231 30976
rect 3911 29888 3919 29952
rect 3983 29888 3999 29952
rect 4063 29888 4079 29952
rect 4143 29888 4159 29952
rect 4223 29888 4231 29952
rect 3911 28864 4231 29888
rect 4294 29205 4354 31859
rect 4291 29204 4357 29205
rect 4291 29140 4292 29204
rect 4356 29140 4357 29204
rect 4291 29139 4357 29140
rect 3911 28800 3919 28864
rect 3983 28800 3999 28864
rect 4063 28800 4079 28864
rect 4143 28800 4159 28864
rect 4223 28800 4231 28864
rect 3911 27776 4231 28800
rect 4475 28796 4541 28797
rect 4475 28732 4476 28796
rect 4540 28732 4541 28796
rect 4475 28731 4541 28732
rect 3911 27712 3919 27776
rect 3983 27712 3999 27776
rect 4063 27712 4079 27776
rect 4143 27712 4159 27776
rect 4223 27712 4231 27776
rect 3911 26688 4231 27712
rect 3911 26624 3919 26688
rect 3983 26624 3999 26688
rect 4063 26624 4079 26688
rect 4143 26624 4159 26688
rect 4223 26624 4231 26688
rect 3911 25600 4231 26624
rect 3911 25536 3919 25600
rect 3983 25536 3999 25600
rect 4063 25536 4079 25600
rect 4143 25536 4159 25600
rect 4223 25536 4231 25600
rect 3739 24988 3805 24989
rect 3739 24924 3740 24988
rect 3804 24924 3805 24988
rect 3739 24923 3805 24924
rect 3742 20501 3802 24923
rect 3911 24512 4231 25536
rect 4291 24716 4357 24717
rect 4291 24652 4292 24716
rect 4356 24652 4357 24716
rect 4291 24651 4357 24652
rect 3911 24448 3919 24512
rect 3983 24448 3999 24512
rect 4063 24448 4079 24512
rect 4143 24448 4159 24512
rect 4223 24448 4231 24512
rect 3911 23424 4231 24448
rect 3911 23360 3919 23424
rect 3983 23360 3999 23424
rect 4063 23360 4079 23424
rect 4143 23360 4159 23424
rect 4223 23360 4231 23424
rect 3911 22336 4231 23360
rect 3911 22272 3919 22336
rect 3983 22272 3999 22336
rect 4063 22272 4079 22336
rect 4143 22272 4159 22336
rect 4223 22272 4231 22336
rect 3911 21248 4231 22272
rect 3911 21184 3919 21248
rect 3983 21184 3999 21248
rect 4063 21184 4079 21248
rect 4143 21184 4159 21248
rect 4223 21184 4231 21248
rect 3739 20500 3805 20501
rect 3739 20436 3740 20500
rect 3804 20436 3805 20500
rect 3739 20435 3805 20436
rect 3911 20160 4231 21184
rect 3911 20096 3919 20160
rect 3983 20096 3999 20160
rect 4063 20096 4079 20160
rect 4143 20096 4159 20160
rect 4223 20096 4231 20160
rect 3911 19072 4231 20096
rect 4294 19277 4354 24651
rect 4478 24309 4538 28731
rect 4662 28661 4722 32675
rect 5030 29069 5090 36211
rect 5398 31925 5458 37027
rect 5950 35597 6010 37299
rect 5947 35596 6013 35597
rect 5947 35532 5948 35596
rect 6012 35532 6013 35596
rect 5947 35531 6013 35532
rect 5395 31924 5461 31925
rect 5395 31860 5396 31924
rect 5460 31860 5461 31924
rect 5395 31859 5461 31860
rect 5027 29068 5093 29069
rect 5027 29004 5028 29068
rect 5092 29004 5093 29068
rect 5027 29003 5093 29004
rect 4659 28660 4725 28661
rect 4659 28596 4660 28660
rect 4724 28596 4725 28660
rect 4659 28595 4725 28596
rect 4475 24308 4541 24309
rect 4475 24244 4476 24308
rect 4540 24244 4541 24308
rect 4475 24243 4541 24244
rect 4291 19276 4357 19277
rect 4291 19212 4292 19276
rect 4356 19212 4357 19276
rect 4291 19211 4357 19212
rect 3911 19008 3919 19072
rect 3983 19008 3999 19072
rect 4063 19008 4079 19072
rect 4143 19008 4159 19072
rect 4223 19008 4231 19072
rect 3911 17984 4231 19008
rect 4475 18052 4541 18053
rect 4475 17988 4476 18052
rect 4540 17988 4541 18052
rect 4475 17987 4541 17988
rect 3911 17920 3919 17984
rect 3983 17920 3999 17984
rect 4063 17920 4079 17984
rect 4143 17920 4159 17984
rect 4223 17920 4231 17984
rect 3911 16896 4231 17920
rect 3911 16832 3919 16896
rect 3983 16832 3999 16896
rect 4063 16832 4079 16896
rect 4143 16832 4159 16896
rect 4223 16832 4231 16896
rect 3555 16284 3621 16285
rect 3555 16220 3556 16284
rect 3620 16220 3621 16284
rect 3555 16219 3621 16220
rect 2267 13700 2333 13701
rect 2267 13636 2268 13700
rect 2332 13636 2333 13700
rect 2267 13635 2333 13636
rect 3558 13293 3618 16219
rect 3911 15808 4231 16832
rect 3911 15744 3919 15808
rect 3983 15744 3999 15808
rect 4063 15744 4079 15808
rect 4143 15744 4159 15808
rect 4223 15744 4231 15808
rect 3911 14720 4231 15744
rect 3911 14656 3919 14720
rect 3983 14656 3999 14720
rect 4063 14656 4079 14720
rect 4143 14656 4159 14720
rect 4223 14656 4231 14720
rect 3911 13632 4231 14656
rect 3911 13568 3919 13632
rect 3983 13568 3999 13632
rect 4063 13568 4079 13632
rect 4143 13568 4159 13632
rect 4223 13568 4231 13632
rect 3555 13292 3621 13293
rect 3555 13228 3556 13292
rect 3620 13228 3621 13292
rect 3555 13227 3621 13228
rect 3187 12476 3253 12477
rect 3187 12412 3188 12476
rect 3252 12412 3253 12476
rect 3187 12411 3253 12412
rect 3003 10300 3069 10301
rect 3003 10236 3004 10300
rect 3068 10236 3069 10300
rect 3003 10235 3069 10236
rect 2083 10164 2149 10165
rect 2083 10100 2084 10164
rect 2148 10100 2149 10164
rect 2083 10099 2149 10100
rect 1899 9892 1965 9893
rect 1899 9828 1900 9892
rect 1964 9828 1965 9892
rect 1899 9827 1965 9828
rect 1163 2276 1229 2277
rect 1163 2212 1164 2276
rect 1228 2212 1229 2276
rect 1163 2211 1229 2212
rect 1902 1325 1962 9827
rect 3006 9757 3066 10235
rect 3190 9757 3250 12411
rect 3003 9756 3069 9757
rect 3003 9692 3004 9756
rect 3068 9692 3069 9756
rect 3003 9691 3069 9692
rect 3187 9756 3253 9757
rect 3187 9692 3188 9756
rect 3252 9692 3253 9756
rect 3187 9691 3253 9692
rect 2635 7716 2701 7717
rect 2635 7652 2636 7716
rect 2700 7652 2701 7716
rect 2635 7651 2701 7652
rect 2638 1325 2698 7651
rect 3558 6221 3618 13227
rect 3911 12544 4231 13568
rect 3911 12480 3919 12544
rect 3983 12480 3999 12544
rect 4063 12480 4079 12544
rect 4143 12480 4159 12544
rect 4223 12480 4231 12544
rect 3911 11456 4231 12480
rect 3911 11392 3919 11456
rect 3983 11392 3999 11456
rect 4063 11392 4079 11456
rect 4143 11392 4159 11456
rect 4223 11392 4231 11456
rect 3911 10368 4231 11392
rect 4478 10981 4538 17987
rect 4662 15605 4722 28595
rect 5030 21453 5090 29003
rect 5579 23220 5645 23221
rect 5579 23156 5580 23220
rect 5644 23156 5645 23220
rect 5579 23155 5645 23156
rect 5395 22812 5461 22813
rect 5395 22748 5396 22812
rect 5460 22748 5461 22812
rect 5395 22747 5461 22748
rect 5027 21452 5093 21453
rect 5027 21388 5028 21452
rect 5092 21388 5093 21452
rect 5027 21387 5093 21388
rect 5398 17642 5458 22747
rect 5214 17582 5458 17642
rect 5027 16556 5093 16557
rect 5027 16492 5028 16556
rect 5092 16492 5093 16556
rect 5027 16491 5093 16492
rect 4659 15604 4725 15605
rect 4659 15540 4660 15604
rect 4724 15540 4725 15604
rect 4659 15539 4725 15540
rect 4662 12069 4722 15539
rect 4843 13836 4909 13837
rect 4843 13772 4844 13836
rect 4908 13772 4909 13836
rect 4843 13771 4909 13772
rect 4659 12068 4725 12069
rect 4659 12004 4660 12068
rect 4724 12004 4725 12068
rect 4659 12003 4725 12004
rect 4475 10980 4541 10981
rect 4475 10916 4476 10980
rect 4540 10916 4541 10980
rect 4475 10915 4541 10916
rect 3911 10304 3919 10368
rect 3983 10304 3999 10368
rect 4063 10304 4079 10368
rect 4143 10304 4159 10368
rect 4223 10304 4231 10368
rect 3911 9280 4231 10304
rect 3911 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4231 9280
rect 3739 8532 3805 8533
rect 3739 8468 3740 8532
rect 3804 8468 3805 8532
rect 3739 8467 3805 8468
rect 3555 6220 3621 6221
rect 3555 6156 3556 6220
rect 3620 6156 3621 6220
rect 3555 6155 3621 6156
rect 3742 2277 3802 8467
rect 3911 8192 4231 9216
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4231 7104
rect 3911 6016 4231 7040
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 4846 5541 4906 13771
rect 4843 5540 4909 5541
rect 4843 5476 4844 5540
rect 4908 5476 4909 5540
rect 4843 5475 4909 5476
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3739 2276 3805 2277
rect 3739 2212 3740 2276
rect 3804 2212 3805 2276
rect 3739 2211 3805 2212
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 1899 1324 1965 1325
rect 1899 1260 1900 1324
rect 1964 1260 1965 1324
rect 1899 1259 1965 1260
rect 2635 1324 2701 1325
rect 2635 1260 2636 1324
rect 2700 1260 2701 1324
rect 2635 1259 2701 1260
rect 3911 1040 4231 1600
rect 5030 1325 5090 16491
rect 5214 15197 5274 17582
rect 5582 17370 5642 23155
rect 5950 22110 6010 35531
rect 6131 30020 6197 30021
rect 6131 29956 6132 30020
rect 6196 29956 6197 30020
rect 6131 29955 6197 29956
rect 6134 27029 6194 29955
rect 6131 27028 6197 27029
rect 6131 26964 6132 27028
rect 6196 26964 6197 27028
rect 6131 26963 6197 26964
rect 6134 24037 6194 26963
rect 6131 24036 6197 24037
rect 6131 23972 6132 24036
rect 6196 23972 6197 24036
rect 6131 23971 6197 23972
rect 5950 22050 6194 22110
rect 5398 17310 5642 17370
rect 5211 15196 5277 15197
rect 5211 15132 5212 15196
rect 5276 15132 5277 15196
rect 5211 15131 5277 15132
rect 5398 12341 5458 17310
rect 5395 12340 5461 12341
rect 5395 12276 5396 12340
rect 5460 12276 5461 12340
rect 5395 12275 5461 12276
rect 6134 1325 6194 22050
rect 6318 20773 6378 41787
rect 6878 41376 7198 42400
rect 9845 43008 10165 43568
rect 9845 42944 9853 43008
rect 9917 42944 9933 43008
rect 9997 42944 10013 43008
rect 10077 42944 10093 43008
rect 10157 42944 10165 43008
rect 9845 41920 10165 42944
rect 12812 43552 13132 43568
rect 12812 43488 12820 43552
rect 12884 43488 12900 43552
rect 12964 43488 12980 43552
rect 13044 43488 13060 43552
rect 13124 43488 13132 43552
rect 10363 42940 10429 42941
rect 10363 42876 10364 42940
rect 10428 42876 10429 42940
rect 10363 42875 10429 42876
rect 9845 41856 9853 41920
rect 9917 41856 9933 41920
rect 9997 41856 10013 41920
rect 10077 41856 10093 41920
rect 10157 41856 10165 41920
rect 7603 41852 7669 41853
rect 7603 41788 7604 41852
rect 7668 41788 7669 41852
rect 7603 41787 7669 41788
rect 8155 41852 8221 41853
rect 8155 41788 8156 41852
rect 8220 41788 8221 41852
rect 8155 41787 8221 41788
rect 6878 41312 6886 41376
rect 6950 41312 6966 41376
rect 7030 41312 7046 41376
rect 7110 41312 7126 41376
rect 7190 41312 7198 41376
rect 6878 40288 7198 41312
rect 6878 40224 6886 40288
rect 6950 40224 6966 40288
rect 7030 40224 7046 40288
rect 7110 40224 7126 40288
rect 7190 40224 7198 40288
rect 6878 39200 7198 40224
rect 6878 39136 6886 39200
rect 6950 39136 6966 39200
rect 7030 39136 7046 39200
rect 7110 39136 7126 39200
rect 7190 39136 7198 39200
rect 6878 38112 7198 39136
rect 6878 38048 6886 38112
rect 6950 38048 6966 38112
rect 7030 38048 7046 38112
rect 7110 38048 7126 38112
rect 7190 38048 7198 38112
rect 6878 37024 7198 38048
rect 6878 36960 6886 37024
rect 6950 36960 6966 37024
rect 7030 36960 7046 37024
rect 7110 36960 7126 37024
rect 7190 36960 7198 37024
rect 6878 35936 7198 36960
rect 6878 35872 6886 35936
rect 6950 35872 6966 35936
rect 7030 35872 7046 35936
rect 7110 35872 7126 35936
rect 7190 35872 7198 35936
rect 6878 34848 7198 35872
rect 6878 34784 6886 34848
rect 6950 34784 6966 34848
rect 7030 34784 7046 34848
rect 7110 34784 7126 34848
rect 7190 34784 7198 34848
rect 6878 33760 7198 34784
rect 6878 33696 6886 33760
rect 6950 33696 6966 33760
rect 7030 33696 7046 33760
rect 7110 33696 7126 33760
rect 7190 33696 7198 33760
rect 6878 32672 7198 33696
rect 6878 32608 6886 32672
rect 6950 32608 6966 32672
rect 7030 32608 7046 32672
rect 7110 32608 7126 32672
rect 7190 32608 7198 32672
rect 6878 31584 7198 32608
rect 6878 31520 6886 31584
rect 6950 31520 6966 31584
rect 7030 31520 7046 31584
rect 7110 31520 7126 31584
rect 7190 31520 7198 31584
rect 6878 30496 7198 31520
rect 6878 30432 6886 30496
rect 6950 30432 6966 30496
rect 7030 30432 7046 30496
rect 7110 30432 7126 30496
rect 7190 30432 7198 30496
rect 6878 29408 7198 30432
rect 6878 29344 6886 29408
rect 6950 29344 6966 29408
rect 7030 29344 7046 29408
rect 7110 29344 7126 29408
rect 7190 29344 7198 29408
rect 6878 28320 7198 29344
rect 6878 28256 6886 28320
rect 6950 28256 6966 28320
rect 7030 28256 7046 28320
rect 7110 28256 7126 28320
rect 7190 28256 7198 28320
rect 6878 27232 7198 28256
rect 7419 27300 7485 27301
rect 7419 27236 7420 27300
rect 7484 27236 7485 27300
rect 7419 27235 7485 27236
rect 6878 27168 6886 27232
rect 6950 27168 6966 27232
rect 7030 27168 7046 27232
rect 7110 27168 7126 27232
rect 7190 27168 7198 27232
rect 6878 26144 7198 27168
rect 6878 26080 6886 26144
rect 6950 26080 6966 26144
rect 7030 26080 7046 26144
rect 7110 26080 7126 26144
rect 7190 26080 7198 26144
rect 6878 25056 7198 26080
rect 6878 24992 6886 25056
rect 6950 24992 6966 25056
rect 7030 24992 7046 25056
rect 7110 24992 7126 25056
rect 7190 24992 7198 25056
rect 6878 23968 7198 24992
rect 6878 23904 6886 23968
rect 6950 23904 6966 23968
rect 7030 23904 7046 23968
rect 7110 23904 7126 23968
rect 7190 23904 7198 23968
rect 6878 22880 7198 23904
rect 7422 23629 7482 27235
rect 7419 23628 7485 23629
rect 7419 23564 7420 23628
rect 7484 23564 7485 23628
rect 7419 23563 7485 23564
rect 6878 22816 6886 22880
rect 6950 22816 6966 22880
rect 7030 22816 7046 22880
rect 7110 22816 7126 22880
rect 7190 22816 7198 22880
rect 6878 21792 7198 22816
rect 6878 21728 6886 21792
rect 6950 21728 6966 21792
rect 7030 21728 7046 21792
rect 7110 21728 7126 21792
rect 7190 21728 7198 21792
rect 6683 20908 6749 20909
rect 6683 20844 6684 20908
rect 6748 20844 6749 20908
rect 6683 20843 6749 20844
rect 6315 20772 6381 20773
rect 6315 20708 6316 20772
rect 6380 20708 6381 20772
rect 6315 20707 6381 20708
rect 6499 15060 6565 15061
rect 6499 14996 6500 15060
rect 6564 14996 6565 15060
rect 6499 14995 6565 14996
rect 6502 12477 6562 14995
rect 6499 12476 6565 12477
rect 6499 12412 6500 12476
rect 6564 12412 6565 12476
rect 6499 12411 6565 12412
rect 6686 2790 6746 20843
rect 6502 2730 6746 2790
rect 6878 20704 7198 21728
rect 7606 20773 7666 41787
rect 8158 22110 8218 41787
rect 9845 40832 10165 41856
rect 9845 40768 9853 40832
rect 9917 40768 9933 40832
rect 9997 40768 10013 40832
rect 10077 40768 10093 40832
rect 10157 40768 10165 40832
rect 9627 40084 9693 40085
rect 9627 40020 9628 40084
rect 9692 40020 9693 40084
rect 9627 40019 9693 40020
rect 8523 36820 8589 36821
rect 8523 36756 8524 36820
rect 8588 36756 8589 36820
rect 8523 36755 8589 36756
rect 8339 36548 8405 36549
rect 8339 36484 8340 36548
rect 8404 36484 8405 36548
rect 8339 36483 8405 36484
rect 8342 30429 8402 36483
rect 8526 31653 8586 36755
rect 8523 31652 8589 31653
rect 8523 31588 8524 31652
rect 8588 31588 8589 31652
rect 8523 31587 8589 31588
rect 8526 30701 8586 31587
rect 8523 30700 8589 30701
rect 8523 30636 8524 30700
rect 8588 30636 8589 30700
rect 8523 30635 8589 30636
rect 9259 30700 9325 30701
rect 9259 30636 9260 30700
rect 9324 30636 9325 30700
rect 9259 30635 9325 30636
rect 9443 30700 9509 30701
rect 9443 30636 9444 30700
rect 9508 30636 9509 30700
rect 9443 30635 9509 30636
rect 8339 30428 8405 30429
rect 8339 30364 8340 30428
rect 8404 30364 8405 30428
rect 8339 30363 8405 30364
rect 8707 30428 8773 30429
rect 8707 30364 8708 30428
rect 8772 30364 8773 30428
rect 8707 30363 8773 30364
rect 8339 25804 8405 25805
rect 8339 25740 8340 25804
rect 8404 25740 8405 25804
rect 8339 25739 8405 25740
rect 7974 22050 8218 22110
rect 7603 20772 7669 20773
rect 7603 20708 7604 20772
rect 7668 20708 7669 20772
rect 7603 20707 7669 20708
rect 6878 20640 6886 20704
rect 6950 20640 6966 20704
rect 7030 20640 7046 20704
rect 7110 20640 7126 20704
rect 7190 20640 7198 20704
rect 6878 19616 7198 20640
rect 6878 19552 6886 19616
rect 6950 19552 6966 19616
rect 7030 19552 7046 19616
rect 7110 19552 7126 19616
rect 7190 19552 7198 19616
rect 6878 18528 7198 19552
rect 6878 18464 6886 18528
rect 6950 18464 6966 18528
rect 7030 18464 7046 18528
rect 7110 18464 7126 18528
rect 7190 18464 7198 18528
rect 6878 17440 7198 18464
rect 6878 17376 6886 17440
rect 6950 17376 6966 17440
rect 7030 17376 7046 17440
rect 7110 17376 7126 17440
rect 7190 17376 7198 17440
rect 6878 16352 7198 17376
rect 6878 16288 6886 16352
rect 6950 16288 6966 16352
rect 7030 16288 7046 16352
rect 7110 16288 7126 16352
rect 7190 16288 7198 16352
rect 6878 15264 7198 16288
rect 6878 15200 6886 15264
rect 6950 15200 6966 15264
rect 7030 15200 7046 15264
rect 7110 15200 7126 15264
rect 7190 15200 7198 15264
rect 6878 14176 7198 15200
rect 6878 14112 6886 14176
rect 6950 14112 6966 14176
rect 7030 14112 7046 14176
rect 7110 14112 7126 14176
rect 7190 14112 7198 14176
rect 6878 13088 7198 14112
rect 6878 13024 6886 13088
rect 6950 13024 6966 13088
rect 7030 13024 7046 13088
rect 7110 13024 7126 13088
rect 7190 13024 7198 13088
rect 6878 12000 7198 13024
rect 6878 11936 6886 12000
rect 6950 11936 6966 12000
rect 7030 11936 7046 12000
rect 7110 11936 7126 12000
rect 7190 11936 7198 12000
rect 6878 10912 7198 11936
rect 6878 10848 6886 10912
rect 6950 10848 6966 10912
rect 7030 10848 7046 10912
rect 7110 10848 7126 10912
rect 7190 10848 7198 10912
rect 6878 9824 7198 10848
rect 6878 9760 6886 9824
rect 6950 9760 6966 9824
rect 7030 9760 7046 9824
rect 7110 9760 7126 9824
rect 7190 9760 7198 9824
rect 6878 8736 7198 9760
rect 6878 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7198 8736
rect 6878 7648 7198 8672
rect 6878 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7198 7648
rect 6878 6560 7198 7584
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6502 2277 6562 2730
rect 6499 2276 6565 2277
rect 6499 2212 6500 2276
rect 6564 2212 6565 2276
rect 6499 2211 6565 2212
rect 6878 2208 7198 3232
rect 7974 2277 8034 22050
rect 8155 19820 8221 19821
rect 8155 19756 8156 19820
rect 8220 19756 8221 19820
rect 8155 19755 8221 19756
rect 8158 16965 8218 19755
rect 8155 16964 8221 16965
rect 8155 16900 8156 16964
rect 8220 16900 8221 16964
rect 8155 16899 8221 16900
rect 8342 15605 8402 25739
rect 8710 16557 8770 30363
rect 8891 28524 8957 28525
rect 8891 28460 8892 28524
rect 8956 28460 8957 28524
rect 8891 28459 8957 28460
rect 8707 16556 8773 16557
rect 8707 16492 8708 16556
rect 8772 16492 8773 16556
rect 8707 16491 8773 16492
rect 8339 15604 8405 15605
rect 8339 15540 8340 15604
rect 8404 15540 8405 15604
rect 8339 15539 8405 15540
rect 8894 12205 8954 28459
rect 9262 21317 9322 30635
rect 9259 21316 9325 21317
rect 9259 21252 9260 21316
rect 9324 21252 9325 21316
rect 9259 21251 9325 21252
rect 9262 19413 9322 21251
rect 9259 19412 9325 19413
rect 9259 19348 9260 19412
rect 9324 19348 9325 19412
rect 9259 19347 9325 19348
rect 9446 17370 9506 30635
rect 9630 20909 9690 40019
rect 9845 39744 10165 40768
rect 9845 39680 9853 39744
rect 9917 39680 9933 39744
rect 9997 39680 10013 39744
rect 10077 39680 10093 39744
rect 10157 39680 10165 39744
rect 9845 38656 10165 39680
rect 9845 38592 9853 38656
rect 9917 38592 9933 38656
rect 9997 38592 10013 38656
rect 10077 38592 10093 38656
rect 10157 38592 10165 38656
rect 9845 37568 10165 38592
rect 9845 37504 9853 37568
rect 9917 37504 9933 37568
rect 9997 37504 10013 37568
rect 10077 37504 10093 37568
rect 10157 37504 10165 37568
rect 9845 36480 10165 37504
rect 9845 36416 9853 36480
rect 9917 36416 9933 36480
rect 9997 36416 10013 36480
rect 10077 36416 10093 36480
rect 10157 36416 10165 36480
rect 9845 35392 10165 36416
rect 9845 35328 9853 35392
rect 9917 35328 9933 35392
rect 9997 35328 10013 35392
rect 10077 35328 10093 35392
rect 10157 35328 10165 35392
rect 9845 34304 10165 35328
rect 9845 34240 9853 34304
rect 9917 34240 9933 34304
rect 9997 34240 10013 34304
rect 10077 34240 10093 34304
rect 10157 34240 10165 34304
rect 9845 33216 10165 34240
rect 9845 33152 9853 33216
rect 9917 33152 9933 33216
rect 9997 33152 10013 33216
rect 10077 33152 10093 33216
rect 10157 33152 10165 33216
rect 9845 32128 10165 33152
rect 9845 32064 9853 32128
rect 9917 32064 9933 32128
rect 9997 32064 10013 32128
rect 10077 32064 10093 32128
rect 10157 32064 10165 32128
rect 9845 31040 10165 32064
rect 9845 30976 9853 31040
rect 9917 30976 9933 31040
rect 9997 30976 10013 31040
rect 10077 30976 10093 31040
rect 10157 30976 10165 31040
rect 9845 29952 10165 30976
rect 10366 30701 10426 42875
rect 12812 42464 13132 43488
rect 15515 43348 15581 43349
rect 15515 43284 15516 43348
rect 15580 43284 15581 43348
rect 15515 43283 15581 43284
rect 14595 43076 14661 43077
rect 14595 43012 14596 43076
rect 14660 43012 14661 43076
rect 14595 43011 14661 43012
rect 13307 42940 13373 42941
rect 13307 42876 13308 42940
rect 13372 42876 13373 42940
rect 13307 42875 13373 42876
rect 12812 42400 12820 42464
rect 12884 42400 12900 42464
rect 12964 42400 12980 42464
rect 13044 42400 13060 42464
rect 13124 42400 13132 42464
rect 11651 42124 11717 42125
rect 11651 42060 11652 42124
rect 11716 42060 11717 42124
rect 11651 42059 11717 42060
rect 11283 36276 11349 36277
rect 11283 36212 11284 36276
rect 11348 36212 11349 36276
rect 11283 36211 11349 36212
rect 10547 34100 10613 34101
rect 10547 34036 10548 34100
rect 10612 34036 10613 34100
rect 10547 34035 10613 34036
rect 10550 30701 10610 34035
rect 11286 32741 11346 36211
rect 11654 33013 11714 42059
rect 11835 41988 11901 41989
rect 11835 41924 11836 41988
rect 11900 41924 11901 41988
rect 11835 41923 11901 41924
rect 11651 33012 11717 33013
rect 11651 32948 11652 33012
rect 11716 32948 11717 33012
rect 11651 32947 11717 32948
rect 11283 32740 11349 32741
rect 11283 32676 11284 32740
rect 11348 32676 11349 32740
rect 11283 32675 11349 32676
rect 11838 32333 11898 41923
rect 12812 41376 13132 42400
rect 12812 41312 12820 41376
rect 12884 41312 12900 41376
rect 12964 41312 12980 41376
rect 13044 41312 13060 41376
rect 13124 41312 13132 41376
rect 12812 40288 13132 41312
rect 12812 40224 12820 40288
rect 12884 40224 12900 40288
rect 12964 40224 12980 40288
rect 13044 40224 13060 40288
rect 13124 40224 13132 40288
rect 12571 39404 12637 39405
rect 12571 39340 12572 39404
rect 12636 39340 12637 39404
rect 12571 39339 12637 39340
rect 12019 35052 12085 35053
rect 12019 34988 12020 35052
rect 12084 34988 12085 35052
rect 12019 34987 12085 34988
rect 11835 32332 11901 32333
rect 11835 32268 11836 32332
rect 11900 32268 11901 32332
rect 11835 32267 11901 32268
rect 10363 30700 10429 30701
rect 10363 30636 10364 30700
rect 10428 30636 10429 30700
rect 10363 30635 10429 30636
rect 10547 30700 10613 30701
rect 10547 30636 10548 30700
rect 10612 30636 10613 30700
rect 10547 30635 10613 30636
rect 10915 30292 10981 30293
rect 10915 30228 10916 30292
rect 10980 30228 10981 30292
rect 10915 30227 10981 30228
rect 9845 29888 9853 29952
rect 9917 29888 9933 29952
rect 9997 29888 10013 29952
rect 10077 29888 10093 29952
rect 10157 29888 10165 29952
rect 9845 28864 10165 29888
rect 10918 28933 10978 30227
rect 11835 29068 11901 29069
rect 11835 29004 11836 29068
rect 11900 29004 11901 29068
rect 11835 29003 11901 29004
rect 10915 28932 10981 28933
rect 10915 28868 10916 28932
rect 10980 28868 10981 28932
rect 10915 28867 10981 28868
rect 9845 28800 9853 28864
rect 9917 28800 9933 28864
rect 9997 28800 10013 28864
rect 10077 28800 10093 28864
rect 10157 28800 10165 28864
rect 9845 27776 10165 28800
rect 9845 27712 9853 27776
rect 9917 27712 9933 27776
rect 9997 27712 10013 27776
rect 10077 27712 10093 27776
rect 10157 27712 10165 27776
rect 9845 26688 10165 27712
rect 11099 27028 11165 27029
rect 11099 26964 11100 27028
rect 11164 26964 11165 27028
rect 11099 26963 11165 26964
rect 9845 26624 9853 26688
rect 9917 26624 9933 26688
rect 9997 26624 10013 26688
rect 10077 26624 10093 26688
rect 10157 26624 10165 26688
rect 9845 25600 10165 26624
rect 9845 25536 9853 25600
rect 9917 25536 9933 25600
rect 9997 25536 10013 25600
rect 10077 25536 10093 25600
rect 10157 25536 10165 25600
rect 9845 24512 10165 25536
rect 9845 24448 9853 24512
rect 9917 24448 9933 24512
rect 9997 24448 10013 24512
rect 10077 24448 10093 24512
rect 10157 24448 10165 24512
rect 9845 23424 10165 24448
rect 10731 23900 10797 23901
rect 10731 23836 10732 23900
rect 10796 23836 10797 23900
rect 10731 23835 10797 23836
rect 9845 23360 9853 23424
rect 9917 23360 9933 23424
rect 9997 23360 10013 23424
rect 10077 23360 10093 23424
rect 10157 23360 10165 23424
rect 9845 22336 10165 23360
rect 9845 22272 9853 22336
rect 9917 22272 9933 22336
rect 9997 22272 10013 22336
rect 10077 22272 10093 22336
rect 10157 22272 10165 22336
rect 9845 21248 10165 22272
rect 9845 21184 9853 21248
rect 9917 21184 9933 21248
rect 9997 21184 10013 21248
rect 10077 21184 10093 21248
rect 10157 21184 10165 21248
rect 9627 20908 9693 20909
rect 9627 20844 9628 20908
rect 9692 20844 9693 20908
rect 9627 20843 9693 20844
rect 9845 20160 10165 21184
rect 9845 20096 9853 20160
rect 9917 20096 9933 20160
rect 9997 20096 10013 20160
rect 10077 20096 10093 20160
rect 10157 20096 10165 20160
rect 9627 19276 9693 19277
rect 9627 19212 9628 19276
rect 9692 19212 9693 19276
rect 9627 19211 9693 19212
rect 9078 17310 9506 17370
rect 8891 12204 8957 12205
rect 8891 12140 8892 12204
rect 8956 12140 8957 12204
rect 8891 12139 8957 12140
rect 8339 11252 8405 11253
rect 8339 11188 8340 11252
rect 8404 11188 8405 11252
rect 8339 11187 8405 11188
rect 8342 2549 8402 11187
rect 9078 10029 9138 17310
rect 9443 16964 9509 16965
rect 9443 16900 9444 16964
rect 9508 16900 9509 16964
rect 9443 16899 9509 16900
rect 9259 13428 9325 13429
rect 9259 13364 9260 13428
rect 9324 13364 9325 13428
rect 9259 13363 9325 13364
rect 9075 10028 9141 10029
rect 9075 9964 9076 10028
rect 9140 9964 9141 10028
rect 9075 9963 9141 9964
rect 9262 8530 9322 13363
rect 9446 8533 9506 16899
rect 9630 13701 9690 19211
rect 9845 19072 10165 20096
rect 10734 19821 10794 23835
rect 10731 19820 10797 19821
rect 10731 19756 10732 19820
rect 10796 19756 10797 19820
rect 10731 19755 10797 19756
rect 9845 19008 9853 19072
rect 9917 19008 9933 19072
rect 9997 19008 10013 19072
rect 10077 19008 10093 19072
rect 10157 19008 10165 19072
rect 9845 17984 10165 19008
rect 10915 18052 10981 18053
rect 10915 17988 10916 18052
rect 10980 17988 10981 18052
rect 10915 17987 10981 17988
rect 9845 17920 9853 17984
rect 9917 17920 9933 17984
rect 9997 17920 10013 17984
rect 10077 17920 10093 17984
rect 10157 17920 10165 17984
rect 9845 16896 10165 17920
rect 9845 16832 9853 16896
rect 9917 16832 9933 16896
rect 9997 16832 10013 16896
rect 10077 16832 10093 16896
rect 10157 16832 10165 16896
rect 9845 15808 10165 16832
rect 10918 16149 10978 17987
rect 10915 16148 10981 16149
rect 10915 16084 10916 16148
rect 10980 16084 10981 16148
rect 10915 16083 10981 16084
rect 9845 15744 9853 15808
rect 9917 15744 9933 15808
rect 9997 15744 10013 15808
rect 10077 15744 10093 15808
rect 10157 15744 10165 15808
rect 9845 14720 10165 15744
rect 10363 15196 10429 15197
rect 10363 15132 10364 15196
rect 10428 15132 10429 15196
rect 10363 15131 10429 15132
rect 9845 14656 9853 14720
rect 9917 14656 9933 14720
rect 9997 14656 10013 14720
rect 10077 14656 10093 14720
rect 10157 14656 10165 14720
rect 9627 13700 9693 13701
rect 9627 13636 9628 13700
rect 9692 13636 9693 13700
rect 9627 13635 9693 13636
rect 9845 13632 10165 14656
rect 9845 13568 9853 13632
rect 9917 13568 9933 13632
rect 9997 13568 10013 13632
rect 10077 13568 10093 13632
rect 10157 13568 10165 13632
rect 9845 12544 10165 13568
rect 9845 12480 9853 12544
rect 9917 12480 9933 12544
rect 9997 12480 10013 12544
rect 10077 12480 10093 12544
rect 10157 12480 10165 12544
rect 9845 11456 10165 12480
rect 9845 11392 9853 11456
rect 9917 11392 9933 11456
rect 9997 11392 10013 11456
rect 10077 11392 10093 11456
rect 10157 11392 10165 11456
rect 9845 10368 10165 11392
rect 9845 10304 9853 10368
rect 9917 10304 9933 10368
rect 9997 10304 10013 10368
rect 10077 10304 10093 10368
rect 10157 10304 10165 10368
rect 9845 9280 10165 10304
rect 10366 10165 10426 15131
rect 10915 12340 10981 12341
rect 10915 12276 10916 12340
rect 10980 12276 10981 12340
rect 10915 12275 10981 12276
rect 10363 10164 10429 10165
rect 10363 10100 10364 10164
rect 10428 10100 10429 10164
rect 10363 10099 10429 10100
rect 9845 9216 9853 9280
rect 9917 9216 9933 9280
rect 9997 9216 10013 9280
rect 10077 9216 10093 9280
rect 10157 9216 10165 9280
rect 8894 8470 9322 8530
rect 9443 8532 9509 8533
rect 8339 2548 8405 2549
rect 8339 2484 8340 2548
rect 8404 2484 8405 2548
rect 8339 2483 8405 2484
rect 7971 2276 8037 2277
rect 7971 2212 7972 2276
rect 8036 2212 8037 2276
rect 7971 2211 8037 2212
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 5027 1324 5093 1325
rect 5027 1260 5028 1324
rect 5092 1260 5093 1324
rect 5027 1259 5093 1260
rect 6131 1324 6197 1325
rect 6131 1260 6132 1324
rect 6196 1260 6197 1324
rect 6131 1259 6197 1260
rect 6878 1120 7198 2144
rect 8894 1733 8954 8470
rect 9443 8468 9444 8532
rect 9508 8468 9509 8532
rect 9443 8467 9509 8468
rect 9075 8396 9141 8397
rect 9075 8332 9076 8396
rect 9140 8332 9141 8396
rect 9075 8331 9141 8332
rect 8891 1732 8957 1733
rect 8891 1668 8892 1732
rect 8956 1668 8957 1732
rect 8891 1667 8957 1668
rect 9078 1325 9138 8331
rect 9845 8192 10165 9216
rect 9845 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10165 8192
rect 9845 7104 10165 8128
rect 9845 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10165 7104
rect 9845 6016 10165 7040
rect 10918 6357 10978 12275
rect 11102 10573 11162 26963
rect 11651 26212 11717 26213
rect 11651 26148 11652 26212
rect 11716 26148 11717 26212
rect 11651 26147 11717 26148
rect 11467 22540 11533 22541
rect 11467 22476 11468 22540
rect 11532 22476 11533 22540
rect 11467 22475 11533 22476
rect 11099 10572 11165 10573
rect 11099 10508 11100 10572
rect 11164 10508 11165 10572
rect 11099 10507 11165 10508
rect 11470 10029 11530 22475
rect 11467 10028 11533 10029
rect 11467 9964 11468 10028
rect 11532 9964 11533 10028
rect 11467 9963 11533 9964
rect 10915 6356 10981 6357
rect 10915 6292 10916 6356
rect 10980 6292 10981 6356
rect 10915 6291 10981 6292
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9845 1664 10165 2688
rect 10918 2277 10978 6291
rect 11654 4045 11714 26147
rect 11838 4045 11898 29003
rect 12022 26077 12082 34987
rect 12203 34644 12269 34645
rect 12203 34580 12204 34644
rect 12268 34580 12269 34644
rect 12203 34579 12269 34580
rect 12019 26076 12085 26077
rect 12019 26012 12020 26076
rect 12084 26012 12085 26076
rect 12019 26011 12085 26012
rect 12206 25125 12266 34579
rect 12203 25124 12269 25125
rect 12203 25060 12204 25124
rect 12268 25060 12269 25124
rect 12203 25059 12269 25060
rect 12574 22218 12634 39339
rect 12812 39200 13132 40224
rect 12812 39136 12820 39200
rect 12884 39136 12900 39200
rect 12964 39136 12980 39200
rect 13044 39136 13060 39200
rect 13124 39136 13132 39200
rect 12812 38112 13132 39136
rect 12812 38048 12820 38112
rect 12884 38048 12900 38112
rect 12964 38048 12980 38112
rect 13044 38048 13060 38112
rect 13124 38048 13132 38112
rect 12812 37024 13132 38048
rect 12812 36960 12820 37024
rect 12884 36960 12900 37024
rect 12964 36960 12980 37024
rect 13044 36960 13060 37024
rect 13124 36960 13132 37024
rect 12812 35936 13132 36960
rect 12812 35872 12820 35936
rect 12884 35872 12900 35936
rect 12964 35872 12980 35936
rect 13044 35872 13060 35936
rect 13124 35872 13132 35936
rect 12812 34848 13132 35872
rect 12812 34784 12820 34848
rect 12884 34784 12900 34848
rect 12964 34784 12980 34848
rect 13044 34784 13060 34848
rect 13124 34784 13132 34848
rect 12812 33760 13132 34784
rect 12812 33696 12820 33760
rect 12884 33696 12900 33760
rect 12964 33696 12980 33760
rect 13044 33696 13060 33760
rect 13124 33696 13132 33760
rect 12812 32672 13132 33696
rect 12812 32608 12820 32672
rect 12884 32608 12900 32672
rect 12964 32608 12980 32672
rect 13044 32608 13060 32672
rect 13124 32608 13132 32672
rect 12812 31584 13132 32608
rect 12812 31520 12820 31584
rect 12884 31520 12900 31584
rect 12964 31520 12980 31584
rect 13044 31520 13060 31584
rect 13124 31520 13132 31584
rect 12812 30496 13132 31520
rect 12812 30432 12820 30496
rect 12884 30432 12900 30496
rect 12964 30432 12980 30496
rect 13044 30432 13060 30496
rect 13124 30432 13132 30496
rect 12812 29408 13132 30432
rect 12812 29344 12820 29408
rect 12884 29344 12900 29408
rect 12964 29344 12980 29408
rect 13044 29344 13060 29408
rect 13124 29344 13132 29408
rect 12812 28320 13132 29344
rect 12812 28256 12820 28320
rect 12884 28256 12900 28320
rect 12964 28256 12980 28320
rect 13044 28256 13060 28320
rect 13124 28256 13132 28320
rect 12812 27232 13132 28256
rect 12812 27168 12820 27232
rect 12884 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13132 27232
rect 12812 26144 13132 27168
rect 12812 26080 12820 26144
rect 12884 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13132 26144
rect 12812 25056 13132 26080
rect 12812 24992 12820 25056
rect 12884 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13132 25056
rect 12812 23968 13132 24992
rect 12812 23904 12820 23968
rect 12884 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13132 23968
rect 12812 22880 13132 23904
rect 12812 22816 12820 22880
rect 12884 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13132 22880
rect 12812 21792 13132 22816
rect 12812 21728 12820 21792
rect 12884 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13132 21792
rect 12571 20908 12637 20909
rect 12571 20844 12572 20908
rect 12636 20844 12637 20908
rect 12571 20843 12637 20844
rect 12574 17645 12634 20843
rect 12812 20704 13132 21728
rect 12812 20640 12820 20704
rect 12884 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13132 20704
rect 12812 19616 13132 20640
rect 12812 19552 12820 19616
rect 12884 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13132 19616
rect 12812 18528 13132 19552
rect 12812 18464 12820 18528
rect 12884 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13132 18528
rect 12571 17644 12637 17645
rect 12571 17580 12572 17644
rect 12636 17580 12637 17644
rect 12571 17579 12637 17580
rect 12812 17440 13132 18464
rect 12812 17376 12820 17440
rect 12884 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13132 17440
rect 12571 16692 12637 16693
rect 12571 16628 12572 16692
rect 12636 16628 12637 16692
rect 12571 16627 12637 16628
rect 12203 9756 12269 9757
rect 12203 9692 12204 9756
rect 12268 9692 12269 9756
rect 12203 9691 12269 9692
rect 11651 4044 11717 4045
rect 11651 3980 11652 4044
rect 11716 3980 11717 4044
rect 11651 3979 11717 3980
rect 11835 4044 11901 4045
rect 11835 3980 11836 4044
rect 11900 3980 11901 4044
rect 11835 3979 11901 3980
rect 12206 3909 12266 9691
rect 12203 3908 12269 3909
rect 12203 3844 12204 3908
rect 12268 3844 12269 3908
rect 12203 3843 12269 3844
rect 12574 2685 12634 16627
rect 12812 16352 13132 17376
rect 12812 16288 12820 16352
rect 12884 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13132 16352
rect 12812 15264 13132 16288
rect 13310 15469 13370 42875
rect 13859 38316 13925 38317
rect 13859 38252 13860 38316
rect 13924 38252 13925 38316
rect 13859 38251 13925 38252
rect 13491 35460 13557 35461
rect 13491 35396 13492 35460
rect 13556 35396 13557 35460
rect 13491 35395 13557 35396
rect 13494 31109 13554 35395
rect 13491 31108 13557 31109
rect 13491 31044 13492 31108
rect 13556 31044 13557 31108
rect 13491 31043 13557 31044
rect 13675 28524 13741 28525
rect 13675 28460 13676 28524
rect 13740 28460 13741 28524
rect 13675 28459 13741 28460
rect 13678 19821 13738 28459
rect 13862 21997 13922 38251
rect 14227 30836 14293 30837
rect 14227 30772 14228 30836
rect 14292 30772 14293 30836
rect 14227 30771 14293 30772
rect 14230 25125 14290 30771
rect 14227 25124 14293 25125
rect 14227 25060 14228 25124
rect 14292 25060 14293 25124
rect 14227 25059 14293 25060
rect 13859 21996 13925 21997
rect 13859 21932 13860 21996
rect 13924 21932 13925 21996
rect 13859 21931 13925 21932
rect 13675 19820 13741 19821
rect 13675 19756 13676 19820
rect 13740 19756 13741 19820
rect 13675 19755 13741 19756
rect 14411 18732 14477 18733
rect 14411 18668 14412 18732
rect 14476 18668 14477 18732
rect 14411 18667 14477 18668
rect 14043 16012 14109 16013
rect 14043 15948 14044 16012
rect 14108 15948 14109 16012
rect 14043 15947 14109 15948
rect 13307 15468 13373 15469
rect 13307 15404 13308 15468
rect 13372 15404 13373 15468
rect 13307 15403 13373 15404
rect 12812 15200 12820 15264
rect 12884 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13132 15264
rect 12812 14176 13132 15200
rect 12812 14112 12820 14176
rect 12884 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13132 14176
rect 12812 13088 13132 14112
rect 12812 13024 12820 13088
rect 12884 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13132 13088
rect 12812 12000 13132 13024
rect 12812 11936 12820 12000
rect 12884 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13132 12000
rect 12812 10912 13132 11936
rect 12812 10848 12820 10912
rect 12884 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13132 10912
rect 12812 9824 13132 10848
rect 12812 9760 12820 9824
rect 12884 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13132 9824
rect 12812 8736 13132 9760
rect 12812 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13132 8736
rect 12812 7648 13132 8672
rect 12812 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13132 7648
rect 12812 6560 13132 7584
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12571 2684 12637 2685
rect 12571 2620 12572 2684
rect 12636 2620 12637 2684
rect 12571 2619 12637 2620
rect 10915 2276 10981 2277
rect 10915 2212 10916 2276
rect 10980 2212 10981 2276
rect 10915 2211 10981 2212
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9075 1324 9141 1325
rect 9075 1260 9076 1324
rect 9140 1260 9141 1324
rect 9075 1259 9141 1260
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 1040 10165 1600
rect 12812 2208 13132 3232
rect 14046 2685 14106 15947
rect 14043 2684 14109 2685
rect 14043 2620 14044 2684
rect 14108 2620 14109 2684
rect 14043 2619 14109 2620
rect 14414 2413 14474 18667
rect 14598 9893 14658 43011
rect 14963 42940 15029 42941
rect 14963 42876 14964 42940
rect 15028 42876 15029 42940
rect 14963 42875 15029 42876
rect 14966 19957 15026 42875
rect 15331 27436 15397 27437
rect 15331 27372 15332 27436
rect 15396 27372 15397 27436
rect 15331 27371 15397 27372
rect 15334 24581 15394 27371
rect 15518 26893 15578 43283
rect 15779 43008 16099 43568
rect 15779 42944 15787 43008
rect 15851 42944 15867 43008
rect 15931 42944 15947 43008
rect 16011 42944 16027 43008
rect 16091 42944 16099 43008
rect 15779 41920 16099 42944
rect 18462 42261 18522 44507
rect 18746 43552 19066 43568
rect 18746 43488 18754 43552
rect 18818 43488 18834 43552
rect 18898 43488 18914 43552
rect 18978 43488 18994 43552
rect 19058 43488 19066 43552
rect 18746 42464 19066 43488
rect 21587 43212 21653 43213
rect 21587 43148 21588 43212
rect 21652 43148 21653 43212
rect 21587 43147 21653 43148
rect 18746 42400 18754 42464
rect 18818 42400 18834 42464
rect 18898 42400 18914 42464
rect 18978 42400 18994 42464
rect 19058 42400 19066 42464
rect 18459 42260 18525 42261
rect 18459 42196 18460 42260
rect 18524 42196 18525 42260
rect 18459 42195 18525 42196
rect 15779 41856 15787 41920
rect 15851 41856 15867 41920
rect 15931 41856 15947 41920
rect 16011 41856 16027 41920
rect 16091 41856 16099 41920
rect 15779 40832 16099 41856
rect 16987 41716 17053 41717
rect 16987 41652 16988 41716
rect 17052 41652 17053 41716
rect 16987 41651 17053 41652
rect 17723 41716 17789 41717
rect 17723 41652 17724 41716
rect 17788 41652 17789 41716
rect 17723 41651 17789 41652
rect 18275 41716 18341 41717
rect 18275 41652 18276 41716
rect 18340 41652 18341 41716
rect 18275 41651 18341 41652
rect 15779 40768 15787 40832
rect 15851 40768 15867 40832
rect 15931 40768 15947 40832
rect 16011 40768 16027 40832
rect 16091 40768 16099 40832
rect 15779 39744 16099 40768
rect 15779 39680 15787 39744
rect 15851 39680 15867 39744
rect 15931 39680 15947 39744
rect 16011 39680 16027 39744
rect 16091 39680 16099 39744
rect 15779 38656 16099 39680
rect 16435 39540 16501 39541
rect 16435 39476 16436 39540
rect 16500 39476 16501 39540
rect 16435 39475 16501 39476
rect 15779 38592 15787 38656
rect 15851 38592 15867 38656
rect 15931 38592 15947 38656
rect 16011 38592 16027 38656
rect 16091 38592 16099 38656
rect 15779 37568 16099 38592
rect 15779 37504 15787 37568
rect 15851 37504 15867 37568
rect 15931 37504 15947 37568
rect 16011 37504 16027 37568
rect 16091 37504 16099 37568
rect 15779 36480 16099 37504
rect 15779 36416 15787 36480
rect 15851 36416 15867 36480
rect 15931 36416 15947 36480
rect 16011 36416 16027 36480
rect 16091 36416 16099 36480
rect 15779 35392 16099 36416
rect 15779 35328 15787 35392
rect 15851 35328 15867 35392
rect 15931 35328 15947 35392
rect 16011 35328 16027 35392
rect 16091 35328 16099 35392
rect 15779 34304 16099 35328
rect 15779 34240 15787 34304
rect 15851 34240 15867 34304
rect 15931 34240 15947 34304
rect 16011 34240 16027 34304
rect 16091 34240 16099 34304
rect 15779 33216 16099 34240
rect 15779 33152 15787 33216
rect 15851 33152 15867 33216
rect 15931 33152 15947 33216
rect 16011 33152 16027 33216
rect 16091 33152 16099 33216
rect 15779 32128 16099 33152
rect 15779 32064 15787 32128
rect 15851 32064 15867 32128
rect 15931 32064 15947 32128
rect 16011 32064 16027 32128
rect 16091 32064 16099 32128
rect 15779 31040 16099 32064
rect 15779 30976 15787 31040
rect 15851 30976 15867 31040
rect 15931 30976 15947 31040
rect 16011 30976 16027 31040
rect 16091 30976 16099 31040
rect 15779 29952 16099 30976
rect 15779 29888 15787 29952
rect 15851 29888 15867 29952
rect 15931 29888 15947 29952
rect 16011 29888 16027 29952
rect 16091 29888 16099 29952
rect 15779 28864 16099 29888
rect 15779 28800 15787 28864
rect 15851 28800 15867 28864
rect 15931 28800 15947 28864
rect 16011 28800 16027 28864
rect 16091 28800 16099 28864
rect 15779 27776 16099 28800
rect 15779 27712 15787 27776
rect 15851 27712 15867 27776
rect 15931 27712 15947 27776
rect 16011 27712 16027 27776
rect 16091 27712 16099 27776
rect 15515 26892 15581 26893
rect 15515 26828 15516 26892
rect 15580 26828 15581 26892
rect 15515 26827 15581 26828
rect 15779 26688 16099 27712
rect 16438 27301 16498 39475
rect 16990 30837 17050 41651
rect 16987 30836 17053 30837
rect 16987 30772 16988 30836
rect 17052 30772 17053 30836
rect 16987 30771 17053 30772
rect 16987 30700 17053 30701
rect 16987 30636 16988 30700
rect 17052 30636 17053 30700
rect 16987 30635 17053 30636
rect 16619 29476 16685 29477
rect 16619 29412 16620 29476
rect 16684 29412 16685 29476
rect 16619 29411 16685 29412
rect 16435 27300 16501 27301
rect 16435 27236 16436 27300
rect 16500 27236 16501 27300
rect 16435 27235 16501 27236
rect 15779 26624 15787 26688
rect 15851 26624 15867 26688
rect 15931 26624 15947 26688
rect 16011 26624 16027 26688
rect 16091 26624 16099 26688
rect 15779 25600 16099 26624
rect 16251 25940 16317 25941
rect 16251 25876 16252 25940
rect 16316 25876 16317 25940
rect 16251 25875 16317 25876
rect 15779 25536 15787 25600
rect 15851 25536 15867 25600
rect 15931 25536 15947 25600
rect 16011 25536 16027 25600
rect 16091 25536 16099 25600
rect 15331 24580 15397 24581
rect 15331 24516 15332 24580
rect 15396 24516 15397 24580
rect 15331 24515 15397 24516
rect 15334 24170 15394 24515
rect 15150 24110 15394 24170
rect 15779 24512 16099 25536
rect 15779 24448 15787 24512
rect 15851 24448 15867 24512
rect 15931 24448 15947 24512
rect 16011 24448 16027 24512
rect 16091 24448 16099 24512
rect 14963 19956 15029 19957
rect 14963 19892 14964 19956
rect 15028 19892 15029 19956
rect 14963 19891 15029 19892
rect 15150 19549 15210 24110
rect 15779 23424 16099 24448
rect 15779 23360 15787 23424
rect 15851 23360 15867 23424
rect 15931 23360 15947 23424
rect 16011 23360 16027 23424
rect 16091 23360 16099 23424
rect 15779 22336 16099 23360
rect 15779 22272 15787 22336
rect 15851 22272 15867 22336
rect 15931 22272 15947 22336
rect 16011 22272 16027 22336
rect 16091 22272 16099 22336
rect 15779 21248 16099 22272
rect 15779 21184 15787 21248
rect 15851 21184 15867 21248
rect 15931 21184 15947 21248
rect 16011 21184 16027 21248
rect 16091 21184 16099 21248
rect 15779 20160 16099 21184
rect 15779 20096 15787 20160
rect 15851 20096 15867 20160
rect 15931 20096 15947 20160
rect 16011 20096 16027 20160
rect 16091 20096 16099 20160
rect 15147 19548 15213 19549
rect 15147 19484 15148 19548
rect 15212 19484 15213 19548
rect 15147 19483 15213 19484
rect 15150 16693 15210 19483
rect 15779 19072 16099 20096
rect 15779 19008 15787 19072
rect 15851 19008 15867 19072
rect 15931 19008 15947 19072
rect 16011 19008 16027 19072
rect 16091 19008 16099 19072
rect 15331 18732 15397 18733
rect 15331 18668 15332 18732
rect 15396 18668 15397 18732
rect 15331 18667 15397 18668
rect 15147 16692 15213 16693
rect 15147 16628 15148 16692
rect 15212 16628 15213 16692
rect 15147 16627 15213 16628
rect 15334 11933 15394 18667
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 15331 11932 15397 11933
rect 15331 11868 15332 11932
rect 15396 11868 15397 11932
rect 15331 11867 15397 11868
rect 14595 9892 14661 9893
rect 14595 9828 14596 9892
rect 14660 9828 14661 9892
rect 14595 9827 14661 9828
rect 15334 9077 15394 11867
rect 15331 9076 15397 9077
rect 15331 9012 15332 9076
rect 15396 9012 15397 9076
rect 15331 9011 15397 9012
rect 15518 7717 15578 17987
rect 15779 17984 16099 19008
rect 15779 17920 15787 17984
rect 15851 17920 15867 17984
rect 15931 17920 15947 17984
rect 16011 17920 16027 17984
rect 16091 17920 16099 17984
rect 15779 16896 16099 17920
rect 16254 17917 16314 25875
rect 16622 24989 16682 29411
rect 16619 24988 16685 24989
rect 16619 24924 16620 24988
rect 16684 24924 16685 24988
rect 16619 24923 16685 24924
rect 16435 24308 16501 24309
rect 16435 24244 16436 24308
rect 16500 24244 16501 24308
rect 16435 24243 16501 24244
rect 16438 21317 16498 24243
rect 16619 21452 16685 21453
rect 16619 21388 16620 21452
rect 16684 21388 16685 21452
rect 16619 21387 16685 21388
rect 16435 21316 16501 21317
rect 16435 21252 16436 21316
rect 16500 21252 16501 21316
rect 16435 21251 16501 21252
rect 16438 18733 16498 21251
rect 16435 18732 16501 18733
rect 16435 18668 16436 18732
rect 16500 18668 16501 18732
rect 16435 18667 16501 18668
rect 16251 17916 16317 17917
rect 16251 17852 16252 17916
rect 16316 17852 16317 17916
rect 16251 17851 16317 17852
rect 16622 17237 16682 21387
rect 16803 19412 16869 19413
rect 16803 19348 16804 19412
rect 16868 19348 16869 19412
rect 16803 19347 16869 19348
rect 16619 17236 16685 17237
rect 16619 17172 16620 17236
rect 16684 17172 16685 17236
rect 16619 17171 16685 17172
rect 15779 16832 15787 16896
rect 15851 16832 15867 16896
rect 15931 16832 15947 16896
rect 16011 16832 16027 16896
rect 16091 16832 16099 16896
rect 15779 15808 16099 16832
rect 15779 15744 15787 15808
rect 15851 15744 15867 15808
rect 15931 15744 15947 15808
rect 16011 15744 16027 15808
rect 16091 15744 16099 15808
rect 15779 14720 16099 15744
rect 15779 14656 15787 14720
rect 15851 14656 15867 14720
rect 15931 14656 15947 14720
rect 16011 14656 16027 14720
rect 16091 14656 16099 14720
rect 15779 13632 16099 14656
rect 15779 13568 15787 13632
rect 15851 13568 15867 13632
rect 15931 13568 15947 13632
rect 16011 13568 16027 13632
rect 16091 13568 16099 13632
rect 15779 12544 16099 13568
rect 15779 12480 15787 12544
rect 15851 12480 15867 12544
rect 15931 12480 15947 12544
rect 16011 12480 16027 12544
rect 16091 12480 16099 12544
rect 15779 11456 16099 12480
rect 15779 11392 15787 11456
rect 15851 11392 15867 11456
rect 15931 11392 15947 11456
rect 16011 11392 16027 11456
rect 16091 11392 16099 11456
rect 15779 10368 16099 11392
rect 15779 10304 15787 10368
rect 15851 10304 15867 10368
rect 15931 10304 15947 10368
rect 16011 10304 16027 10368
rect 16091 10304 16099 10368
rect 15779 9280 16099 10304
rect 16806 9757 16866 19347
rect 16990 19277 17050 30635
rect 17726 29749 17786 41651
rect 18278 35869 18338 41651
rect 18459 41444 18525 41445
rect 18459 41380 18460 41444
rect 18524 41380 18525 41444
rect 18459 41379 18525 41380
rect 18275 35868 18341 35869
rect 18275 35804 18276 35868
rect 18340 35804 18341 35868
rect 18275 35803 18341 35804
rect 18091 33148 18157 33149
rect 18091 33084 18092 33148
rect 18156 33084 18157 33148
rect 18091 33083 18157 33084
rect 17723 29748 17789 29749
rect 17723 29684 17724 29748
rect 17788 29684 17789 29748
rect 17723 29683 17789 29684
rect 17539 27708 17605 27709
rect 17539 27644 17540 27708
rect 17604 27644 17605 27708
rect 17539 27643 17605 27644
rect 17355 26756 17421 26757
rect 17355 26692 17356 26756
rect 17420 26692 17421 26756
rect 17355 26691 17421 26692
rect 17171 25668 17237 25669
rect 17171 25604 17172 25668
rect 17236 25604 17237 25668
rect 17171 25603 17237 25604
rect 17174 21861 17234 25603
rect 17171 21860 17237 21861
rect 17171 21796 17172 21860
rect 17236 21796 17237 21860
rect 17171 21795 17237 21796
rect 17358 21181 17418 26691
rect 17542 25261 17602 27643
rect 17539 25260 17605 25261
rect 17539 25196 17540 25260
rect 17604 25196 17605 25260
rect 17539 25195 17605 25196
rect 17542 21589 17602 25195
rect 17723 24172 17789 24173
rect 17723 24108 17724 24172
rect 17788 24108 17789 24172
rect 17723 24107 17789 24108
rect 17539 21588 17605 21589
rect 17539 21524 17540 21588
rect 17604 21524 17605 21588
rect 17539 21523 17605 21524
rect 17355 21180 17421 21181
rect 17355 21116 17356 21180
rect 17420 21116 17421 21180
rect 17355 21115 17421 21116
rect 16987 19276 17053 19277
rect 16987 19212 16988 19276
rect 17052 19212 17053 19276
rect 16987 19211 17053 19212
rect 17171 18868 17237 18869
rect 17171 18804 17172 18868
rect 17236 18804 17237 18868
rect 17171 18803 17237 18804
rect 16987 17236 17053 17237
rect 16987 17172 16988 17236
rect 17052 17172 17053 17236
rect 16987 17171 17053 17172
rect 16803 9756 16869 9757
rect 16803 9692 16804 9756
rect 16868 9692 16869 9756
rect 16803 9691 16869 9692
rect 15779 9216 15787 9280
rect 15851 9216 15867 9280
rect 15931 9216 15947 9280
rect 16011 9216 16027 9280
rect 16091 9216 16099 9280
rect 15779 8192 16099 9216
rect 15779 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16099 8192
rect 15515 7716 15581 7717
rect 15515 7652 15516 7716
rect 15580 7652 15581 7716
rect 15515 7651 15581 7652
rect 15779 7104 16099 8128
rect 15779 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16099 7104
rect 15779 6016 16099 7040
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15779 3840 16099 4864
rect 16990 4861 17050 17171
rect 17174 16149 17234 18803
rect 17171 16148 17237 16149
rect 17171 16084 17172 16148
rect 17236 16084 17237 16148
rect 17171 16083 17237 16084
rect 17355 15468 17421 15469
rect 17355 15404 17356 15468
rect 17420 15404 17421 15468
rect 17355 15403 17421 15404
rect 16987 4860 17053 4861
rect 16987 4796 16988 4860
rect 17052 4796 17053 4860
rect 16987 4795 17053 4796
rect 17358 3909 17418 15403
rect 17726 3909 17786 24107
rect 18094 3909 18154 33083
rect 18462 3909 18522 41379
rect 18746 41376 19066 42400
rect 20667 42124 20733 42125
rect 20667 42060 20668 42124
rect 20732 42060 20733 42124
rect 20667 42059 20733 42060
rect 19563 41716 19629 41717
rect 19563 41652 19564 41716
rect 19628 41652 19629 41716
rect 19563 41651 19629 41652
rect 18746 41312 18754 41376
rect 18818 41312 18834 41376
rect 18898 41312 18914 41376
rect 18978 41312 18994 41376
rect 19058 41312 19066 41376
rect 18746 40288 19066 41312
rect 18746 40224 18754 40288
rect 18818 40224 18834 40288
rect 18898 40224 18914 40288
rect 18978 40224 18994 40288
rect 19058 40224 19066 40288
rect 18746 39200 19066 40224
rect 18746 39136 18754 39200
rect 18818 39136 18834 39200
rect 18898 39136 18914 39200
rect 18978 39136 18994 39200
rect 19058 39136 19066 39200
rect 18746 38112 19066 39136
rect 18746 38048 18754 38112
rect 18818 38048 18834 38112
rect 18898 38048 18914 38112
rect 18978 38048 18994 38112
rect 19058 38048 19066 38112
rect 18746 37024 19066 38048
rect 18746 36960 18754 37024
rect 18818 36960 18834 37024
rect 18898 36960 18914 37024
rect 18978 36960 18994 37024
rect 19058 36960 19066 37024
rect 18746 35936 19066 36960
rect 18746 35872 18754 35936
rect 18818 35872 18834 35936
rect 18898 35872 18914 35936
rect 18978 35872 18994 35936
rect 19058 35872 19066 35936
rect 18746 34848 19066 35872
rect 18746 34784 18754 34848
rect 18818 34784 18834 34848
rect 18898 34784 18914 34848
rect 18978 34784 18994 34848
rect 19058 34784 19066 34848
rect 18746 33760 19066 34784
rect 18746 33696 18754 33760
rect 18818 33696 18834 33760
rect 18898 33696 18914 33760
rect 18978 33696 18994 33760
rect 19058 33696 19066 33760
rect 18746 32672 19066 33696
rect 18746 32608 18754 32672
rect 18818 32608 18834 32672
rect 18898 32608 18914 32672
rect 18978 32608 18994 32672
rect 19058 32608 19066 32672
rect 18746 31584 19066 32608
rect 18746 31520 18754 31584
rect 18818 31520 18834 31584
rect 18898 31520 18914 31584
rect 18978 31520 18994 31584
rect 19058 31520 19066 31584
rect 18746 30496 19066 31520
rect 18746 30432 18754 30496
rect 18818 30432 18834 30496
rect 18898 30432 18914 30496
rect 18978 30432 18994 30496
rect 19058 30432 19066 30496
rect 18746 29408 19066 30432
rect 18746 29344 18754 29408
rect 18818 29344 18834 29408
rect 18898 29344 18914 29408
rect 18978 29344 18994 29408
rect 19058 29344 19066 29408
rect 18746 28320 19066 29344
rect 18746 28256 18754 28320
rect 18818 28256 18834 28320
rect 18898 28256 18914 28320
rect 18978 28256 18994 28320
rect 19058 28256 19066 28320
rect 18746 27232 19066 28256
rect 18746 27168 18754 27232
rect 18818 27168 18834 27232
rect 18898 27168 18914 27232
rect 18978 27168 18994 27232
rect 19058 27168 19066 27232
rect 18746 26144 19066 27168
rect 18746 26080 18754 26144
rect 18818 26080 18834 26144
rect 18898 26080 18914 26144
rect 18978 26080 18994 26144
rect 19058 26080 19066 26144
rect 18746 25056 19066 26080
rect 18746 24992 18754 25056
rect 18818 24992 18834 25056
rect 18898 24992 18914 25056
rect 18978 24992 18994 25056
rect 19058 24992 19066 25056
rect 18746 23968 19066 24992
rect 18746 23904 18754 23968
rect 18818 23904 18834 23968
rect 18898 23904 18914 23968
rect 18978 23904 18994 23968
rect 19058 23904 19066 23968
rect 18746 22880 19066 23904
rect 18746 22816 18754 22880
rect 18818 22816 18834 22880
rect 18898 22816 18914 22880
rect 18978 22816 18994 22880
rect 19058 22816 19066 22880
rect 18746 21792 19066 22816
rect 19566 22110 19626 41651
rect 19747 38860 19813 38861
rect 19747 38796 19748 38860
rect 19812 38796 19813 38860
rect 19747 38795 19813 38796
rect 18746 21728 18754 21792
rect 18818 21728 18834 21792
rect 18898 21728 18914 21792
rect 18978 21728 18994 21792
rect 19058 21728 19066 21792
rect 18746 20704 19066 21728
rect 19382 22050 19626 22110
rect 19382 20773 19442 22050
rect 19563 21180 19629 21181
rect 19563 21116 19564 21180
rect 19628 21116 19629 21180
rect 19563 21115 19629 21116
rect 19379 20772 19445 20773
rect 19379 20708 19380 20772
rect 19444 20708 19445 20772
rect 19379 20707 19445 20708
rect 18746 20640 18754 20704
rect 18818 20640 18834 20704
rect 18898 20640 18914 20704
rect 18978 20640 18994 20704
rect 19058 20640 19066 20704
rect 18746 19616 19066 20640
rect 18746 19552 18754 19616
rect 18818 19552 18834 19616
rect 18898 19552 18914 19616
rect 18978 19552 18994 19616
rect 19058 19552 19066 19616
rect 18746 18528 19066 19552
rect 18746 18464 18754 18528
rect 18818 18464 18834 18528
rect 18898 18464 18914 18528
rect 18978 18464 18994 18528
rect 19058 18464 19066 18528
rect 18746 17440 19066 18464
rect 18746 17376 18754 17440
rect 18818 17376 18834 17440
rect 18898 17376 18914 17440
rect 18978 17376 18994 17440
rect 19058 17376 19066 17440
rect 18746 16352 19066 17376
rect 19379 16556 19445 16557
rect 19379 16492 19380 16556
rect 19444 16492 19445 16556
rect 19379 16491 19445 16492
rect 18746 16288 18754 16352
rect 18818 16288 18834 16352
rect 18898 16288 18914 16352
rect 18978 16288 18994 16352
rect 19058 16288 19066 16352
rect 18746 15264 19066 16288
rect 18746 15200 18754 15264
rect 18818 15200 18834 15264
rect 18898 15200 18914 15264
rect 18978 15200 18994 15264
rect 19058 15200 19066 15264
rect 18746 14176 19066 15200
rect 18746 14112 18754 14176
rect 18818 14112 18834 14176
rect 18898 14112 18914 14176
rect 18978 14112 18994 14176
rect 19058 14112 19066 14176
rect 18746 13088 19066 14112
rect 18746 13024 18754 13088
rect 18818 13024 18834 13088
rect 18898 13024 18914 13088
rect 18978 13024 18994 13088
rect 19058 13024 19066 13088
rect 18746 12000 19066 13024
rect 18746 11936 18754 12000
rect 18818 11936 18834 12000
rect 18898 11936 18914 12000
rect 18978 11936 18994 12000
rect 19058 11936 19066 12000
rect 18746 10912 19066 11936
rect 18746 10848 18754 10912
rect 18818 10848 18834 10912
rect 18898 10848 18914 10912
rect 18978 10848 18994 10912
rect 19058 10848 19066 10912
rect 18746 9824 19066 10848
rect 18746 9760 18754 9824
rect 18818 9760 18834 9824
rect 18898 9760 18914 9824
rect 18978 9760 18994 9824
rect 19058 9760 19066 9824
rect 18746 8736 19066 9760
rect 18746 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19066 8736
rect 18746 7648 19066 8672
rect 18746 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19066 7648
rect 18746 6560 19066 7584
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 17355 3908 17421 3909
rect 17355 3844 17356 3908
rect 17420 3844 17421 3908
rect 17355 3843 17421 3844
rect 17723 3908 17789 3909
rect 17723 3844 17724 3908
rect 17788 3844 17789 3908
rect 17723 3843 17789 3844
rect 18091 3908 18157 3909
rect 18091 3844 18092 3908
rect 18156 3844 18157 3908
rect 18091 3843 18157 3844
rect 18459 3908 18525 3909
rect 18459 3844 18460 3908
rect 18524 3844 18525 3908
rect 18459 3843 18525 3844
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 14411 2412 14477 2413
rect 14411 2348 14412 2412
rect 14476 2348 14477 2412
rect 14411 2347 14477 2348
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 1664 16099 2688
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 18746 3296 19066 4320
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18746 2208 19066 3232
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 18746 1120 19066 2144
rect 19382 1325 19442 16491
rect 19566 8397 19626 21115
rect 19750 9485 19810 38795
rect 20115 38724 20181 38725
rect 20115 38660 20116 38724
rect 20180 38660 20181 38724
rect 20115 38659 20181 38660
rect 19931 24580 19997 24581
rect 19931 24516 19932 24580
rect 19996 24516 19997 24580
rect 19931 24515 19997 24516
rect 19934 21181 19994 24515
rect 19931 21180 19997 21181
rect 19931 21116 19932 21180
rect 19996 21116 19997 21180
rect 19931 21115 19997 21116
rect 20118 17237 20178 38659
rect 20299 26892 20365 26893
rect 20299 26828 20300 26892
rect 20364 26828 20365 26892
rect 20299 26827 20365 26828
rect 20115 17236 20181 17237
rect 20115 17172 20116 17236
rect 20180 17172 20181 17236
rect 20115 17171 20181 17172
rect 20302 17101 20362 26827
rect 20299 17100 20365 17101
rect 20299 17036 20300 17100
rect 20364 17036 20365 17100
rect 20299 17035 20365 17036
rect 20670 16693 20730 42059
rect 21590 41037 21650 43147
rect 21713 43008 22033 43568
rect 21713 42944 21721 43008
rect 21785 42944 21801 43008
rect 21865 42944 21881 43008
rect 21945 42944 21961 43008
rect 22025 42944 22033 43008
rect 21713 41920 22033 42944
rect 21713 41856 21721 41920
rect 21785 41856 21801 41920
rect 21865 41856 21881 41920
rect 21945 41856 21961 41920
rect 22025 41856 22033 41920
rect 21587 41036 21653 41037
rect 21587 40972 21588 41036
rect 21652 40972 21653 41036
rect 21587 40971 21653 40972
rect 21713 40832 22033 41856
rect 21713 40768 21721 40832
rect 21785 40768 21801 40832
rect 21865 40768 21881 40832
rect 21945 40768 21961 40832
rect 22025 40768 22033 40832
rect 21713 39744 22033 40768
rect 21713 39680 21721 39744
rect 21785 39680 21801 39744
rect 21865 39680 21881 39744
rect 21945 39680 21961 39744
rect 22025 39680 22033 39744
rect 21713 38656 22033 39680
rect 21713 38592 21721 38656
rect 21785 38592 21801 38656
rect 21865 38592 21881 38656
rect 21945 38592 21961 38656
rect 22025 38592 22033 38656
rect 21713 37568 22033 38592
rect 21713 37504 21721 37568
rect 21785 37504 21801 37568
rect 21865 37504 21881 37568
rect 21945 37504 21961 37568
rect 22025 37504 22033 37568
rect 21713 36480 22033 37504
rect 21713 36416 21721 36480
rect 21785 36416 21801 36480
rect 21865 36416 21881 36480
rect 21945 36416 21961 36480
rect 22025 36416 22033 36480
rect 21713 35392 22033 36416
rect 24680 43552 25000 43568
rect 24680 43488 24688 43552
rect 24752 43488 24768 43552
rect 24832 43488 24848 43552
rect 24912 43488 24928 43552
rect 24992 43488 25000 43552
rect 24680 42464 25000 43488
rect 24680 42400 24688 42464
rect 24752 42400 24768 42464
rect 24832 42400 24848 42464
rect 24912 42400 24928 42464
rect 24992 42400 25000 42464
rect 24680 41376 25000 42400
rect 24680 41312 24688 41376
rect 24752 41312 24768 41376
rect 24832 41312 24848 41376
rect 24912 41312 24928 41376
rect 24992 41312 25000 41376
rect 24680 40288 25000 41312
rect 24680 40224 24688 40288
rect 24752 40224 24768 40288
rect 24832 40224 24848 40288
rect 24912 40224 24928 40288
rect 24992 40224 25000 40288
rect 24680 39200 25000 40224
rect 24680 39136 24688 39200
rect 24752 39136 24768 39200
rect 24832 39136 24848 39200
rect 24912 39136 24928 39200
rect 24992 39136 25000 39200
rect 24680 38112 25000 39136
rect 24680 38048 24688 38112
rect 24752 38048 24768 38112
rect 24832 38048 24848 38112
rect 24912 38048 24928 38112
rect 24992 38048 25000 38112
rect 24680 37024 25000 38048
rect 24680 36960 24688 37024
rect 24752 36960 24768 37024
rect 24832 36960 24848 37024
rect 24912 36960 24928 37024
rect 24992 36960 25000 37024
rect 22875 36004 22941 36005
rect 22875 35940 22876 36004
rect 22940 35940 22941 36004
rect 22875 35939 22941 35940
rect 22323 35596 22389 35597
rect 22323 35532 22324 35596
rect 22388 35532 22389 35596
rect 22323 35531 22389 35532
rect 21713 35328 21721 35392
rect 21785 35328 21801 35392
rect 21865 35328 21881 35392
rect 21945 35328 21961 35392
rect 22025 35328 22033 35392
rect 21713 34304 22033 35328
rect 21713 34240 21721 34304
rect 21785 34240 21801 34304
rect 21865 34240 21881 34304
rect 21945 34240 21961 34304
rect 22025 34240 22033 34304
rect 21713 33216 22033 34240
rect 21713 33152 21721 33216
rect 21785 33152 21801 33216
rect 21865 33152 21881 33216
rect 21945 33152 21961 33216
rect 22025 33152 22033 33216
rect 21713 32128 22033 33152
rect 21713 32064 21721 32128
rect 21785 32064 21801 32128
rect 21865 32064 21881 32128
rect 21945 32064 21961 32128
rect 22025 32064 22033 32128
rect 21713 31040 22033 32064
rect 21713 30976 21721 31040
rect 21785 30976 21801 31040
rect 21865 30976 21881 31040
rect 21945 30976 21961 31040
rect 22025 30976 22033 31040
rect 21713 29952 22033 30976
rect 21713 29888 21721 29952
rect 21785 29888 21801 29952
rect 21865 29888 21881 29952
rect 21945 29888 21961 29952
rect 22025 29888 22033 29952
rect 20851 29068 20917 29069
rect 20851 29004 20852 29068
rect 20916 29004 20917 29068
rect 20851 29003 20917 29004
rect 20667 16692 20733 16693
rect 20667 16628 20668 16692
rect 20732 16628 20733 16692
rect 20667 16627 20733 16628
rect 19931 13700 19997 13701
rect 19931 13636 19932 13700
rect 19996 13636 19997 13700
rect 19931 13635 19997 13636
rect 19747 9484 19813 9485
rect 19747 9420 19748 9484
rect 19812 9420 19813 9484
rect 19747 9419 19813 9420
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 19379 1324 19445 1325
rect 19379 1260 19380 1324
rect 19444 1260 19445 1324
rect 19379 1259 19445 1260
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 19934 917 19994 13635
rect 20854 13565 20914 29003
rect 21713 28864 22033 29888
rect 21713 28800 21721 28864
rect 21785 28800 21801 28864
rect 21865 28800 21881 28864
rect 21945 28800 21961 28864
rect 22025 28800 22033 28864
rect 21713 27776 22033 28800
rect 21713 27712 21721 27776
rect 21785 27712 21801 27776
rect 21865 27712 21881 27776
rect 21945 27712 21961 27776
rect 22025 27712 22033 27776
rect 21219 27028 21285 27029
rect 21219 26964 21220 27028
rect 21284 26964 21285 27028
rect 21219 26963 21285 26964
rect 21222 19685 21282 26963
rect 21713 26688 22033 27712
rect 21713 26624 21721 26688
rect 21785 26624 21801 26688
rect 21865 26624 21881 26688
rect 21945 26624 21961 26688
rect 22025 26624 22033 26688
rect 21713 25600 22033 26624
rect 21713 25536 21721 25600
rect 21785 25536 21801 25600
rect 21865 25536 21881 25600
rect 21945 25536 21961 25600
rect 22025 25536 22033 25600
rect 21713 24512 22033 25536
rect 21713 24448 21721 24512
rect 21785 24448 21801 24512
rect 21865 24448 21881 24512
rect 21945 24448 21961 24512
rect 22025 24448 22033 24512
rect 21713 23424 22033 24448
rect 21713 23360 21721 23424
rect 21785 23360 21801 23424
rect 21865 23360 21881 23424
rect 21945 23360 21961 23424
rect 22025 23360 22033 23424
rect 21713 22336 22033 23360
rect 21713 22272 21721 22336
rect 21785 22272 21801 22336
rect 21865 22272 21881 22336
rect 21945 22272 21961 22336
rect 22025 22272 22033 22336
rect 21713 21248 22033 22272
rect 21713 21184 21721 21248
rect 21785 21184 21801 21248
rect 21865 21184 21881 21248
rect 21945 21184 21961 21248
rect 22025 21184 22033 21248
rect 21713 20160 22033 21184
rect 21713 20096 21721 20160
rect 21785 20096 21801 20160
rect 21865 20096 21881 20160
rect 21945 20096 21961 20160
rect 22025 20096 22033 20160
rect 21219 19684 21285 19685
rect 21219 19620 21220 19684
rect 21284 19620 21285 19684
rect 21219 19619 21285 19620
rect 21713 19072 22033 20096
rect 21713 19008 21721 19072
rect 21785 19008 21801 19072
rect 21865 19008 21881 19072
rect 21945 19008 21961 19072
rect 22025 19008 22033 19072
rect 21713 17984 22033 19008
rect 21713 17920 21721 17984
rect 21785 17920 21801 17984
rect 21865 17920 21881 17984
rect 21945 17920 21961 17984
rect 22025 17920 22033 17984
rect 21713 16896 22033 17920
rect 21713 16832 21721 16896
rect 21785 16832 21801 16896
rect 21865 16832 21881 16896
rect 21945 16832 21961 16896
rect 22025 16832 22033 16896
rect 21713 15808 22033 16832
rect 21713 15744 21721 15808
rect 21785 15744 21801 15808
rect 21865 15744 21881 15808
rect 21945 15744 21961 15808
rect 22025 15744 22033 15808
rect 21713 14720 22033 15744
rect 21713 14656 21721 14720
rect 21785 14656 21801 14720
rect 21865 14656 21881 14720
rect 21945 14656 21961 14720
rect 22025 14656 22033 14720
rect 21713 13632 22033 14656
rect 21713 13568 21721 13632
rect 21785 13568 21801 13632
rect 21865 13568 21881 13632
rect 21945 13568 21961 13632
rect 22025 13568 22033 13632
rect 20851 13564 20917 13565
rect 20851 13500 20852 13564
rect 20916 13500 20917 13564
rect 20851 13499 20917 13500
rect 21713 12544 22033 13568
rect 21713 12480 21721 12544
rect 21785 12480 21801 12544
rect 21865 12480 21881 12544
rect 21945 12480 21961 12544
rect 22025 12480 22033 12544
rect 21713 11456 22033 12480
rect 21713 11392 21721 11456
rect 21785 11392 21801 11456
rect 21865 11392 21881 11456
rect 21945 11392 21961 11456
rect 22025 11392 22033 11456
rect 21713 10368 22033 11392
rect 21713 10304 21721 10368
rect 21785 10304 21801 10368
rect 21865 10304 21881 10368
rect 21945 10304 21961 10368
rect 22025 10304 22033 10368
rect 21587 10164 21653 10165
rect 21587 10100 21588 10164
rect 21652 10100 21653 10164
rect 21587 10099 21653 10100
rect 20483 8396 20549 8397
rect 20483 8332 20484 8396
rect 20548 8332 20549 8396
rect 20483 8331 20549 8332
rect 20299 3772 20365 3773
rect 20299 3708 20300 3772
rect 20364 3708 20365 3772
rect 20299 3707 20365 3708
rect 20302 2549 20362 3707
rect 20299 2548 20365 2549
rect 20299 2484 20300 2548
rect 20364 2484 20365 2548
rect 20299 2483 20365 2484
rect 20486 1325 20546 8331
rect 21590 4045 21650 10099
rect 21713 9280 22033 10304
rect 21713 9216 21721 9280
rect 21785 9216 21801 9280
rect 21865 9216 21881 9280
rect 21945 9216 21961 9280
rect 22025 9216 22033 9280
rect 21713 8192 22033 9216
rect 21713 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22033 8192
rect 21713 7104 22033 8128
rect 21713 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22033 7104
rect 21713 6016 22033 7040
rect 22326 6357 22386 35531
rect 22691 33284 22757 33285
rect 22691 33220 22692 33284
rect 22756 33220 22757 33284
rect 22691 33219 22757 33220
rect 22507 24852 22573 24853
rect 22507 24788 22508 24852
rect 22572 24788 22573 24852
rect 22507 24787 22573 24788
rect 22323 6356 22389 6357
rect 22323 6292 22324 6356
rect 22388 6292 22389 6356
rect 22323 6291 22389 6292
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21587 4044 21653 4045
rect 21587 3980 21588 4044
rect 21652 3980 21653 4044
rect 21587 3979 21653 3980
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 22510 3229 22570 24787
rect 22694 23629 22754 33219
rect 22878 24309 22938 35939
rect 24680 35936 25000 36960
rect 24680 35872 24688 35936
rect 24752 35872 24768 35936
rect 24832 35872 24848 35936
rect 24912 35872 24928 35936
rect 24992 35872 25000 35936
rect 24680 34848 25000 35872
rect 24680 34784 24688 34848
rect 24752 34784 24768 34848
rect 24832 34784 24848 34848
rect 24912 34784 24928 34848
rect 24992 34784 25000 34848
rect 24680 33760 25000 34784
rect 24680 33696 24688 33760
rect 24752 33696 24768 33760
rect 24832 33696 24848 33760
rect 24912 33696 24928 33760
rect 24992 33696 25000 33760
rect 24680 32672 25000 33696
rect 24680 32608 24688 32672
rect 24752 32608 24768 32672
rect 24832 32608 24848 32672
rect 24912 32608 24928 32672
rect 24992 32608 25000 32672
rect 23243 31788 23309 31789
rect 23243 31724 23244 31788
rect 23308 31724 23309 31788
rect 23243 31723 23309 31724
rect 22875 24308 22941 24309
rect 22875 24244 22876 24308
rect 22940 24244 22941 24308
rect 22875 24243 22941 24244
rect 22691 23628 22757 23629
rect 22691 23564 22692 23628
rect 22756 23564 22757 23628
rect 22691 23563 22757 23564
rect 22691 23492 22757 23493
rect 22691 23428 22692 23492
rect 22756 23428 22757 23492
rect 22691 23427 22757 23428
rect 22694 15469 22754 23427
rect 22691 15468 22757 15469
rect 22691 15404 22692 15468
rect 22756 15404 22757 15468
rect 22691 15403 22757 15404
rect 22507 3228 22573 3229
rect 22507 3164 22508 3228
rect 22572 3164 22573 3228
rect 22507 3163 22573 3164
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 21713 1664 22033 2688
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 20483 1324 20549 1325
rect 20483 1260 20484 1324
rect 20548 1260 20549 1324
rect 20483 1259 20549 1260
rect 21713 1040 22033 1600
rect 23246 1189 23306 31723
rect 24680 31584 25000 32608
rect 24680 31520 24688 31584
rect 24752 31520 24768 31584
rect 24832 31520 24848 31584
rect 24912 31520 24928 31584
rect 24992 31520 25000 31584
rect 24680 30496 25000 31520
rect 24680 30432 24688 30496
rect 24752 30432 24768 30496
rect 24832 30432 24848 30496
rect 24912 30432 24928 30496
rect 24992 30432 25000 30496
rect 24680 29408 25000 30432
rect 24680 29344 24688 29408
rect 24752 29344 24768 29408
rect 24832 29344 24848 29408
rect 24912 29344 24928 29408
rect 24992 29344 25000 29408
rect 24680 28320 25000 29344
rect 24680 28256 24688 28320
rect 24752 28256 24768 28320
rect 24832 28256 24848 28320
rect 24912 28256 24928 28320
rect 24992 28256 25000 28320
rect 24680 27232 25000 28256
rect 24680 27168 24688 27232
rect 24752 27168 24768 27232
rect 24832 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 25000 27232
rect 24680 26144 25000 27168
rect 24680 26080 24688 26144
rect 24752 26080 24768 26144
rect 24832 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 25000 26144
rect 24680 25056 25000 26080
rect 24680 24992 24688 25056
rect 24752 24992 24768 25056
rect 24832 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 25000 25056
rect 24680 23968 25000 24992
rect 24680 23904 24688 23968
rect 24752 23904 24768 23968
rect 24832 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 25000 23968
rect 24680 22880 25000 23904
rect 24680 22816 24688 22880
rect 24752 22816 24768 22880
rect 24832 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 25000 22880
rect 24680 21792 25000 22816
rect 24680 21728 24688 21792
rect 24752 21728 24768 21792
rect 24832 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 25000 21792
rect 24680 20704 25000 21728
rect 24680 20640 24688 20704
rect 24752 20640 24768 20704
rect 24832 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 25000 20704
rect 24680 19616 25000 20640
rect 24680 19552 24688 19616
rect 24752 19552 24768 19616
rect 24832 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 25000 19616
rect 24680 18528 25000 19552
rect 24680 18464 24688 18528
rect 24752 18464 24768 18528
rect 24832 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 25000 18528
rect 24680 17440 25000 18464
rect 24680 17376 24688 17440
rect 24752 17376 24768 17440
rect 24832 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 25000 17440
rect 24680 16352 25000 17376
rect 24680 16288 24688 16352
rect 24752 16288 24768 16352
rect 24832 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 25000 16352
rect 24680 15264 25000 16288
rect 24680 15200 24688 15264
rect 24752 15200 24768 15264
rect 24832 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 25000 15264
rect 24680 14176 25000 15200
rect 24680 14112 24688 14176
rect 24752 14112 24768 14176
rect 24832 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 25000 14176
rect 24680 13088 25000 14112
rect 24680 13024 24688 13088
rect 24752 13024 24768 13088
rect 24832 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 25000 13088
rect 24680 12000 25000 13024
rect 24680 11936 24688 12000
rect 24752 11936 24768 12000
rect 24832 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 25000 12000
rect 24680 10912 25000 11936
rect 24680 10848 24688 10912
rect 24752 10848 24768 10912
rect 24832 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 25000 10912
rect 24680 9824 25000 10848
rect 24680 9760 24688 9824
rect 24752 9760 24768 9824
rect 24832 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 25000 9824
rect 24680 8736 25000 9760
rect 24680 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25000 8736
rect 24680 7648 25000 8672
rect 24680 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25000 7648
rect 24680 6560 25000 7584
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 23243 1188 23309 1189
rect 23243 1124 23244 1188
rect 23308 1124 23309 1188
rect 23243 1123 23309 1124
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
rect 19931 916 19997 917
rect 19931 852 19932 916
rect 19996 852 19997 916
rect 19931 851 19997 852
<< via4 >>
rect 3102 21982 3338 22218
rect 12486 21982 12722 22218
<< metal5 >>
rect 3060 22218 12764 22260
rect 3060 21982 3102 22218
rect 3338 21982 12486 22218
rect 12722 21982 12764 22218
rect 3060 21940 12764 21982
use sky130_fd_sc_hd__clkbuf_1  _000_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _001_
timestamp 1688980957
transform 1 0 23276 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp 1688980957
transform 1 0 23184 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp 1688980957
transform 1 0 23184 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _004_
timestamp 1688980957
transform 1 0 23368 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp 1688980957
transform 1 0 23276 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp 1688980957
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp 1688980957
transform 1 0 22816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp 1688980957
transform 1 0 23552 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _009_
timestamp 1688980957
transform 1 0 21620 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp 1688980957
transform 1 0 23092 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp 1688980957
transform 1 0 23644 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _013_
timestamp 1688980957
transform 1 0 23092 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _014_
timestamp 1688980957
transform 1 0 23736 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _015_
timestamp 1688980957
transform 1 0 20792 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _016_
timestamp 1688980957
transform 1 0 22356 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _017_
timestamp 1688980957
transform 1 0 22816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _018_
timestamp 1688980957
transform 1 0 22356 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp 1688980957
transform 1 0 20608 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _020_
timestamp 1688980957
transform 1 0 21620 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _021_
timestamp 1688980957
transform 1 0 23644 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp 1688980957
transform 1 0 23368 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp 1688980957
transform 1 0 23644 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp 1688980957
transform 1 0 19780 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp 1688980957
transform 1 0 20056 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp 1688980957
transform 1 0 23460 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp 1688980957
transform 1 0 21160 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp 1688980957
transform 1 0 21344 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform 1 0 22356 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform 1 0 20240 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1688980957
transform 1 0 20516 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1688980957
transform 1 0 20332 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform 1 0 23000 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform 1 0 22080 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform 1 0 20792 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp 1688980957
transform 1 0 17296 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1688980957
transform 1 0 22356 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform 1 0 21160 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform 1 0 21620 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform 1 0 21068 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform 1 0 23644 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform 1 0 20884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 22080 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1688980957
transform 1 0 20608 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp 1688980957
transform 1 0 23092 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1688980957
transform 1 0 12696 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp 1688980957
transform 1 0 15272 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform 1 0 4140 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform 1 0 8372 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 3036 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 3404 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform 1 0 3128 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 5152 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 4048 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 4600 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 4324 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 5704 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform 1 0 5428 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 7176 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 7544 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 7820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 8096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 7728 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 9936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 10580 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform 1 0 13340 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform 1 0 11316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1688980957
transform 1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1688980957
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1688980957
transform 1 0 18308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 16744 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1688980957
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1688980957
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1688980957
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1688980957
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1688980957
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform 1 0 1472 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _145_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1688980957
transform 1 0 1472 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1688980957
transform 1 0 3220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp 1688980957
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform 1 0 2576 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1688980957
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 4232 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 2944 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 4600 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 12972 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 6808 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 2944 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 3128 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 23552 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 23092 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1688980957
transform 1 0 8188 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1688980957
transform 1 0 9384 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1688980957
transform 1 0 9292 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1688980957
transform 1 0 5612 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1688980957
transform 1 0 7360 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1688980957
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1688980957
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1688980957
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1688980957
transform 1 0 6164 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1688980957
transform 1 0 7084 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0._0_
timestamp 1688980957
transform 1 0 22724 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1._0_
timestamp 1688980957
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2._0_
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3._0_
timestamp 1688980957
transform 1 0 22632 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4._0_
timestamp 1688980957
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5._0_
timestamp 1688980957
transform 1 0 23184 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6._0_
timestamp 1688980957
transform 1 0 23460 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7._0_
timestamp 1688980957
transform 1 0 23092 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8._0_
timestamp 1688980957
transform 1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9._0_
timestamp 1688980957
transform 1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10._0_
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11._0_
timestamp 1688980957
transform 1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12._0_
timestamp 1688980957
transform 1 0 21896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13._0_
timestamp 1688980957
transform 1 0 23460 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14._0_
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15._0_
timestamp 1688980957
transform 1 0 18768 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16._0_
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17._0_
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18._0_
timestamp 1688980957
transform 1 0 20976 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19._0_
timestamp 1688980957
transform 1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20._0_
timestamp 1688980957
transform 1 0 20056 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21._0_
timestamp 1688980957
transform 1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22._0_
timestamp 1688980957
transform 1 0 22816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23._0_
timestamp 1688980957
transform 1 0 21896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24._0_
timestamp 1688980957
transform 1 0 19872 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25._0_
timestamp 1688980957
transform 1 0 22080 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26._0_
timestamp 1688980957
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27._0_
timestamp 1688980957
transform 1 0 22448 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28._0_
timestamp 1688980957
transform 1 0 19320 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29._0_
timestamp 1688980957
transform 1 0 20608 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30._0_
timestamp 1688980957
transform 1 0 23184 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31._0_
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0._0_
timestamp 1688980957
transform 1 0 23552 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1._0_
timestamp 1688980957
transform 1 0 23736 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2._0_
timestamp 1688980957
transform 1 0 23460 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3._0_
timestamp 1688980957
transform 1 0 23460 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4._0_
timestamp 1688980957
transform 1 0 23644 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5._0_
timestamp 1688980957
transform 1 0 23552 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6._0_
timestamp 1688980957
transform 1 0 23736 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7._0_
timestamp 1688980957
transform 1 0 23460 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8._0_
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9._0_
timestamp 1688980957
transform 1 0 21160 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10._0_
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11._0_
timestamp 1688980957
transform 1 0 23368 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12._0_
timestamp 1688980957
transform 1 0 22816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13._0_
timestamp 1688980957
transform 1 0 23368 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14._0_
timestamp 1688980957
transform 1 0 23184 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15._0_
timestamp 1688980957
transform 1 0 19872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16._0_
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17._0_
timestamp 1688980957
transform 1 0 23092 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18._0_
timestamp 1688980957
transform 1 0 21620 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19._0_
timestamp 1688980957
transform 1 0 19596 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20._0_
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21._0_
timestamp 1688980957
transform 1 0 23644 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22._0_
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23._0_
timestamp 1688980957
transform 1 0 23000 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24._0_
timestamp 1688980957
transform 1 0 20424 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25._0_
timestamp 1688980957
transform 1 0 22816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26._0_
timestamp 1688980957
transform 1 0 20884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27._0_
timestamp 1688980957
transform 1 0 20240 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28._0_
timestamp 1688980957
transform 1 0 19964 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29._0_
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30._0_
timestamp 1688980957
transform 1 0 21160 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31._0_
timestamp 1688980957
transform 1 0 20332 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_35
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_88
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_98
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_21
timestamp 1688980957
transform 1 0 3036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_127
timestamp 1688980957
transform 1 0 12788 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_131
timestamp 1688980957
transform 1 0 13156 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_139
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_233
timestamp 1688980957
transform 1 0 22540 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_11
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_36
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_43
timestamp 1688980957
transform 1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_66
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_88
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_110
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_120
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_124
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_129
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_151
timestamp 1688980957
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_162 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_241
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_13
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_21
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_88
timestamp 1688980957
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_92
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_116
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_135
timestamp 1688980957
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_155
timestamp 1688980957
transform 1 0 15364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_159
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_173
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_199
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_210
timestamp 1688980957
transform 1 0 20424 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_235
timestamp 1688980957
transform 1 0 22724 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1688980957
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_58
timestamp 1688980957
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_64
timestamp 1688980957
transform 1 0 6992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_106
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_110
timestamp 1688980957
transform 1 0 11224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_156
timestamp 1688980957
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_168
timestamp 1688980957
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_172
timestamp 1688980957
transform 1 0 16928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_176
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_180
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_38
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_128
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_183
timestamp 1688980957
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1688980957
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_250
timestamp 1688980957
transform 1 0 24104 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_35
timestamp 1688980957
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_52
timestamp 1688980957
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_64
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_170
timestamp 1688980957
transform 1 0 16744 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_176
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_224
timestamp 1688980957
transform 1 0 21712 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_231
timestamp 1688980957
transform 1 0 22356 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_72
timestamp 1688980957
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_103
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_52
timestamp 1688980957
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_125
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 1688980957
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_212
timestamp 1688980957
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_238
timestamp 1688980957
transform 1 0 23000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_29
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_177
timestamp 1688980957
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_184
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_196
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_202
timestamp 1688980957
transform 1 0 19688 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_35
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_52
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_64
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_76
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_106
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_118
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_238
timestamp 1688980957
transform 1 0 23000 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp 1688980957
transform 1 0 23736 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_148
timestamp 1688980957
transform 1 0 14720 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_160
timestamp 1688980957
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_201
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_228
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_245
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_35
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_207
timestamp 1688980957
transform 1 0 20148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_83
timestamp 1688980957
transform 1 0 8740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_131
timestamp 1688980957
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_135
timestamp 1688980957
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_238
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_35
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_47
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_59
timestamp 1688980957
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_67
timestamp 1688980957
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_186
timestamp 1688980957
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1688980957
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_217
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_24
timestamp 1688980957
transform 1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_143
timestamp 1688980957
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_218
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_234
timestamp 1688980957
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_253
timestamp 1688980957
transform 1 0 24380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_71
timestamp 1688980957
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_129
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_156
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_180
timestamp 1688980957
transform 1 0 17664 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_186
timestamp 1688980957
transform 1 0 18216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_190
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_205
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_229
timestamp 1688980957
transform 1 0 22172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_72
timestamp 1688980957
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_84
timestamp 1688980957
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_103
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1688980957
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_152
timestamp 1688980957
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1688980957
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_231
timestamp 1688980957
transform 1 0 22356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_250
timestamp 1688980957
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_254
timestamp 1688980957
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_58
timestamp 1688980957
transform 1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_79
timestamp 1688980957
transform 1 0 8372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_106
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_110
timestamp 1688980957
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_114
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_126
timestamp 1688980957
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_200
timestamp 1688980957
transform 1 0 19504 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_217
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_229
timestamp 1688980957
transform 1 0 22172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_143
timestamp 1688980957
transform 1 0 14260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_199
timestamp 1688980957
transform 1 0 19412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_211
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_219
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_238
timestamp 1688980957
transform 1 0 23000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_159
timestamp 1688980957
transform 1 0 15732 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_203
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_72
timestamp 1688980957
transform 1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_130
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_154
timestamp 1688980957
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_185
timestamp 1688980957
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_246
timestamp 1688980957
transform 1 0 23736 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_253
timestamp 1688980957
transform 1 0 24380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_44
timestamp 1688980957
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_56
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_68
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_92
timestamp 1688980957
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_123
timestamp 1688980957
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_183
timestamp 1688980957
transform 1 0 17940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_61
timestamp 1688980957
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_121
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_144
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_162
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_202
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_233
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_248
timestamp 1688980957
transform 1 0 23920 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_35
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_39
timestamp 1688980957
transform 1 0 4692 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_218
timestamp 1688980957
transform 1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_224
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_235
timestamp 1688980957
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_50
timestamp 1688980957
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_86
timestamp 1688980957
transform 1 0 9016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_103
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_131
timestamp 1688980957
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_154
timestamp 1688980957
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_190
timestamp 1688980957
transform 1 0 18584 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_198
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_240
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_44
timestamp 1688980957
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_185
timestamp 1688980957
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_212
timestamp 1688980957
transform 1 0 20608 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_224
timestamp 1688980957
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_99
timestamp 1688980957
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_134
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_142
timestamp 1688980957
transform 1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_204
timestamp 1688980957
transform 1 0 19872 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1688980957
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_233
timestamp 1688980957
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_253
timestamp 1688980957
transform 1 0 24380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_17
timestamp 1688980957
transform 1 0 2668 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_35
timestamp 1688980957
transform 1 0 4324 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_47
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_59
timestamp 1688980957
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_183
timestamp 1688980957
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_222
timestamp 1688980957
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_230
timestamp 1688980957
transform 1 0 22264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_30
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_38
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_75
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_79
timestamp 1688980957
transform 1 0 8372 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_91
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_124
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_140
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_184
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_196
timestamp 1688980957
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_203
timestamp 1688980957
transform 1 0 19780 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_209
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_214
timestamp 1688980957
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_219
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_240
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_118
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_144
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_156
timestamp 1688980957
transform 1 0 15456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_168
timestamp 1688980957
transform 1 0 16560 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_192
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_9
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_29
timestamp 1688980957
transform 1 0 3772 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_131
timestamp 1688980957
transform 1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_139
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_157
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_173
timestamp 1688980957
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_207
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_219
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_24
timestamp 1688980957
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_44
timestamp 1688980957
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_56
timestamp 1688980957
transform 1 0 6256 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_64
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_125
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_159
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_204
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_208
timestamp 1688980957
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_220
timestamp 1688980957
transform 1 0 21344 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_232
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_241
timestamp 1688980957
transform 1 0 23276 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_99
timestamp 1688980957
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_128
timestamp 1688980957
transform 1 0 12880 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_184
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_235
timestamp 1688980957
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_239
timestamp 1688980957
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_32
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_38
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_78
timestamp 1688980957
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_113
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_179
timestamp 1688980957
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_191
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_250
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_18
timestamp 1688980957
transform 1 0 2760 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_143
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 1688980957
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_196
timestamp 1688980957
transform 1 0 19136 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_208
timestamp 1688980957
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1688980957
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_56
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_68
timestamp 1688980957
transform 1 0 7360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_115
timestamp 1688980957
transform 1 0 11684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_147
timestamp 1688980957
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_169
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_187
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_200
timestamp 1688980957
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_208
timestamp 1688980957
transform 1 0 20240 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_212
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_216
timestamp 1688980957
transform 1 0 20976 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_228
timestamp 1688980957
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_232
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_24
timestamp 1688980957
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_36
timestamp 1688980957
transform 1 0 4416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1688980957
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_75
timestamp 1688980957
transform 1 0 8004 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_96
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 1688980957
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_131
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_147
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_196
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_200
timestamp 1688980957
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_228
timestamp 1688980957
transform 1 0 22080 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_240
timestamp 1688980957
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_26
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_32
timestamp 1688980957
transform 1 0 4048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_36
timestamp 1688980957
transform 1 0 4416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_55
timestamp 1688980957
transform 1 0 6164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_75
timestamp 1688980957
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_130
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_162
timestamp 1688980957
transform 1 0 16008 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_180
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_213
timestamp 1688980957
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_217
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_225
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_234
timestamp 1688980957
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_238
timestamp 1688980957
transform 1 0 23000 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_18
timestamp 1688980957
transform 1 0 2760 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_25
timestamp 1688980957
transform 1 0 3404 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_48
timestamp 1688980957
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_72
timestamp 1688980957
transform 1 0 7728 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_84
timestamp 1688980957
transform 1 0 8832 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_96
timestamp 1688980957
transform 1 0 9936 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_145
timestamp 1688980957
transform 1 0 14444 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_150
timestamp 1688980957
transform 1 0 14904 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_190
timestamp 1688980957
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_214
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_220
timestamp 1688980957
transform 1 0 21344 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_9
timestamp 1688980957
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_44
timestamp 1688980957
transform 1 0 5152 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_56
timestamp 1688980957
transform 1 0 6256 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_68
timestamp 1688980957
transform 1 0 7360 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_100
timestamp 1688980957
transform 1 0 10304 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_119
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_131
timestamp 1688980957
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_156
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_168
timestamp 1688980957
transform 1 0 16560 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_180
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_191
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_200
timestamp 1688980957
transform 1 0 19504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_205
timestamp 1688980957
transform 1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_211
timestamp 1688980957
transform 1 0 20516 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_247
timestamp 1688980957
transform 1 0 23828 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_13
timestamp 1688980957
transform 1 0 2300 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_33
timestamp 1688980957
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 1688980957
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_100
timestamp 1688980957
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_120
timestamp 1688980957
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_124
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_146
timestamp 1688980957
transform 1 0 14536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_213
timestamp 1688980957
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_233
timestamp 1688980957
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_239
timestamp 1688980957
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_21
timestamp 1688980957
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_68
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_75
timestamp 1688980957
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_100
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_118
timestamp 1688980957
transform 1 0 11960 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_124
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_149
timestamp 1688980957
transform 1 0 14812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_187
timestamp 1688980957
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_206
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_212
timestamp 1688980957
transform 1 0 20608 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_218
timestamp 1688980957
transform 1 0 21160 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_230
timestamp 1688980957
transform 1 0 22264 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_77
timestamp 1688980957
transform 1 0 8188 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_95
timestamp 1688980957
transform 1 0 9844 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_119
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_135
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_159
timestamp 1688980957
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_199
timestamp 1688980957
transform 1 0 19412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_203
timestamp 1688980957
transform 1 0 19780 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_228
timestamp 1688980957
transform 1 0 22080 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_247
timestamp 1688980957
transform 1 0 23828 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_12
timestamp 1688980957
transform 1 0 2208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_62
timestamp 1688980957
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_66
timestamp 1688980957
transform 1 0 7176 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_82
timestamp 1688980957
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_106
timestamp 1688980957
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_128
timestamp 1688980957
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_200
timestamp 1688980957
transform 1 0 19504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_204
timestamp 1688980957
transform 1 0 19872 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_208
timestamp 1688980957
transform 1 0 20240 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_224
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_241
timestamp 1688980957
transform 1 0 23276 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_107
timestamp 1688980957
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_128
timestamp 1688980957
transform 1 0 12880 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_151
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_163
timestamp 1688980957
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_212
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_234
timestamp 1688980957
transform 1 0 22632 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_241
timestamp 1688980957
transform 1 0 23276 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_20
timestamp 1688980957
transform 1 0 2944 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_35
timestamp 1688980957
transform 1 0 4324 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_47
timestamp 1688980957
transform 1 0 5428 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_74
timestamp 1688980957
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_82
timestamp 1688980957
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_129
timestamp 1688980957
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_172
timestamp 1688980957
transform 1 0 16928 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_200
timestamp 1688980957
transform 1 0 19504 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_212
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_224
timestamp 1688980957
transform 1 0 21712 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_232
timestamp 1688980957
transform 1 0 22448 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_238
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_242
timestamp 1688980957
transform 1 0 23368 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_7
timestamp 1688980957
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_29
timestamp 1688980957
transform 1 0 3772 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_52
timestamp 1688980957
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_87
timestamp 1688980957
transform 1 0 9108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_99
timestamp 1688980957
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1688980957
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_190
timestamp 1688980957
transform 1 0 18584 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_202
timestamp 1688980957
transform 1 0 19688 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_214
timestamp 1688980957
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_240
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_247
timestamp 1688980957
transform 1 0 23828 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_24
timestamp 1688980957
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_73
timestamp 1688980957
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_106
timestamp 1688980957
transform 1 0 10856 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_112
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_128
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_149
timestamp 1688980957
transform 1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_154
timestamp 1688980957
transform 1 0 15272 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_162
timestamp 1688980957
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_208
timestamp 1688980957
transform 1 0 20240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_214
timestamp 1688980957
transform 1 0 20792 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_247
timestamp 1688980957
transform 1 0 23828 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_11
timestamp 1688980957
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_34
timestamp 1688980957
transform 1 0 4232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1688980957
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_72
timestamp 1688980957
transform 1 0 7728 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_84
timestamp 1688980957
transform 1 0 8832 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_96
timestamp 1688980957
transform 1 0 9936 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_148
timestamp 1688980957
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_152
timestamp 1688980957
transform 1 0 15088 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_198
timestamp 1688980957
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_231
timestamp 1688980957
transform 1 0 22356 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_45
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_57
timestamp 1688980957
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_69
timestamp 1688980957
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_100
timestamp 1688980957
transform 1 0 10304 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_114
timestamp 1688980957
transform 1 0 11592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_130
timestamp 1688980957
transform 1 0 13064 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_156
timestamp 1688980957
transform 1 0 15456 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_183
timestamp 1688980957
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_187
timestamp 1688980957
transform 1 0 18308 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_191
timestamp 1688980957
transform 1 0 18676 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_200
timestamp 1688980957
transform 1 0 19504 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_220
timestamp 1688980957
transform 1 0 21344 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_232
timestamp 1688980957
transform 1 0 22448 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_237
timestamp 1688980957
transform 1 0 22908 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_246
timestamp 1688980957
transform 1 0 23736 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_11
timestamp 1688980957
transform 1 0 2116 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_30
timestamp 1688980957
transform 1 0 3864 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_38
timestamp 1688980957
transform 1 0 4600 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_83
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_87
timestamp 1688980957
transform 1 0 9108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_107
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_117
timestamp 1688980957
transform 1 0 11868 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_123
timestamp 1688980957
transform 1 0 12420 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_139
timestamp 1688980957
transform 1 0 13892 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_159
timestamp 1688980957
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_184
timestamp 1688980957
transform 1 0 18032 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_192
timestamp 1688980957
transform 1 0 18768 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_211
timestamp 1688980957
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_248
timestamp 1688980957
transform 1 0 23920 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_24
timestamp 1688980957
transform 1 0 3312 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_39
timestamp 1688980957
transform 1 0 4692 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_58
timestamp 1688980957
transform 1 0 6440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_62
timestamp 1688980957
transform 1 0 6808 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_101
timestamp 1688980957
transform 1 0 10396 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_178
timestamp 1688980957
transform 1 0 17480 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_190
timestamp 1688980957
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_215
timestamp 1688980957
transform 1 0 20884 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_219
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_226
timestamp 1688980957
transform 1 0 21896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_234
timestamp 1688980957
transform 1 0 22632 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_240
timestamp 1688980957
transform 1 0 23184 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_247
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_28
timestamp 1688980957
transform 1 0 3680 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_32
timestamp 1688980957
transform 1 0 4048 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_48
timestamp 1688980957
transform 1 0 5520 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_61
timestamp 1688980957
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_89
timestamp 1688980957
transform 1 0 9292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_95
timestamp 1688980957
transform 1 0 9844 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_154
timestamp 1688980957
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_166
timestamp 1688980957
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_198
timestamp 1688980957
transform 1 0 19320 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_206
timestamp 1688980957
transform 1 0 20056 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_7
timestamp 1688980957
transform 1 0 1748 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_32
timestamp 1688980957
transform 1 0 4048 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_49
timestamp 1688980957
transform 1 0 5612 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_72
timestamp 1688980957
transform 1 0 7728 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_100
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_123
timestamp 1688980957
transform 1 0 12420 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 1688980957
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_154
timestamp 1688980957
transform 1 0 15272 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_158
timestamp 1688980957
transform 1 0 15640 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_207
timestamp 1688980957
transform 1 0 20148 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_211
timestamp 1688980957
transform 1 0 20516 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_215
timestamp 1688980957
transform 1 0 20884 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_227
timestamp 1688980957
transform 1 0 21988 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_231
timestamp 1688980957
transform 1 0 22356 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_235
timestamp 1688980957
transform 1 0 22724 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_242
timestamp 1688980957
transform 1 0 23368 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_49
timestamp 1688980957
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_75
timestamp 1688980957
transform 1 0 8004 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_79
timestamp 1688980957
transform 1 0 8372 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_98
timestamp 1688980957
transform 1 0 10120 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_117
timestamp 1688980957
transform 1 0 11868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_142
timestamp 1688980957
transform 1 0 14168 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_150
timestamp 1688980957
transform 1 0 14904 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_187
timestamp 1688980957
transform 1 0 18308 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_192
timestamp 1688980957
transform 1 0 18768 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1688980957
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_229
timestamp 1688980957
transform 1 0 22172 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_233
timestamp 1688980957
transform 1 0 22540 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_240
timestamp 1688980957
transform 1 0 23184 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_247
timestamp 1688980957
transform 1 0 23828 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_24
timestamp 1688980957
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_42
timestamp 1688980957
transform 1 0 4968 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_50
timestamp 1688980957
transform 1 0 5704 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_66
timestamp 1688980957
transform 1 0 7176 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_78
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_105
timestamp 1688980957
transform 1 0 10764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_123
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_129
timestamp 1688980957
transform 1 0 12972 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_156
timestamp 1688980957
transform 1 0 15456 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_178
timestamp 1688980957
transform 1 0 17480 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_190
timestamp 1688980957
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_203
timestamp 1688980957
transform 1 0 19780 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_226
timestamp 1688980957
transform 1 0 21896 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_238
timestamp 1688980957
transform 1 0 23000 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_241
timestamp 1688980957
transform 1 0 23276 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_90
timestamp 1688980957
transform 1 0 9384 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_96
timestamp 1688980957
transform 1 0 9936 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_157
timestamp 1688980957
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_165
timestamp 1688980957
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_212
timestamp 1688980957
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_228
timestamp 1688980957
transform 1 0 22080 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_9
timestamp 1688980957
transform 1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_58
timestamp 1688980957
transform 1 0 6440 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_81
timestamp 1688980957
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_93
timestamp 1688980957
transform 1 0 9660 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_132
timestamp 1688980957
transform 1 0 13248 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_162
timestamp 1688980957
transform 1 0 16008 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_174
timestamp 1688980957
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_178
timestamp 1688980957
transform 1 0 17480 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_194
timestamp 1688980957
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_225
timestamp 1688980957
transform 1 0 21804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_232
timestamp 1688980957
transform 1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_239
timestamp 1688980957
transform 1 0 23092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_37
timestamp 1688980957
transform 1 0 4508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_90
timestamp 1688980957
transform 1 0 9384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_106
timestamp 1688980957
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_201
timestamp 1688980957
transform 1 0 19596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_213
timestamp 1688980957
transform 1 0 20700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_248
timestamp 1688980957
transform 1 0 23920 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_24
timestamp 1688980957
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_35
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_52
timestamp 1688980957
transform 1 0 5888 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_60
timestamp 1688980957
transform 1 0 6624 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_100
timestamp 1688980957
transform 1 0 10304 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_112
timestamp 1688980957
transform 1 0 11408 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_156
timestamp 1688980957
transform 1 0 15456 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_160
timestamp 1688980957
transform 1 0 15824 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_179
timestamp 1688980957
transform 1 0 17572 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_183
timestamp 1688980957
transform 1 0 17940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_188
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_223
timestamp 1688980957
transform 1 0 21620 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_237
timestamp 1688980957
transform 1 0 22908 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_24
timestamp 1688980957
transform 1 0 3312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_47
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_72
timestamp 1688980957
transform 1 0 7728 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_80
timestamp 1688980957
transform 1 0 8464 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_87
timestamp 1688980957
transform 1 0 9108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_95
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_141
timestamp 1688980957
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_157
timestamp 1688980957
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_165
timestamp 1688980957
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_179
timestamp 1688980957
transform 1 0 17572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_191
timestamp 1688980957
transform 1 0 18676 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_243
timestamp 1688980957
transform 1 0 23460 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_248
timestamp 1688980957
transform 1 0 23920 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_9
timestamp 1688980957
transform 1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_62
timestamp 1688980957
transform 1 0 6808 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_74
timestamp 1688980957
transform 1 0 7912 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_82
timestamp 1688980957
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_93
timestamp 1688980957
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_131
timestamp 1688980957
transform 1 0 13156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_156
timestamp 1688980957
transform 1 0 15456 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_173
timestamp 1688980957
transform 1 0 17020 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_188
timestamp 1688980957
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_203
timestamp 1688980957
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_207
timestamp 1688980957
transform 1 0 20148 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_213
timestamp 1688980957
transform 1 0 20700 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_217
timestamp 1688980957
transform 1 0 21068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_229
timestamp 1688980957
transform 1 0 22172 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_237
timestamp 1688980957
transform 1 0 22908 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_246
timestamp 1688980957
transform 1 0 23736 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_31
timestamp 1688980957
transform 1 0 3956 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_108
timestamp 1688980957
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_146
timestamp 1688980957
transform 1 0 14536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_158
timestamp 1688980957
transform 1 0 15640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_166
timestamp 1688980957
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_177
timestamp 1688980957
transform 1 0 17388 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_201
timestamp 1688980957
transform 1 0 19596 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_213
timestamp 1688980957
transform 1 0 20700 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_220
timestamp 1688980957
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_228
timestamp 1688980957
transform 1 0 22080 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_242
timestamp 1688980957
transform 1 0 23368 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_25
timestamp 1688980957
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_67
timestamp 1688980957
transform 1 0 7268 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_79
timestamp 1688980957
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_173
timestamp 1688980957
transform 1 0 17020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_215
timestamp 1688980957
transform 1 0 20884 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_219
timestamp 1688980957
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_226
timestamp 1688980957
transform 1 0 21896 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_230
timestamp 1688980957
transform 1 0 22264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_234
timestamp 1688980957
transform 1 0 22632 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_84
timestamp 1688980957
transform 1 0 8832 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_96
timestamp 1688980957
transform 1 0 9936 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_108
timestamp 1688980957
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_128
timestamp 1688980957
transform 1 0 12880 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_140
timestamp 1688980957
transform 1 0 13984 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_152
timestamp 1688980957
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_164
timestamp 1688980957
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_177
timestamp 1688980957
transform 1 0 17388 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_182
timestamp 1688980957
transform 1 0 17848 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_197
timestamp 1688980957
transform 1 0 19228 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_204
timestamp 1688980957
transform 1 0 19872 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_218
timestamp 1688980957
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_233
timestamp 1688980957
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_242
timestamp 1688980957
transform 1 0 23368 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_246
timestamp 1688980957
transform 1 0 23736 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_14
timestamp 1688980957
transform 1 0 2392 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_35
timestamp 1688980957
transform 1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_54
timestamp 1688980957
transform 1 0 6072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_58
timestamp 1688980957
transform 1 0 6440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_81
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_112
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_124
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_136
timestamp 1688980957
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_214
timestamp 1688980957
transform 1 0 20792 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_222
timestamp 1688980957
transform 1 0 21528 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_229
timestamp 1688980957
transform 1 0 22172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_54
timestamp 1688980957
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_72
timestamp 1688980957
transform 1 0 7728 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_80
timestamp 1688980957
transform 1 0 8464 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_101
timestamp 1688980957
transform 1 0 10396 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_109
timestamp 1688980957
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_134
timestamp 1688980957
transform 1 0 13432 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_146
timestamp 1688980957
transform 1 0 14536 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_158
timestamp 1688980957
transform 1 0 15640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_166
timestamp 1688980957
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_250
timestamp 1688980957
transform 1 0 24104 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_25
timestamp 1688980957
transform 1 0 3404 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_44
timestamp 1688980957
transform 1 0 5152 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_67
timestamp 1688980957
transform 1 0 7268 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_79
timestamp 1688980957
transform 1 0 8372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_102
timestamp 1688980957
transform 1 0 10488 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_110
timestamp 1688980957
transform 1 0 11224 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_203
timestamp 1688980957
transform 1 0 19780 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_207
timestamp 1688980957
transform 1 0 20148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_219
timestamp 1688980957
transform 1 0 21252 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_227
timestamp 1688980957
transform 1 0 21988 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_231
timestamp 1688980957
transform 1 0 22356 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_244
timestamp 1688980957
transform 1 0 23552 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_44
timestamp 1688980957
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_75
timestamp 1688980957
transform 1 0 8004 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_91
timestamp 1688980957
transform 1 0 9476 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_103
timestamp 1688980957
transform 1 0 10580 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_128
timestamp 1688980957
transform 1 0 12880 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_140
timestamp 1688980957
transform 1 0 13984 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_152
timestamp 1688980957
transform 1 0 15088 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_164
timestamp 1688980957
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_209
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_216
timestamp 1688980957
transform 1 0 20976 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_220
timestamp 1688980957
transform 1 0 21344 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_241
timestamp 1688980957
transform 1 0 23276 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_248
timestamp 1688980957
transform 1 0 23920 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_106
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_118
timestamp 1688980957
transform 1 0 11960 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_137
timestamp 1688980957
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_216
timestamp 1688980957
transform 1 0 20976 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_220
timestamp 1688980957
transform 1 0 21344 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_234
timestamp 1688980957
transform 1 0 22632 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_239
timestamp 1688980957
transform 1 0 23092 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_243
timestamp 1688980957
transform 1 0 23460 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_36
timestamp 1688980957
transform 1 0 4416 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_40
timestamp 1688980957
transform 1 0 4784 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_65
timestamp 1688980957
transform 1 0 7084 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_103
timestamp 1688980957
transform 1 0 10580 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_109
timestamp 1688980957
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_200
timestamp 1688980957
transform 1 0 19504 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_243
timestamp 1688980957
transform 1 0 23460 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_248
timestamp 1688980957
transform 1 0 23920 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_44
timestamp 1688980957
transform 1 0 5152 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_78
timestamp 1688980957
transform 1 0 8280 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_93
timestamp 1688980957
transform 1 0 9660 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_134
timestamp 1688980957
transform 1 0 13432 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_204
timestamp 1688980957
transform 1 0 19872 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_241
timestamp 1688980957
transform 1 0 23276 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_14
timestamp 1688980957
transform 1 0 2392 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_19
timestamp 1688980957
transform 1 0 2852 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_24
timestamp 1688980957
transform 1 0 3312 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_61
timestamp 1688980957
transform 1 0 6716 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_64
timestamp 1688980957
transform 1 0 6992 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_70
timestamp 1688980957
transform 1 0 7544 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_75
timestamp 1688980957
transform 1 0 8004 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_96
timestamp 1688980957
transform 1 0 9936 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_198
timestamp 1688980957
transform 1 0 19320 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_234
timestamp 1688980957
transform 1 0 22632 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_253
timestamp 1688980957
transform 1 0 24380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_18
timestamp 1688980957
transform 1 0 2760 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_57
timestamp 1688980957
transform 1 0 6348 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_62
timestamp 1688980957
transform 1 0 6808 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_69
timestamp 1688980957
transform 1 0 7452 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_82
timestamp 1688980957
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_88
timestamp 1688980957
transform 1 0 9200 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_92
timestamp 1688980957
transform 1 0 9568 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_108
timestamp 1688980957
transform 1 0 11040 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_120
timestamp 1688980957
transform 1 0 12144 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_132
timestamp 1688980957
transform 1 0 13248 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_190
timestamp 1688980957
transform 1 0 18584 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_204
timestamp 1688980957
transform 1 0 19872 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_214
timestamp 1688980957
transform 1 0 20792 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_227
timestamp 1688980957
transform 1 0 21988 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_22
timestamp 1688980957
transform 1 0 3128 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_35
timestamp 1688980957
transform 1 0 4324 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_47
timestamp 1688980957
transform 1 0 5428 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_63
timestamp 1688980957
transform 1 0 6900 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_70
timestamp 1688980957
transform 1 0 7544 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_87
timestamp 1688980957
transform 1 0 9108 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_91
timestamp 1688980957
transform 1 0 9476 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_99
timestamp 1688980957
transform 1 0 10212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_201
timestamp 1688980957
transform 1 0 19596 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_228
timestamp 1688980957
transform 1 0 22080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_247
timestamp 1688980957
transform 1 0 23828 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_254
timestamp 1688980957
transform 1 0 24472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_9
timestamp 1688980957
transform 1 0 1932 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_58
timestamp 1688980957
transform 1 0 6440 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_76
timestamp 1688980957
transform 1 0 8096 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_88
timestamp 1688980957
transform 1 0 9200 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_96
timestamp 1688980957
transform 1 0 9936 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_106
timestamp 1688980957
transform 1 0 10856 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_120
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_132
timestamp 1688980957
transform 1 0 13248 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_150
timestamp 1688980957
transform 1 0 14904 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_160
timestamp 1688980957
transform 1 0 15824 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_164
timestamp 1688980957
transform 1 0 16192 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_220
timestamp 1688980957
transform 1 0 21344 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1688980957
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_12
timestamp 1688980957
transform 1 0 2208 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_26
timestamp 1688980957
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_32
timestamp 1688980957
transform 1 0 4048 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_42
timestamp 1688980957
transform 1 0 4968 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_50
timestamp 1688980957
transform 1 0 5704 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_85
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_117
timestamp 1688980957
transform 1 0 11868 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_130
timestamp 1688980957
transform 1 0 13064 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_145
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_155
timestamp 1688980957
transform 1 0 15364 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_173
timestamp 1688980957
transform 1 0 17020 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_194
timestamp 1688980957
transform 1 0 18952 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_203
timestamp 1688980957
transform 1 0 19780 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_247
timestamp 1688980957
transform 1 0 23828 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_253
timestamp 1688980957
transform 1 0 24380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform 1 0 3404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 2944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 2300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 2760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 3220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 3128 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 2024 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 3312 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 2576 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 3404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1688980957
transform 1 0 2760 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 3036 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2760 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3036 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 4048 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 3312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input50
timestamp 1688980957
transform 1 0 2852 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input51
timestamp 1688980957
transform 1 0 3404 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input52
timestamp 1688980957
transform 1 0 4876 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input53
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input54
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input55
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1688980957
transform 1 0 3312 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1688980957
transform 1 0 4968 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1688980957
transform 1 0 5520 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1688980957
transform 1 0 4048 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input66 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input67
timestamp 1688980957
transform 1 0 2392 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input68
timestamp 1688980957
transform 1 0 3036 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input69
timestamp 1688980957
transform 1 0 4600 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input70
timestamp 1688980957
transform 1 0 2392 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input71
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input72
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input73
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input74
timestamp 1688980957
transform 1 0 3312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input75
timestamp 1688980957
transform 1 0 3864 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input76
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1688980957
transform 1 0 2760 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input78
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1688980957
transform 1 0 2760 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input80
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1688980957
transform 1 0 22172 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1688980957
transform 1 0 23644 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1688980957
transform 1 0 21252 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1688980957
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1688980957
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1688980957
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1688980957
transform 1 0 18584 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1688980957
transform 1 0 21068 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input93
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input94
timestamp 1688980957
transform 1 0 22724 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input95
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input96
timestamp 1688980957
transform 1 0 19320 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input97
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input98
timestamp 1688980957
transform 1 0 21988 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input99
timestamp 1688980957
transform 1 0 23000 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input100
timestamp 1688980957
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1688980957
transform 1 0 4048 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1688980957
transform 1 0 3496 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1688980957
transform 1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1688980957
transform 1 0 5244 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1688980957
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1688980957
transform 1 0 2944 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1688980957
transform 1 0 4508 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1688980957
transform 1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1688980957
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input128
timestamp 1688980957
transform 1 0 4416 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input129
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1688980957
transform 1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1688980957
transform 1 0 8004 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1688980957
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1688980957
transform 1 0 22724 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1688980957
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1688980957
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1688980957
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1688980957
transform 1 0 10304 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input155
timestamp 1688980957
transform 1 0 10672 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1688980957
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input157
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1688980957
transform 1 0 11592 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1688980957
transform 1 0 11868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1688980957
transform 1 0 12328 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1688980957
transform 1 0 12696 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1688980957
transform 1 0 12972 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input165
timestamp 1688980957
transform 1 0 13616 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1688980957
transform 1 0 14628 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1688980957
transform 1 0 14352 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1688980957
transform 1 0 14628 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1688980957
transform 1 0 14996 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1688980957
transform 1 0 15548 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input172
timestamp 1688980957
transform 1 0 15456 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input173
timestamp 1688980957
transform 1 0 15824 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1688980957
transform 1 0 20792 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1688980957
transform 1 0 18768 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1688980957
transform 1 0 19596 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1688980957
transform 1 0 20516 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1688980957
transform 1 0 19504 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1688980957
transform 1 0 17940 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1688980957
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input181
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input182
timestamp 1688980957
transform 1 0 16560 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1688980957
transform 1 0 17572 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1688980957
transform 1 0 17848 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1688980957
transform 1 0 18124 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1688980957
transform 1 0 18400 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1688980957
transform 1 0 19228 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1688980957
transform 1 0 21068 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._0_
timestamp 1688980957
transform 1 0 24104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._1_
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._2_
timestamp 1688980957
transform 1 0 22448 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._3_
timestamp 1688980957
transform 1 0 23092 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 20700 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19596 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 24288 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 23000 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 22080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21160 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22172 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17112 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22356 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 22724 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22448 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19596 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20240 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19136 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20056 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 20608 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20884 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22080 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22724 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23184 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20240 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19412 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17112 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17848 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 21620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21988 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20976 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22080 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20884 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18124 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19320 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17572 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20240 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18400 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20608 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17204 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 22080 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23000 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23460 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23368 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22356 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18124 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19044 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21160 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19044 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17664 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23000 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23276 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22080 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22632 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20516 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 21344 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20976 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20792 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18492 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19596 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18032 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19872 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17848 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22356 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19872 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23184 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22632 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 21344 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20148 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19688 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 21252 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19872 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23092 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21252 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 23092 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 21528 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23092 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19596 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18952 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22816 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 22816 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 17664 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23276 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 23368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23920 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit1
timestamp 1688980957
transform 1 0 11224 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit2
timestamp 1688980957
transform 1 0 1932 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit3
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit4
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit5
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit6
timestamp 1688980957
transform 1 0 12512 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit7
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit8
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit10
timestamp 1688980957
transform 1 0 2300 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit11
timestamp 1688980957
transform 1 0 4232 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit12
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit13
timestamp 1688980957
transform 1 0 4876 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit14
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit15
timestamp 1688980957
transform 1 0 10580 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit16
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit17
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit18
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit19
timestamp 1688980957
transform 1 0 5704 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit20
timestamp 1688980957
transform 1 0 8004 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit21
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit22
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit23
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit24
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit25
timestamp 1688980957
transform 1 0 11224 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit26
timestamp 1688980957
transform 1 0 1656 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit27
timestamp 1688980957
transform 1 0 1932 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit28
timestamp 1688980957
transform 1 0 9660 0 1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit30
timestamp 1688980957
transform 1 0 12604 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit31
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit0
timestamp 1688980957
transform 1 0 12052 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit1
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit2
timestamp 1688980957
transform 1 0 1472 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit3
timestamp 1688980957
transform 1 0 2300 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit4
timestamp 1688980957
transform 1 0 11776 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit5
timestamp 1688980957
transform 1 0 12328 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit6
timestamp 1688980957
transform 1 0 17112 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit7
timestamp 1688980957
transform 1 0 17572 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit8
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit9
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit10
timestamp 1688980957
transform 1 0 2300 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit11
timestamp 1688980957
transform 1 0 3496 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit12
timestamp 1688980957
transform 1 0 8096 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit13
timestamp 1688980957
transform 1 0 9108 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit14
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit15
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit17
timestamp 1688980957
transform 1 0 11684 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit18
timestamp 1688980957
transform 1 0 1840 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit19
timestamp 1688980957
transform 1 0 4876 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit20
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit21
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit22
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit23
timestamp 1688980957
transform 1 0 13892 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit24
timestamp 1688980957
transform 1 0 10856 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit25
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit26
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit27
timestamp 1688980957
transform 1 0 3496 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit28
timestamp 1688980957
transform 1 0 6900 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit29
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit30
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit31
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit0
timestamp 1688980957
transform 1 0 10028 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit1
timestamp 1688980957
transform 1 0 11684 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit2
timestamp 1688980957
transform 1 0 3864 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit3
timestamp 1688980957
transform 1 0 4508 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit4
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit5
timestamp 1688980957
transform 1 0 10028 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit6
timestamp 1688980957
transform 1 0 15088 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit7
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit8
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit9
timestamp 1688980957
transform 1 0 12604 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit10
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit11
timestamp 1688980957
transform 1 0 3404 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit12
timestamp 1688980957
transform 1 0 11868 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit13
timestamp 1688980957
transform 1 0 12512 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit14
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit15
timestamp 1688980957
transform 1 0 18032 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit16
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit17
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit18
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit19
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit20
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit21
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit22
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit23
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit24
timestamp 1688980957
transform 1 0 14628 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit25
timestamp 1688980957
transform 1 0 16928 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit26
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit27
timestamp 1688980957
transform 1 0 6624 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit28
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit29
timestamp 1688980957
transform 1 0 7268 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit30
timestamp 1688980957
transform 1 0 13248 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit31
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit0
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit1
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit2
timestamp 1688980957
transform 1 0 6624 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit3
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit4
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit5
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit6
timestamp 1688980957
transform 1 0 8832 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit7
timestamp 1688980957
transform 1 0 9200 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit8
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit10
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit11
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit12
timestamp 1688980957
transform 1 0 2300 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit13
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit14
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit15
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit17
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit18
timestamp 1688980957
transform 1 0 2208 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit19
timestamp 1688980957
transform 1 0 2300 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit20
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit21
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit22
timestamp 1688980957
transform 1 0 15180 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit23
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit24
timestamp 1688980957
transform 1 0 12420 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit25
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit26
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit27
timestamp 1688980957
transform 1 0 2300 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit28
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit30
timestamp 1688980957
transform 1 0 16192 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit31
timestamp 1688980957
transform 1 0 17572 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit0
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit1
timestamp 1688980957
transform 1 0 17112 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit3
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit4
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit5
timestamp 1688980957
transform 1 0 3496 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit6
timestamp 1688980957
transform 1 0 9568 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit7
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit8
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit9
timestamp 1688980957
transform 1 0 16744 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit10
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit11
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit12
timestamp 1688980957
transform 1 0 1656 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit13
timestamp 1688980957
transform 1 0 2024 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit14
timestamp 1688980957
transform 1 0 6808 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit15
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit16
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit17
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit18
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit19
timestamp 1688980957
transform 1 0 6808 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit20
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit21
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit22
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit23
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit24
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit25
timestamp 1688980957
transform 1 0 14628 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit26
timestamp 1688980957
transform 1 0 4876 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit27
timestamp 1688980957
transform 1 0 5520 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit28
timestamp 1688980957
transform 1 0 4876 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit29
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit30
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit31
timestamp 1688980957
transform 1 0 12604 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit0
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit1
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit2
timestamp 1688980957
transform 1 0 1840 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit3
timestamp 1688980957
transform 1 0 2300 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit4
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit5
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit6
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit7
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit8
timestamp 1688980957
transform 1 0 7452 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit9
timestamp 1688980957
transform 1 0 9200 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit10
timestamp 1688980957
transform 1 0 3956 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit11
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit12
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit13
timestamp 1688980957
transform 1 0 1564 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit14
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit15
timestamp 1688980957
transform 1 0 6440 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit16
timestamp 1688980957
transform 1 0 14536 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit17
timestamp 1688980957
transform 1 0 15364 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit18
timestamp 1688980957
transform 1 0 1840 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit19
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit20
timestamp 1688980957
transform 1 0 1656 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit21
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit22
timestamp 1688980957
transform 1 0 6716 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit23
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit24
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit25
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit26
timestamp 1688980957
transform 1 0 4324 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit27
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit28
timestamp 1688980957
transform 1 0 1656 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit29
timestamp 1688980957
transform 1 0 2208 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit30
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit31
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit0
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit1
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit2
timestamp 1688980957
transform 1 0 13432 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit3
timestamp 1688980957
transform 1 0 14168 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit4
timestamp 1688980957
transform 1 0 12512 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit5
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit6
timestamp 1688980957
transform 1 0 14904 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit7
timestamp 1688980957
transform 1 0 4784 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit8
timestamp 1688980957
transform 1 0 5428 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit9
timestamp 1688980957
transform 1 0 6900 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit10
timestamp 1688980957
transform 1 0 9936 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit11
timestamp 1688980957
transform 1 0 11040 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit12
timestamp 1688980957
transform 1 0 12512 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit13
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit14
timestamp 1688980957
transform 1 0 16928 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit15
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit16
timestamp 1688980957
transform 1 0 9844 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit17
timestamp 1688980957
transform 1 0 11224 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit18
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit19
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit20
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit21
timestamp 1688980957
transform 1 0 9200 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit22
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit23
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit24
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit25
timestamp 1688980957
transform 1 0 9384 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit26
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit27
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit28
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit29
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit30
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit31
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit0
timestamp 1688980957
transform 1 0 8464 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit1
timestamp 1688980957
transform 1 0 9476 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit2
timestamp 1688980957
transform 1 0 9200 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit3
timestamp 1688980957
transform 1 0 4692 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit4
timestamp 1688980957
transform 1 0 5428 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit5
timestamp 1688980957
transform 1 0 6532 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit6
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit7
timestamp 1688980957
transform 1 0 7176 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit8
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit9
timestamp 1688980957
transform 1 0 15180 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit10
timestamp 1688980957
transform 1 0 15916 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit11
timestamp 1688980957
transform 1 0 15640 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit12
timestamp 1688980957
transform 1 0 10304 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit13
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit14
timestamp 1688980957
transform 1 0 4508 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit15
timestamp 1688980957
transform 1 0 4876 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit16
timestamp 1688980957
transform 1 0 11776 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit17
timestamp 1688980957
transform 1 0 13156 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit18
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit19
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit20
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit21
timestamp 1688980957
transform 1 0 11776 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit22
timestamp 1688980957
transform 1 0 4784 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit23
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit24
timestamp 1688980957
transform 1 0 5796 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit25
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit26
timestamp 1688980957
transform 1 0 13892 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit27
timestamp 1688980957
transform 1 0 14168 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit28
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit29
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit30
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit31
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit0
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit1
timestamp 1688980957
transform 1 0 19504 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit2
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit3
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit4
timestamp 1688980957
transform 1 0 22724 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit5
timestamp 1688980957
transform 1 0 22724 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit6
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit7
timestamp 1688980957
transform 1 0 22724 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit8
timestamp 1688980957
transform 1 0 7728 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit9
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit10
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit11
timestamp 1688980957
transform 1 0 1472 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit12
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit13
timestamp 1688980957
transform 1 0 12052 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit14
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit15
timestamp 1688980957
transform 1 0 14168 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit16
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit17
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit19
timestamp 1688980957
transform 1 0 1656 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit20
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit21
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit22
timestamp 1688980957
transform 1 0 6808 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit23
timestamp 1688980957
transform 1 0 7360 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit24
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit25
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit26
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit27
timestamp 1688980957
transform 1 0 1472 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit28
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit29
timestamp 1688980957
transform 1 0 1564 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit30
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit31
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit0
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit1
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit2
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit3
timestamp 1688980957
transform 1 0 18216 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit4
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit5
timestamp 1688980957
transform 1 0 22356 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit6
timestamp 1688980957
transform 1 0 21252 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit7
timestamp 1688980957
transform 1 0 22632 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit8
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit9
timestamp 1688980957
transform 1 0 19964 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit10
timestamp 1688980957
transform 1 0 17572 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit11
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit12
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit13
timestamp 1688980957
transform 1 0 22448 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit14
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit15
timestamp 1688980957
transform 1 0 18584 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit16
timestamp 1688980957
transform 1 0 19872 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit17
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit18
timestamp 1688980957
transform 1 0 19596 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit19
timestamp 1688980957
transform 1 0 17940 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit20
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit21
timestamp 1688980957
transform 1 0 23184 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit22
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit23
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit24
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit25
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit26
timestamp 1688980957
transform 1 0 22724 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit27
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit28
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit29
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit30
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit31
timestamp 1688980957
transform 1 0 19136 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit24
timestamp 1688980957
transform 1 0 19320 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit25
timestamp 1688980957
transform 1 0 19228 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit26
timestamp 1688980957
transform 1 0 22264 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit27
timestamp 1688980957
transform 1 0 20792 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit28
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit29
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit30
timestamp 1688980957
transform 1 0 22448 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit31
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 3680 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 3864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._36_
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._37_
timestamp 1688980957
transform 1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._38_
timestamp 1688980957
transform 1 0 4692 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._39_
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._40_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._41_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._42_
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._43_
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._44_
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._45_
timestamp 1688980957
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._46_
timestamp 1688980957
transform 1 0 12144 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._47_
timestamp 1688980957
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396
timestamp 1688980957
transform 1 0 8004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397
timestamp 1688980957
transform 1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3
timestamp 1688980957
transform 1 0 14720 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0
timestamp 1688980957
transform 1 0 14996 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399
timestamp 1688980957
transform 1 0 16008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400
timestamp 1688980957
transform 1 0 6348 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401
timestamp 1688980957
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2
timestamp 1688980957
transform 1 0 6900 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402
timestamp 1688980957
transform 1 0 14628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1
timestamp 1688980957
transform 1 0 2852 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404
timestamp 1688980957
transform 1 0 4416 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405
timestamp 1688980957
transform 1 0 13156 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2
timestamp 1688980957
transform 1 0 11776 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3
timestamp 1688980957
transform 1 0 17112 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0
timestamp 1688980957
transform 1 0 11224 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1
timestamp 1688980957
transform 1 0 2576 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2
timestamp 1688980957
transform 1 0 10304 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0
timestamp 1688980957
transform 1 0 12788 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1
timestamp 1688980957
transform 1 0 2668 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2
timestamp 1688980957
transform 1 0 9936 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0
timestamp 1688980957
transform 1 0 11316 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1
timestamp 1688980957
transform 1 0 4324 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2
timestamp 1688980957
transform 1 0 9844 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3
timestamp 1688980957
transform 1 0 15732 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2
timestamp 1688980957
transform 1 0 11776 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3
timestamp 1688980957
transform 1 0 16652 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406
timestamp 1688980957
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407
timestamp 1688980957
transform 1 0 3864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1
timestamp 1688980957
transform 1 0 1748 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2
timestamp 1688980957
transform 1 0 9844 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408
timestamp 1688980957
transform 1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2
timestamp 1688980957
transform 1 0 4784 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6
timestamp 1688980957
transform 1 0 8464 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0
timestamp 1688980957
transform 1 0 11316 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2
timestamp 1688980957
transform 1 0 8740 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4
timestamp 1688980957
transform 1 0 11316 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5
timestamp 1688980957
transform 1 0 3220 0 -1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6
timestamp 1688980957
transform 1 0 8004 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10
timestamp 1688980957
transform 1 0 7268 0 -1 40256
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11
timestamp 1688980957
transform 1 0 13432 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13
timestamp 1688980957
transform 1 0 3312 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14
timestamp 1688980957
transform 1 0 8924 0 -1 40256
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1
timestamp 1688980957
transform 1 0 1472 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2
timestamp 1688980957
transform 1 0 11408 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0
timestamp 1688980957
transform 1 0 8648 0 -1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1
timestamp 1688980957
transform 1 0 1472 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3
timestamp 1688980957
transform 1 0 6900 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4
timestamp 1688980957
transform 1 0 1564 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6
timestamp 1688980957
transform 1 0 1840 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1
timestamp 1688980957
transform 1 0 4784 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3
timestamp 1688980957
transform 1 0 13892 0 -1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0
timestamp 1688980957
transform 1 0 11408 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1
timestamp 1688980957
transform 1 0 6164 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3
timestamp 1688980957
transform 1 0 14076 0 -1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4
timestamp 1688980957
transform 1 0 15272 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5
timestamp 1688980957
transform 1 0 1748 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6
timestamp 1688980957
transform 1 0 2392 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3
timestamp 1688980957
transform 1 0 6256 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5
timestamp 1688980957
transform 1 0 1748 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6
timestamp 1688980957
transform 1 0 1748 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7
timestamp 1688980957
transform 1 0 8096 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1
timestamp 1688980957
transform 1 0 5428 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2
timestamp 1688980957
transform 1 0 5336 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4
timestamp 1688980957
transform 1 0 16192 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5
timestamp 1688980957
transform 1 0 6808 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8
timestamp 1688980957
transform 1 0 15732 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9
timestamp 1688980957
transform 1 0 6900 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10
timestamp 1688980957
transform 1 0 2852 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2
timestamp 1688980957
transform 1 0 1748 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6
timestamp 1688980957
transform 1 0 3680 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8
timestamp 1688980957
transform 1 0 16376 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9
timestamp 1688980957
transform 1 0 5704 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14
timestamp 1688980957
transform 1 0 2392 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 11040 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 11316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 10580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10488 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9016 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9200 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 6900 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 8280 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6992 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7176 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4324 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5060 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 9292 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 9108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 8832 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6900 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6808 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 17020 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 17296 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16928 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 15548 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 15548 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 15824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14996 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 12788 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 13064 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 7452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7636 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 13892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 12512 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 12788 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 10488 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 10488 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18216 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 4508 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 5152 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 6532 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 6900 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 6624 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 7268 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 7728 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 8004 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 4784 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 5152 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 5520 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 6624 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 6992 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 7360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 7728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 7360 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output189
timestamp 1688980957
transform 1 0 23552 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 23000 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1688980957
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 23736 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1688980957
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 23644 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output200
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 23552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output206
timestamp 1688980957
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output208
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output209
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output211
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output213
timestamp 1688980957
transform 1 0 23552 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output216
timestamp 1688980957
transform 1 0 23460 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output217
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output219
timestamp 1688980957
transform 1 0 23460 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output220
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1688980957
transform 1 0 24196 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1688980957
transform 1 0 24196 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1688980957
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output224
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output226
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1688980957
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output228
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output229
timestamp 1688980957
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1688980957
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output231
timestamp 1688980957
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1688980957
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1688980957
transform 1 0 24196 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1688980957
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output235
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1688980957
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output237
timestamp 1688980957
transform 1 0 24012 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output238
timestamp 1688980957
transform 1 0 23736 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output239
timestamp 1688980957
transform 1 0 23276 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output240
timestamp 1688980957
transform 1 0 23920 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1688980957
transform 1 0 23920 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output242
timestamp 1688980957
transform 1 0 23092 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output243
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output244
timestamp 1688980957
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output245
timestamp 1688980957
transform 1 0 22724 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1688980957
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output247
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1688980957
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output250
timestamp 1688980957
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1688980957
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output252
timestamp 1688980957
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1688980957
transform 1 0 19872 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output254
timestamp 1688980957
transform 1 0 23276 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output255
timestamp 1688980957
transform 1 0 22724 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output256
timestamp 1688980957
transform 1 0 22080 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output257
timestamp 1688980957
transform 1 0 22632 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output258
timestamp 1688980957
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output259
timestamp 1688980957
transform 1 0 23276 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output260
timestamp 1688980957
transform 1 0 21988 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output261
timestamp 1688980957
transform 1 0 23828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output262
timestamp 1688980957
transform 1 0 23184 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output263
timestamp 1688980957
transform 1 0 22172 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output264
timestamp 1688980957
transform 1 0 20792 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1688980957
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output267
timestamp 1688980957
transform 1 0 22172 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output268
timestamp 1688980957
transform 1 0 22724 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output269
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output270
timestamp 1688980957
transform 1 0 22540 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output271
timestamp 1688980957
transform 1 0 20240 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output272
timestamp 1688980957
transform 1 0 21160 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output273
timestamp 1688980957
transform 1 0 2944 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output274
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output275
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output276
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output277
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output278
timestamp 1688980957
transform 1 0 1932 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output279
timestamp 1688980957
transform 1 0 1656 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output280
timestamp 1688980957
transform 1 0 2024 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output282
timestamp 1688980957
transform 1 0 2576 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output283
timestamp 1688980957
transform 1 0 2392 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output284
timestamp 1688980957
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1688980957
transform 1 0 2760 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1688980957
transform 1 0 3956 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output287
timestamp 1688980957
transform 1 0 3956 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output288
timestamp 1688980957
transform 1 0 4416 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output289
timestamp 1688980957
transform 1 0 4508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output290
timestamp 1688980957
transform 1 0 4968 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1688980957
transform 1 0 4784 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output292
timestamp 1688980957
transform 1 0 5152 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output293
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output294
timestamp 1688980957
transform 1 0 7912 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output295
timestamp 1688980957
transform 1 0 8280 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output296
timestamp 1688980957
transform 1 0 8464 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output297
timestamp 1688980957
transform 1 0 9384 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output298
timestamp 1688980957
transform 1 0 9016 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output299
timestamp 1688980957
transform 1 0 9384 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output300
timestamp 1688980957
transform 1 0 5888 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output301
timestamp 1688980957
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output302
timestamp 1688980957
transform 1 0 6624 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output303
timestamp 1688980957
transform 1 0 6624 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output304
timestamp 1688980957
transform 1 0 7176 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output306
timestamp 1688980957
transform 1 0 7176 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output307
timestamp 1688980957
transform 1 0 7544 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output308
timestamp 1688980957
transform 1 0 8280 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output309
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output310
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output311
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output312
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output313
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output314
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output315
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output316
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output317
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output318
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output319
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output320
timestamp 1688980957
transform 1 0 16100 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output321
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output322
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output323
timestamp 1688980957
transform 1 0 11684 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output324
timestamp 1688980957
transform 1 0 8464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output325
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output326
timestamp 1688980957
transform 1 0 12236 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output327
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output328
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output329
timestamp 1688980957
transform 1 0 15548 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output330
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output331
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output332
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output333
timestamp 1688980957
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output334
timestamp 1688980957
transform 1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output335
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output336
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output337
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output338
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output339
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output340
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output341
timestamp 1688980957
transform 1 0 17204 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output342
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output343
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output344
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output345
timestamp 1688980957
transform 1 0 20516 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output346
timestamp 1688980957
transform 1 0 1932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output347
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output348
timestamp 1688980957
transform 1 0 1564 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output349
timestamp 1688980957
transform 1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output350
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output351
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output352
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output353
timestamp 1688980957
transform 1 0 2116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output354
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output355
timestamp 1688980957
transform 1 0 1564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output356
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output357
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output358
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output359
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output360
timestamp 1688980957
transform 1 0 1564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output361
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output362
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output363
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output364
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output365
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output366
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output367
timestamp 1688980957
transform 1 0 1564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output368
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output369
timestamp 1688980957
transform 1 0 2116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output370
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output371
timestamp 1688980957
transform 1 0 3220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output372
timestamp 1688980957
transform 1 0 3772 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output373
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output374
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output375
timestamp 1688980957
transform 1 0 2668 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output376
timestamp 1688980957
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output377
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output378
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output379
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output380
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output381
timestamp 1688980957
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output382
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output383
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output384
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output385
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output386
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output387
timestamp 1688980957
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output388
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output389
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output390
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output391
timestamp 1688980957
transform 1 0 4324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output392
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output393
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 24840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 24840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 24840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 24840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 24840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 24840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 24840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 24840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 24840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 24840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 24840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 24840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 24840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 24840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 24840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 24840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 24840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 24840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 24840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 24840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 24840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 24840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 24840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 24840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 24840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 24840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 24840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 24840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 24840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 24840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 24840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 24840 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 24840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 24840 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 24840 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 24840 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 24840 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 24840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 24840 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 24840 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 24840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 24840 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 24840 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 16100 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 17020 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 17388 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 18124 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 18492 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 18216 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 19136 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 16928 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 17204 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 17480 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 17756 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 18032 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 18308 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 18584 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 18676 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 19504 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 19044 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 19596 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 19688 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 20056 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 20700 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 20884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 22356 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 19780 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 23460 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 23368 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 22356 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 23920 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 23460 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 20240 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 20516 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 20700 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 21712 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 21804 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 21528 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 22172 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 22724 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 22632 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 21896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 23368 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 23736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 23368 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 22448 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 23184 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 23828 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 23920 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 24288 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 25840 9256 26000 9376 0 FreeSans 480 0 0 0 Config_accessC_bit0
port 0 nsew signal tristate
flabel metal3 s 25840 9800 26000 9920 0 FreeSans 480 0 0 0 Config_accessC_bit1
port 1 nsew signal tristate
flabel metal3 s 25840 10344 26000 10464 0 FreeSans 480 0 0 0 Config_accessC_bit2
port 2 nsew signal tristate
flabel metal3 s 25840 10888 26000 11008 0 FreeSans 480 0 0 0 Config_accessC_bit3
port 3 nsew signal tristate
flabel metal3 s 0 17960 160 18080 0 FreeSans 480 0 0 0 E1END[0]
port 4 nsew signal input
flabel metal3 s 0 18232 160 18352 0 FreeSans 480 0 0 0 E1END[1]
port 5 nsew signal input
flabel metal3 s 0 18504 160 18624 0 FreeSans 480 0 0 0 E1END[2]
port 6 nsew signal input
flabel metal3 s 0 18776 160 18896 0 FreeSans 480 0 0 0 E1END[3]
port 7 nsew signal input
flabel metal3 s 0 21224 160 21344 0 FreeSans 480 0 0 0 E2END[0]
port 8 nsew signal input
flabel metal3 s 0 21496 160 21616 0 FreeSans 480 0 0 0 E2END[1]
port 9 nsew signal input
flabel metal3 s 0 21768 160 21888 0 FreeSans 480 0 0 0 E2END[2]
port 10 nsew signal input
flabel metal3 s 0 22040 160 22160 0 FreeSans 480 0 0 0 E2END[3]
port 11 nsew signal input
flabel metal3 s 0 22312 160 22432 0 FreeSans 480 0 0 0 E2END[4]
port 12 nsew signal input
flabel metal3 s 0 22584 160 22704 0 FreeSans 480 0 0 0 E2END[5]
port 13 nsew signal input
flabel metal3 s 0 22856 160 22976 0 FreeSans 480 0 0 0 E2END[6]
port 14 nsew signal input
flabel metal3 s 0 23128 160 23248 0 FreeSans 480 0 0 0 E2END[7]
port 15 nsew signal input
flabel metal3 s 0 19048 160 19168 0 FreeSans 480 0 0 0 E2MID[0]
port 16 nsew signal input
flabel metal3 s 0 19320 160 19440 0 FreeSans 480 0 0 0 E2MID[1]
port 17 nsew signal input
flabel metal3 s 0 19592 160 19712 0 FreeSans 480 0 0 0 E2MID[2]
port 18 nsew signal input
flabel metal3 s 0 19864 160 19984 0 FreeSans 480 0 0 0 E2MID[3]
port 19 nsew signal input
flabel metal3 s 0 20136 160 20256 0 FreeSans 480 0 0 0 E2MID[4]
port 20 nsew signal input
flabel metal3 s 0 20408 160 20528 0 FreeSans 480 0 0 0 E2MID[5]
port 21 nsew signal input
flabel metal3 s 0 20680 160 20800 0 FreeSans 480 0 0 0 E2MID[6]
port 22 nsew signal input
flabel metal3 s 0 20952 160 21072 0 FreeSans 480 0 0 0 E2MID[7]
port 23 nsew signal input
flabel metal3 s 0 27752 160 27872 0 FreeSans 480 0 0 0 E6END[0]
port 24 nsew signal input
flabel metal3 s 0 30472 160 30592 0 FreeSans 480 0 0 0 E6END[10]
port 25 nsew signal input
flabel metal3 s 0 30744 160 30864 0 FreeSans 480 0 0 0 E6END[11]
port 26 nsew signal input
flabel metal3 s 0 28024 160 28144 0 FreeSans 480 0 0 0 E6END[1]
port 27 nsew signal input
flabel metal3 s 0 28296 160 28416 0 FreeSans 480 0 0 0 E6END[2]
port 28 nsew signal input
flabel metal3 s 0 28568 160 28688 0 FreeSans 480 0 0 0 E6END[3]
port 29 nsew signal input
flabel metal3 s 0 28840 160 28960 0 FreeSans 480 0 0 0 E6END[4]
port 30 nsew signal input
flabel metal3 s 0 29112 160 29232 0 FreeSans 480 0 0 0 E6END[5]
port 31 nsew signal input
flabel metal3 s 0 29384 160 29504 0 FreeSans 480 0 0 0 E6END[6]
port 32 nsew signal input
flabel metal3 s 0 29656 160 29776 0 FreeSans 480 0 0 0 E6END[7]
port 33 nsew signal input
flabel metal3 s 0 29928 160 30048 0 FreeSans 480 0 0 0 E6END[8]
port 34 nsew signal input
flabel metal3 s 0 30200 160 30320 0 FreeSans 480 0 0 0 E6END[9]
port 35 nsew signal input
flabel metal3 s 0 23400 160 23520 0 FreeSans 480 0 0 0 EE4END[0]
port 36 nsew signal input
flabel metal3 s 0 26120 160 26240 0 FreeSans 480 0 0 0 EE4END[10]
port 37 nsew signal input
flabel metal3 s 0 26392 160 26512 0 FreeSans 480 0 0 0 EE4END[11]
port 38 nsew signal input
flabel metal3 s 0 26664 160 26784 0 FreeSans 480 0 0 0 EE4END[12]
port 39 nsew signal input
flabel metal3 s 0 26936 160 27056 0 FreeSans 480 0 0 0 EE4END[13]
port 40 nsew signal input
flabel metal3 s 0 27208 160 27328 0 FreeSans 480 0 0 0 EE4END[14]
port 41 nsew signal input
flabel metal3 s 0 27480 160 27600 0 FreeSans 480 0 0 0 EE4END[15]
port 42 nsew signal input
flabel metal3 s 0 23672 160 23792 0 FreeSans 480 0 0 0 EE4END[1]
port 43 nsew signal input
flabel metal3 s 0 23944 160 24064 0 FreeSans 480 0 0 0 EE4END[2]
port 44 nsew signal input
flabel metal3 s 0 24216 160 24336 0 FreeSans 480 0 0 0 EE4END[3]
port 45 nsew signal input
flabel metal3 s 0 24488 160 24608 0 FreeSans 480 0 0 0 EE4END[4]
port 46 nsew signal input
flabel metal3 s 0 24760 160 24880 0 FreeSans 480 0 0 0 EE4END[5]
port 47 nsew signal input
flabel metal3 s 0 25032 160 25152 0 FreeSans 480 0 0 0 EE4END[6]
port 48 nsew signal input
flabel metal3 s 0 25304 160 25424 0 FreeSans 480 0 0 0 EE4END[7]
port 49 nsew signal input
flabel metal3 s 0 25576 160 25696 0 FreeSans 480 0 0 0 EE4END[8]
port 50 nsew signal input
flabel metal3 s 0 25848 160 25968 0 FreeSans 480 0 0 0 EE4END[9]
port 51 nsew signal input
flabel metal3 s 25840 15784 26000 15904 0 FreeSans 480 0 0 0 FAB2RAM_A0_O0
port 52 nsew signal tristate
flabel metal3 s 25840 16328 26000 16448 0 FreeSans 480 0 0 0 FAB2RAM_A0_O1
port 53 nsew signal tristate
flabel metal3 s 25840 16872 26000 16992 0 FreeSans 480 0 0 0 FAB2RAM_A0_O2
port 54 nsew signal tristate
flabel metal3 s 25840 17416 26000 17536 0 FreeSans 480 0 0 0 FAB2RAM_A0_O3
port 55 nsew signal tristate
flabel metal3 s 25840 13608 26000 13728 0 FreeSans 480 0 0 0 FAB2RAM_A1_O0
port 56 nsew signal tristate
flabel metal3 s 25840 14152 26000 14272 0 FreeSans 480 0 0 0 FAB2RAM_A1_O1
port 57 nsew signal tristate
flabel metal3 s 25840 14696 26000 14816 0 FreeSans 480 0 0 0 FAB2RAM_A1_O2
port 58 nsew signal tristate
flabel metal3 s 25840 15240 26000 15360 0 FreeSans 480 0 0 0 FAB2RAM_A1_O3
port 59 nsew signal tristate
flabel metal3 s 25840 11432 26000 11552 0 FreeSans 480 0 0 0 FAB2RAM_C_O0
port 60 nsew signal tristate
flabel metal3 s 25840 11976 26000 12096 0 FreeSans 480 0 0 0 FAB2RAM_C_O1
port 61 nsew signal tristate
flabel metal3 s 25840 12520 26000 12640 0 FreeSans 480 0 0 0 FAB2RAM_C_O2
port 62 nsew signal tristate
flabel metal3 s 25840 13064 26000 13184 0 FreeSans 480 0 0 0 FAB2RAM_C_O3
port 63 nsew signal tristate
flabel metal3 s 25840 24488 26000 24608 0 FreeSans 480 0 0 0 FAB2RAM_D0_O0
port 64 nsew signal tristate
flabel metal3 s 25840 25032 26000 25152 0 FreeSans 480 0 0 0 FAB2RAM_D0_O1
port 65 nsew signal tristate
flabel metal3 s 25840 25576 26000 25696 0 FreeSans 480 0 0 0 FAB2RAM_D0_O2
port 66 nsew signal tristate
flabel metal3 s 25840 26120 26000 26240 0 FreeSans 480 0 0 0 FAB2RAM_D0_O3
port 67 nsew signal tristate
flabel metal3 s 25840 22312 26000 22432 0 FreeSans 480 0 0 0 FAB2RAM_D1_O0
port 68 nsew signal tristate
flabel metal3 s 25840 22856 26000 22976 0 FreeSans 480 0 0 0 FAB2RAM_D1_O1
port 69 nsew signal tristate
flabel metal3 s 25840 23400 26000 23520 0 FreeSans 480 0 0 0 FAB2RAM_D1_O2
port 70 nsew signal tristate
flabel metal3 s 25840 23944 26000 24064 0 FreeSans 480 0 0 0 FAB2RAM_D1_O3
port 71 nsew signal tristate
flabel metal3 s 25840 20136 26000 20256 0 FreeSans 480 0 0 0 FAB2RAM_D2_O0
port 72 nsew signal tristate
flabel metal3 s 25840 20680 26000 20800 0 FreeSans 480 0 0 0 FAB2RAM_D2_O1
port 73 nsew signal tristate
flabel metal3 s 25840 21224 26000 21344 0 FreeSans 480 0 0 0 FAB2RAM_D2_O2
port 74 nsew signal tristate
flabel metal3 s 25840 21768 26000 21888 0 FreeSans 480 0 0 0 FAB2RAM_D2_O3
port 75 nsew signal tristate
flabel metal3 s 25840 17960 26000 18080 0 FreeSans 480 0 0 0 FAB2RAM_D3_O0
port 76 nsew signal tristate
flabel metal3 s 25840 18504 26000 18624 0 FreeSans 480 0 0 0 FAB2RAM_D3_O1
port 77 nsew signal tristate
flabel metal3 s 25840 19048 26000 19168 0 FreeSans 480 0 0 0 FAB2RAM_D3_O2
port 78 nsew signal tristate
flabel metal3 s 25840 19592 26000 19712 0 FreeSans 480 0 0 0 FAB2RAM_D3_O3
port 79 nsew signal tristate
flabel metal3 s 0 31016 160 31136 0 FreeSans 480 0 0 0 FrameData[0]
port 80 nsew signal input
flabel metal3 s 0 33736 160 33856 0 FreeSans 480 0 0 0 FrameData[10]
port 81 nsew signal input
flabel metal3 s 0 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[11]
port 82 nsew signal input
flabel metal3 s 0 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[12]
port 83 nsew signal input
flabel metal3 s 0 34552 160 34672 0 FreeSans 480 0 0 0 FrameData[13]
port 84 nsew signal input
flabel metal3 s 0 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[14]
port 85 nsew signal input
flabel metal3 s 0 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[15]
port 86 nsew signal input
flabel metal3 s 0 35368 160 35488 0 FreeSans 480 0 0 0 FrameData[16]
port 87 nsew signal input
flabel metal3 s 0 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s 0 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[18]
port 89 nsew signal input
flabel metal3 s 0 36184 160 36304 0 FreeSans 480 0 0 0 FrameData[19]
port 90 nsew signal input
flabel metal3 s 0 31288 160 31408 0 FreeSans 480 0 0 0 FrameData[1]
port 91 nsew signal input
flabel metal3 s 0 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[20]
port 92 nsew signal input
flabel metal3 s 0 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[21]
port 93 nsew signal input
flabel metal3 s 0 37000 160 37120 0 FreeSans 480 0 0 0 FrameData[22]
port 94 nsew signal input
flabel metal3 s 0 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[23]
port 95 nsew signal input
flabel metal3 s 0 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[24]
port 96 nsew signal input
flabel metal3 s 0 37816 160 37936 0 FreeSans 480 0 0 0 FrameData[25]
port 97 nsew signal input
flabel metal3 s 0 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[26]
port 98 nsew signal input
flabel metal3 s 0 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[27]
port 99 nsew signal input
flabel metal3 s 0 38632 160 38752 0 FreeSans 480 0 0 0 FrameData[28]
port 100 nsew signal input
flabel metal3 s 0 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 101 nsew signal input
flabel metal3 s 0 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[2]
port 102 nsew signal input
flabel metal3 s 0 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[30]
port 103 nsew signal input
flabel metal3 s 0 39448 160 39568 0 FreeSans 480 0 0 0 FrameData[31]
port 104 nsew signal input
flabel metal3 s 0 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[3]
port 105 nsew signal input
flabel metal3 s 0 32104 160 32224 0 FreeSans 480 0 0 0 FrameData[4]
port 106 nsew signal input
flabel metal3 s 0 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[5]
port 107 nsew signal input
flabel metal3 s 0 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[6]
port 108 nsew signal input
flabel metal3 s 0 32920 160 33040 0 FreeSans 480 0 0 0 FrameData[7]
port 109 nsew signal input
flabel metal3 s 0 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[8]
port 110 nsew signal input
flabel metal3 s 0 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[9]
port 111 nsew signal input
flabel metal3 s 25840 26664 26000 26784 0 FreeSans 480 0 0 0 FrameData_O[0]
port 112 nsew signal tristate
flabel metal3 s 25840 32104 26000 32224 0 FreeSans 480 0 0 0 FrameData_O[10]
port 113 nsew signal tristate
flabel metal3 s 25840 32648 26000 32768 0 FreeSans 480 0 0 0 FrameData_O[11]
port 114 nsew signal tristate
flabel metal3 s 25840 33192 26000 33312 0 FreeSans 480 0 0 0 FrameData_O[12]
port 115 nsew signal tristate
flabel metal3 s 25840 33736 26000 33856 0 FreeSans 480 0 0 0 FrameData_O[13]
port 116 nsew signal tristate
flabel metal3 s 25840 34280 26000 34400 0 FreeSans 480 0 0 0 FrameData_O[14]
port 117 nsew signal tristate
flabel metal3 s 25840 34824 26000 34944 0 FreeSans 480 0 0 0 FrameData_O[15]
port 118 nsew signal tristate
flabel metal3 s 25840 35368 26000 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 119 nsew signal tristate
flabel metal3 s 25840 35912 26000 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 120 nsew signal tristate
flabel metal3 s 25840 36456 26000 36576 0 FreeSans 480 0 0 0 FrameData_O[18]
port 121 nsew signal tristate
flabel metal3 s 25840 37000 26000 37120 0 FreeSans 480 0 0 0 FrameData_O[19]
port 122 nsew signal tristate
flabel metal3 s 25840 27208 26000 27328 0 FreeSans 480 0 0 0 FrameData_O[1]
port 123 nsew signal tristate
flabel metal3 s 25840 37544 26000 37664 0 FreeSans 480 0 0 0 FrameData_O[20]
port 124 nsew signal tristate
flabel metal3 s 25840 38088 26000 38208 0 FreeSans 480 0 0 0 FrameData_O[21]
port 125 nsew signal tristate
flabel metal3 s 25840 38632 26000 38752 0 FreeSans 480 0 0 0 FrameData_O[22]
port 126 nsew signal tristate
flabel metal3 s 25840 39176 26000 39296 0 FreeSans 480 0 0 0 FrameData_O[23]
port 127 nsew signal tristate
flabel metal3 s 25840 39720 26000 39840 0 FreeSans 480 0 0 0 FrameData_O[24]
port 128 nsew signal tristate
flabel metal3 s 25840 40264 26000 40384 0 FreeSans 480 0 0 0 FrameData_O[25]
port 129 nsew signal tristate
flabel metal3 s 25840 40808 26000 40928 0 FreeSans 480 0 0 0 FrameData_O[26]
port 130 nsew signal tristate
flabel metal3 s 25840 41352 26000 41472 0 FreeSans 480 0 0 0 FrameData_O[27]
port 131 nsew signal tristate
flabel metal3 s 25840 41896 26000 42016 0 FreeSans 480 0 0 0 FrameData_O[28]
port 132 nsew signal tristate
flabel metal3 s 25840 42440 26000 42560 0 FreeSans 480 0 0 0 FrameData_O[29]
port 133 nsew signal tristate
flabel metal3 s 25840 27752 26000 27872 0 FreeSans 480 0 0 0 FrameData_O[2]
port 134 nsew signal tristate
flabel metal3 s 25840 42984 26000 43104 0 FreeSans 480 0 0 0 FrameData_O[30]
port 135 nsew signal tristate
flabel metal3 s 25840 43528 26000 43648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 136 nsew signal tristate
flabel metal3 s 25840 28296 26000 28416 0 FreeSans 480 0 0 0 FrameData_O[3]
port 137 nsew signal tristate
flabel metal3 s 25840 28840 26000 28960 0 FreeSans 480 0 0 0 FrameData_O[4]
port 138 nsew signal tristate
flabel metal3 s 25840 29384 26000 29504 0 FreeSans 480 0 0 0 FrameData_O[5]
port 139 nsew signal tristate
flabel metal3 s 25840 29928 26000 30048 0 FreeSans 480 0 0 0 FrameData_O[6]
port 140 nsew signal tristate
flabel metal3 s 25840 30472 26000 30592 0 FreeSans 480 0 0 0 FrameData_O[7]
port 141 nsew signal tristate
flabel metal3 s 25840 31016 26000 31136 0 FreeSans 480 0 0 0 FrameData_O[8]
port 142 nsew signal tristate
flabel metal3 s 25840 31560 26000 31680 0 FreeSans 480 0 0 0 FrameData_O[9]
port 143 nsew signal tristate
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 144 nsew signal input
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 145 nsew signal input
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 146 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 147 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 148 nsew signal input
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 149 nsew signal input
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 150 nsew signal input
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 151 nsew signal input
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 152 nsew signal input
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 153 nsew signal input
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 154 nsew signal input
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 155 nsew signal input
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 156 nsew signal input
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 157 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 158 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 159 nsew signal input
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 160 nsew signal input
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 161 nsew signal input
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 162 nsew signal input
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 163 nsew signal input
flabel metal2 s 20350 44463 20406 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 164 nsew signal tristate
flabel metal2 s 23110 44463 23166 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 165 nsew signal tristate
flabel metal2 s 23386 44463 23442 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 166 nsew signal tristate
flabel metal2 s 23662 44463 23718 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 167 nsew signal tristate
flabel metal2 s 23938 44463 23994 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 168 nsew signal tristate
flabel metal2 s 24214 44463 24270 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 169 nsew signal tristate
flabel metal2 s 24490 44463 24546 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 170 nsew signal tristate
flabel metal2 s 24766 44463 24822 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 171 nsew signal tristate
flabel metal2 s 25042 44463 25098 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 172 nsew signal tristate
flabel metal2 s 25318 44463 25374 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 173 nsew signal tristate
flabel metal2 s 25594 44463 25650 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 174 nsew signal tristate
flabel metal2 s 20626 44463 20682 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 175 nsew signal tristate
flabel metal2 s 20902 44463 20958 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 176 nsew signal tristate
flabel metal2 s 21178 44463 21234 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 177 nsew signal tristate
flabel metal2 s 21454 44463 21510 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 178 nsew signal tristate
flabel metal2 s 21730 44463 21786 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 179 nsew signal tristate
flabel metal2 s 22006 44463 22062 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 180 nsew signal tristate
flabel metal2 s 22282 44463 22338 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 181 nsew signal tristate
flabel metal2 s 22558 44463 22614 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 182 nsew signal tristate
flabel metal2 s 22834 44463 22890 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 183 nsew signal tristate
flabel metal2 s 202 44463 258 44623 0 FreeSans 224 90 0 0 N1BEG[0]
port 184 nsew signal tristate
flabel metal2 s 478 44463 534 44623 0 FreeSans 224 90 0 0 N1BEG[1]
port 185 nsew signal tristate
flabel metal2 s 754 44463 810 44623 0 FreeSans 224 90 0 0 N1BEG[2]
port 186 nsew signal tristate
flabel metal2 s 1030 44463 1086 44623 0 FreeSans 224 90 0 0 N1BEG[3]
port 187 nsew signal tristate
flabel metal2 s 202 0 258 160 0 FreeSans 224 90 0 0 N1END[0]
port 188 nsew signal input
flabel metal2 s 478 0 534 160 0 FreeSans 224 90 0 0 N1END[1]
port 189 nsew signal input
flabel metal2 s 754 0 810 160 0 FreeSans 224 90 0 0 N1END[2]
port 190 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[3]
port 191 nsew signal input
flabel metal2 s 1306 44463 1362 44623 0 FreeSans 224 90 0 0 N2BEG[0]
port 192 nsew signal tristate
flabel metal2 s 1582 44463 1638 44623 0 FreeSans 224 90 0 0 N2BEG[1]
port 193 nsew signal tristate
flabel metal2 s 1858 44463 1914 44623 0 FreeSans 224 90 0 0 N2BEG[2]
port 194 nsew signal tristate
flabel metal2 s 2134 44463 2190 44623 0 FreeSans 224 90 0 0 N2BEG[3]
port 195 nsew signal tristate
flabel metal2 s 2410 44463 2466 44623 0 FreeSans 224 90 0 0 N2BEG[4]
port 196 nsew signal tristate
flabel metal2 s 2686 44463 2742 44623 0 FreeSans 224 90 0 0 N2BEG[5]
port 197 nsew signal tristate
flabel metal2 s 2962 44463 3018 44623 0 FreeSans 224 90 0 0 N2BEG[6]
port 198 nsew signal tristate
flabel metal2 s 3238 44463 3294 44623 0 FreeSans 224 90 0 0 N2BEG[7]
port 199 nsew signal tristate
flabel metal2 s 3514 44463 3570 44623 0 FreeSans 224 90 0 0 N2BEGb[0]
port 200 nsew signal tristate
flabel metal2 s 3790 44463 3846 44623 0 FreeSans 224 90 0 0 N2BEGb[1]
port 201 nsew signal tristate
flabel metal2 s 4066 44463 4122 44623 0 FreeSans 224 90 0 0 N2BEGb[2]
port 202 nsew signal tristate
flabel metal2 s 4342 44463 4398 44623 0 FreeSans 224 90 0 0 N2BEGb[3]
port 203 nsew signal tristate
flabel metal2 s 4618 44463 4674 44623 0 FreeSans 224 90 0 0 N2BEGb[4]
port 204 nsew signal tristate
flabel metal2 s 4894 44463 4950 44623 0 FreeSans 224 90 0 0 N2BEGb[5]
port 205 nsew signal tristate
flabel metal2 s 5170 44463 5226 44623 0 FreeSans 224 90 0 0 N2BEGb[6]
port 206 nsew signal tristate
flabel metal2 s 5446 44463 5502 44623 0 FreeSans 224 90 0 0 N2BEGb[7]
port 207 nsew signal tristate
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 N2END[0]
port 208 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 N2END[1]
port 209 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2END[2]
port 210 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2END[3]
port 211 nsew signal input
flabel metal2 s 4618 0 4674 160 0 FreeSans 224 90 0 0 N2END[4]
port 212 nsew signal input
flabel metal2 s 4894 0 4950 160 0 FreeSans 224 90 0 0 N2END[5]
port 213 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2END[6]
port 214 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[7]
port 215 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 N2MID[0]
port 216 nsew signal input
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 N2MID[1]
port 217 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N2MID[2]
port 218 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[3]
port 219 nsew signal input
flabel metal2 s 2410 0 2466 160 0 FreeSans 224 90 0 0 N2MID[4]
port 220 nsew signal input
flabel metal2 s 2686 0 2742 160 0 FreeSans 224 90 0 0 N2MID[5]
port 221 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[6]
port 222 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[7]
port 223 nsew signal input
flabel metal2 s 5722 44463 5778 44623 0 FreeSans 224 90 0 0 N4BEG[0]
port 224 nsew signal tristate
flabel metal2 s 8482 44463 8538 44623 0 FreeSans 224 90 0 0 N4BEG[10]
port 225 nsew signal tristate
flabel metal2 s 8758 44463 8814 44623 0 FreeSans 224 90 0 0 N4BEG[11]
port 226 nsew signal tristate
flabel metal2 s 9034 44463 9090 44623 0 FreeSans 224 90 0 0 N4BEG[12]
port 227 nsew signal tristate
flabel metal2 s 9310 44463 9366 44623 0 FreeSans 224 90 0 0 N4BEG[13]
port 228 nsew signal tristate
flabel metal2 s 9586 44463 9642 44623 0 FreeSans 224 90 0 0 N4BEG[14]
port 229 nsew signal tristate
flabel metal2 s 9862 44463 9918 44623 0 FreeSans 224 90 0 0 N4BEG[15]
port 230 nsew signal tristate
flabel metal2 s 5998 44463 6054 44623 0 FreeSans 224 90 0 0 N4BEG[1]
port 231 nsew signal tristate
flabel metal2 s 6274 44463 6330 44623 0 FreeSans 224 90 0 0 N4BEG[2]
port 232 nsew signal tristate
flabel metal2 s 6550 44463 6606 44623 0 FreeSans 224 90 0 0 N4BEG[3]
port 233 nsew signal tristate
flabel metal2 s 6826 44463 6882 44623 0 FreeSans 224 90 0 0 N4BEG[4]
port 234 nsew signal tristate
flabel metal2 s 7102 44463 7158 44623 0 FreeSans 224 90 0 0 N4BEG[5]
port 235 nsew signal tristate
flabel metal2 s 7378 44463 7434 44623 0 FreeSans 224 90 0 0 N4BEG[6]
port 236 nsew signal tristate
flabel metal2 s 7654 44463 7710 44623 0 FreeSans 224 90 0 0 N4BEG[7]
port 237 nsew signal tristate
flabel metal2 s 7930 44463 7986 44623 0 FreeSans 224 90 0 0 N4BEG[8]
port 238 nsew signal tristate
flabel metal2 s 8206 44463 8262 44623 0 FreeSans 224 90 0 0 N4BEG[9]
port 239 nsew signal tristate
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N4END[0]
port 240 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 241 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[11]
port 242 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N4END[12]
port 243 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N4END[13]
port 244 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[14]
port 245 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[15]
port 246 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N4END[1]
port 247 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N4END[2]
port 248 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N4END[3]
port 249 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 250 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N4END[5]
port 251 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N4END[6]
port 252 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N4END[7]
port 253 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N4END[8]
port 254 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N4END[9]
port 255 nsew signal input
flabel metal3 s 25840 7080 26000 7200 0 FreeSans 480 0 0 0 RAM2FAB_D0_I0
port 256 nsew signal input
flabel metal3 s 25840 7624 26000 7744 0 FreeSans 480 0 0 0 RAM2FAB_D0_I1
port 257 nsew signal input
flabel metal3 s 25840 8168 26000 8288 0 FreeSans 480 0 0 0 RAM2FAB_D0_I2
port 258 nsew signal input
flabel metal3 s 25840 8712 26000 8832 0 FreeSans 480 0 0 0 RAM2FAB_D0_I3
port 259 nsew signal input
flabel metal3 s 25840 4904 26000 5024 0 FreeSans 480 0 0 0 RAM2FAB_D1_I0
port 260 nsew signal input
flabel metal3 s 25840 5448 26000 5568 0 FreeSans 480 0 0 0 RAM2FAB_D1_I1
port 261 nsew signal input
flabel metal3 s 25840 5992 26000 6112 0 FreeSans 480 0 0 0 RAM2FAB_D1_I2
port 262 nsew signal input
flabel metal3 s 25840 6536 26000 6656 0 FreeSans 480 0 0 0 RAM2FAB_D1_I3
port 263 nsew signal input
flabel metal3 s 25840 2728 26000 2848 0 FreeSans 480 0 0 0 RAM2FAB_D2_I0
port 264 nsew signal input
flabel metal3 s 25840 3272 26000 3392 0 FreeSans 480 0 0 0 RAM2FAB_D2_I1
port 265 nsew signal input
flabel metal3 s 25840 3816 26000 3936 0 FreeSans 480 0 0 0 RAM2FAB_D2_I2
port 266 nsew signal input
flabel metal3 s 25840 4360 26000 4480 0 FreeSans 480 0 0 0 RAM2FAB_D2_I3
port 267 nsew signal input
flabel metal3 s 25840 552 26000 672 0 FreeSans 480 0 0 0 RAM2FAB_D3_I0
port 268 nsew signal input
flabel metal3 s 25840 1096 26000 1216 0 FreeSans 480 0 0 0 RAM2FAB_D3_I1
port 269 nsew signal input
flabel metal3 s 25840 1640 26000 1760 0 FreeSans 480 0 0 0 RAM2FAB_D3_I2
port 270 nsew signal input
flabel metal3 s 25840 2184 26000 2304 0 FreeSans 480 0 0 0 RAM2FAB_D3_I3
port 271 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 272 nsew signal tristate
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 273 nsew signal tristate
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 274 nsew signal tristate
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 275 nsew signal tristate
flabel metal2 s 10138 44463 10194 44623 0 FreeSans 224 90 0 0 S1END[0]
port 276 nsew signal input
flabel metal2 s 10414 44463 10470 44623 0 FreeSans 224 90 0 0 S1END[1]
port 277 nsew signal input
flabel metal2 s 10690 44463 10746 44623 0 FreeSans 224 90 0 0 S1END[2]
port 278 nsew signal input
flabel metal2 s 10966 44463 11022 44623 0 FreeSans 224 90 0 0 S1END[3]
port 279 nsew signal input
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 280 nsew signal tristate
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 281 nsew signal tristate
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 282 nsew signal tristate
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 283 nsew signal tristate
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 284 nsew signal tristate
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 285 nsew signal tristate
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 286 nsew signal tristate
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 287 nsew signal tristate
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 288 nsew signal tristate
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 289 nsew signal tristate
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 290 nsew signal tristate
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 291 nsew signal tristate
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 292 nsew signal tristate
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 293 nsew signal tristate
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 294 nsew signal tristate
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 295 nsew signal tristate
flabel metal2 s 11242 44463 11298 44623 0 FreeSans 224 90 0 0 S2END[0]
port 296 nsew signal input
flabel metal2 s 11518 44463 11574 44623 0 FreeSans 224 90 0 0 S2END[1]
port 297 nsew signal input
flabel metal2 s 11794 44463 11850 44623 0 FreeSans 224 90 0 0 S2END[2]
port 298 nsew signal input
flabel metal2 s 12070 44463 12126 44623 0 FreeSans 224 90 0 0 S2END[3]
port 299 nsew signal input
flabel metal2 s 12346 44463 12402 44623 0 FreeSans 224 90 0 0 S2END[4]
port 300 nsew signal input
flabel metal2 s 12622 44463 12678 44623 0 FreeSans 224 90 0 0 S2END[5]
port 301 nsew signal input
flabel metal2 s 12898 44463 12954 44623 0 FreeSans 224 90 0 0 S2END[6]
port 302 nsew signal input
flabel metal2 s 13174 44463 13230 44623 0 FreeSans 224 90 0 0 S2END[7]
port 303 nsew signal input
flabel metal2 s 13450 44463 13506 44623 0 FreeSans 224 90 0 0 S2MID[0]
port 304 nsew signal input
flabel metal2 s 13726 44463 13782 44623 0 FreeSans 224 90 0 0 S2MID[1]
port 305 nsew signal input
flabel metal2 s 14002 44463 14058 44623 0 FreeSans 224 90 0 0 S2MID[2]
port 306 nsew signal input
flabel metal2 s 14278 44463 14334 44623 0 FreeSans 224 90 0 0 S2MID[3]
port 307 nsew signal input
flabel metal2 s 14554 44463 14610 44623 0 FreeSans 224 90 0 0 S2MID[4]
port 308 nsew signal input
flabel metal2 s 14830 44463 14886 44623 0 FreeSans 224 90 0 0 S2MID[5]
port 309 nsew signal input
flabel metal2 s 15106 44463 15162 44623 0 FreeSans 224 90 0 0 S2MID[6]
port 310 nsew signal input
flabel metal2 s 15382 44463 15438 44623 0 FreeSans 224 90 0 0 S2MID[7]
port 311 nsew signal input
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 312 nsew signal tristate
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 313 nsew signal tristate
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 314 nsew signal tristate
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 315 nsew signal tristate
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 316 nsew signal tristate
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 317 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 318 nsew signal tristate
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 319 nsew signal tristate
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 320 nsew signal tristate
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 321 nsew signal tristate
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 322 nsew signal tristate
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 323 nsew signal tristate
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 324 nsew signal tristate
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 325 nsew signal tristate
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 326 nsew signal tristate
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 327 nsew signal tristate
flabel metal2 s 15658 44463 15714 44623 0 FreeSans 224 90 0 0 S4END[0]
port 328 nsew signal input
flabel metal2 s 18418 44463 18474 44623 0 FreeSans 224 90 0 0 S4END[10]
port 329 nsew signal input
flabel metal2 s 18694 44463 18750 44623 0 FreeSans 224 90 0 0 S4END[11]
port 330 nsew signal input
flabel metal2 s 18970 44463 19026 44623 0 FreeSans 224 90 0 0 S4END[12]
port 331 nsew signal input
flabel metal2 s 19246 44463 19302 44623 0 FreeSans 224 90 0 0 S4END[13]
port 332 nsew signal input
flabel metal2 s 19522 44463 19578 44623 0 FreeSans 224 90 0 0 S4END[14]
port 333 nsew signal input
flabel metal2 s 19798 44463 19854 44623 0 FreeSans 224 90 0 0 S4END[15]
port 334 nsew signal input
flabel metal2 s 15934 44463 15990 44623 0 FreeSans 224 90 0 0 S4END[1]
port 335 nsew signal input
flabel metal2 s 16210 44463 16266 44623 0 FreeSans 224 90 0 0 S4END[2]
port 336 nsew signal input
flabel metal2 s 16486 44463 16542 44623 0 FreeSans 224 90 0 0 S4END[3]
port 337 nsew signal input
flabel metal2 s 16762 44463 16818 44623 0 FreeSans 224 90 0 0 S4END[4]
port 338 nsew signal input
flabel metal2 s 17038 44463 17094 44623 0 FreeSans 224 90 0 0 S4END[5]
port 339 nsew signal input
flabel metal2 s 17314 44463 17370 44623 0 FreeSans 224 90 0 0 S4END[6]
port 340 nsew signal input
flabel metal2 s 17590 44463 17646 44623 0 FreeSans 224 90 0 0 S4END[7]
port 341 nsew signal input
flabel metal2 s 17866 44463 17922 44623 0 FreeSans 224 90 0 0 S4END[8]
port 342 nsew signal input
flabel metal2 s 18142 44463 18198 44623 0 FreeSans 224 90 0 0 S4END[9]
port 343 nsew signal input
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 UserCLK
port 344 nsew signal input
flabel metal2 s 20074 44463 20130 44623 0 FreeSans 224 90 0 0 UserCLKo
port 345 nsew signal tristate
flabel metal4 s 6878 1040 7198 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 9845 1040 10165 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 15779 1040 16099 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 21713 1040 22033 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal3 s 0 4904 160 5024 0 FreeSans 480 0 0 0 W1BEG[0]
port 348 nsew signal tristate
flabel metal3 s 0 5176 160 5296 0 FreeSans 480 0 0 0 W1BEG[1]
port 349 nsew signal tristate
flabel metal3 s 0 5448 160 5568 0 FreeSans 480 0 0 0 W1BEG[2]
port 350 nsew signal tristate
flabel metal3 s 0 5720 160 5840 0 FreeSans 480 0 0 0 W1BEG[3]
port 351 nsew signal tristate
flabel metal3 s 0 5992 160 6112 0 FreeSans 480 0 0 0 W2BEG[0]
port 352 nsew signal tristate
flabel metal3 s 0 6264 160 6384 0 FreeSans 480 0 0 0 W2BEG[1]
port 353 nsew signal tristate
flabel metal3 s 0 6536 160 6656 0 FreeSans 480 0 0 0 W2BEG[2]
port 354 nsew signal tristate
flabel metal3 s 0 6808 160 6928 0 FreeSans 480 0 0 0 W2BEG[3]
port 355 nsew signal tristate
flabel metal3 s 0 7080 160 7200 0 FreeSans 480 0 0 0 W2BEG[4]
port 356 nsew signal tristate
flabel metal3 s 0 7352 160 7472 0 FreeSans 480 0 0 0 W2BEG[5]
port 357 nsew signal tristate
flabel metal3 s 0 7624 160 7744 0 FreeSans 480 0 0 0 W2BEG[6]
port 358 nsew signal tristate
flabel metal3 s 0 7896 160 8016 0 FreeSans 480 0 0 0 W2BEG[7]
port 359 nsew signal tristate
flabel metal3 s 0 8168 160 8288 0 FreeSans 480 0 0 0 W2BEGb[0]
port 360 nsew signal tristate
flabel metal3 s 0 8440 160 8560 0 FreeSans 480 0 0 0 W2BEGb[1]
port 361 nsew signal tristate
flabel metal3 s 0 8712 160 8832 0 FreeSans 480 0 0 0 W2BEGb[2]
port 362 nsew signal tristate
flabel metal3 s 0 8984 160 9104 0 FreeSans 480 0 0 0 W2BEGb[3]
port 363 nsew signal tristate
flabel metal3 s 0 9256 160 9376 0 FreeSans 480 0 0 0 W2BEGb[4]
port 364 nsew signal tristate
flabel metal3 s 0 9528 160 9648 0 FreeSans 480 0 0 0 W2BEGb[5]
port 365 nsew signal tristate
flabel metal3 s 0 9800 160 9920 0 FreeSans 480 0 0 0 W2BEGb[6]
port 366 nsew signal tristate
flabel metal3 s 0 10072 160 10192 0 FreeSans 480 0 0 0 W2BEGb[7]
port 367 nsew signal tristate
flabel metal3 s 0 14696 160 14816 0 FreeSans 480 0 0 0 W6BEG[0]
port 368 nsew signal tristate
flabel metal3 s 0 17416 160 17536 0 FreeSans 480 0 0 0 W6BEG[10]
port 369 nsew signal tristate
flabel metal3 s 0 17688 160 17808 0 FreeSans 480 0 0 0 W6BEG[11]
port 370 nsew signal tristate
flabel metal3 s 0 14968 160 15088 0 FreeSans 480 0 0 0 W6BEG[1]
port 371 nsew signal tristate
flabel metal3 s 0 15240 160 15360 0 FreeSans 480 0 0 0 W6BEG[2]
port 372 nsew signal tristate
flabel metal3 s 0 15512 160 15632 0 FreeSans 480 0 0 0 W6BEG[3]
port 373 nsew signal tristate
flabel metal3 s 0 15784 160 15904 0 FreeSans 480 0 0 0 W6BEG[4]
port 374 nsew signal tristate
flabel metal3 s 0 16056 160 16176 0 FreeSans 480 0 0 0 W6BEG[5]
port 375 nsew signal tristate
flabel metal3 s 0 16328 160 16448 0 FreeSans 480 0 0 0 W6BEG[6]
port 376 nsew signal tristate
flabel metal3 s 0 16600 160 16720 0 FreeSans 480 0 0 0 W6BEG[7]
port 377 nsew signal tristate
flabel metal3 s 0 16872 160 16992 0 FreeSans 480 0 0 0 W6BEG[8]
port 378 nsew signal tristate
flabel metal3 s 0 17144 160 17264 0 FreeSans 480 0 0 0 W6BEG[9]
port 379 nsew signal tristate
flabel metal3 s 0 10344 160 10464 0 FreeSans 480 0 0 0 WW4BEG[0]
port 380 nsew signal tristate
flabel metal3 s 0 13064 160 13184 0 FreeSans 480 0 0 0 WW4BEG[10]
port 381 nsew signal tristate
flabel metal3 s 0 13336 160 13456 0 FreeSans 480 0 0 0 WW4BEG[11]
port 382 nsew signal tristate
flabel metal3 s 0 13608 160 13728 0 FreeSans 480 0 0 0 WW4BEG[12]
port 383 nsew signal tristate
flabel metal3 s 0 13880 160 14000 0 FreeSans 480 0 0 0 WW4BEG[13]
port 384 nsew signal tristate
flabel metal3 s 0 14152 160 14272 0 FreeSans 480 0 0 0 WW4BEG[14]
port 385 nsew signal tristate
flabel metal3 s 0 14424 160 14544 0 FreeSans 480 0 0 0 WW4BEG[15]
port 386 nsew signal tristate
flabel metal3 s 0 10616 160 10736 0 FreeSans 480 0 0 0 WW4BEG[1]
port 387 nsew signal tristate
flabel metal3 s 0 10888 160 11008 0 FreeSans 480 0 0 0 WW4BEG[2]
port 388 nsew signal tristate
flabel metal3 s 0 11160 160 11280 0 FreeSans 480 0 0 0 WW4BEG[3]
port 389 nsew signal tristate
flabel metal3 s 0 11432 160 11552 0 FreeSans 480 0 0 0 WW4BEG[4]
port 390 nsew signal tristate
flabel metal3 s 0 11704 160 11824 0 FreeSans 480 0 0 0 WW4BEG[5]
port 391 nsew signal tristate
flabel metal3 s 0 11976 160 12096 0 FreeSans 480 0 0 0 WW4BEG[6]
port 392 nsew signal tristate
flabel metal3 s 0 12248 160 12368 0 FreeSans 480 0 0 0 WW4BEG[7]
port 393 nsew signal tristate
flabel metal3 s 0 12520 160 12640 0 FreeSans 480 0 0 0 WW4BEG[8]
port 394 nsew signal tristate
flabel metal3 s 0 12792 160 12912 0 FreeSans 480 0 0 0 WW4BEG[9]
port 395 nsew signal tristate
rlabel via1 13052 43520 13052 43520 0 VGND
rlabel metal1 12972 42976 12972 42976 0 VPWR
rlabel metal1 24012 9146 24012 9146 0 Config_accessC_bit0
rlabel metal1 24656 7514 24656 7514 0 Config_accessC_bit1
rlabel metal1 23368 9146 23368 9146 0 Config_accessC_bit2
rlabel metal3 25572 10948 25572 10948 0 Config_accessC_bit3
rlabel metal3 682 18020 682 18020 0 E1END[0]
rlabel metal3 728 18292 728 18292 0 E1END[1]
rlabel metal3 912 18564 912 18564 0 E1END[2]
rlabel metal3 774 18836 774 18836 0 E1END[3]
rlabel metal3 682 21284 682 21284 0 E2END[0]
rlabel metal3 682 21556 682 21556 0 E2END[1]
rlabel metal3 728 21828 728 21828 0 E2END[2]
rlabel metal3 1694 22100 1694 22100 0 E2END[3]
rlabel metal3 820 22372 820 22372 0 E2END[4]
rlabel metal3 728 22644 728 22644 0 E2END[5]
rlabel metal3 590 22916 590 22916 0 E2END[6]
rlabel metal3 820 23188 820 23188 0 E2END[7]
rlabel metal2 3358 19227 3358 19227 0 E2MID[0]
rlabel metal3 958 19380 958 19380 0 E2MID[1]
rlabel metal3 728 19652 728 19652 0 E2MID[2]
rlabel metal3 498 19924 498 19924 0 E2MID[3]
rlabel metal3 452 20196 452 20196 0 E2MID[4]
rlabel metal3 774 20468 774 20468 0 E2MID[5]
rlabel metal3 728 20740 728 20740 0 E2MID[6]
rlabel metal3 728 21012 728 21012 0 E2MID[7]
rlabel metal3 452 27812 452 27812 0 E6END[0]
rlabel metal2 3450 30379 3450 30379 0 E6END[10]
rlabel metal3 728 30804 728 30804 0 E6END[11]
rlabel metal3 498 28084 498 28084 0 E6END[1]
rlabel metal3 820 28356 820 28356 0 E6END[2]
rlabel metal3 544 28628 544 28628 0 E6END[3]
rlabel metal2 3634 29019 3634 29019 0 E6END[4]
rlabel metal3 728 29172 728 29172 0 E6END[5]
rlabel metal3 636 29444 636 29444 0 E6END[6]
rlabel metal3 544 29716 544 29716 0 E6END[7]
rlabel metal3 820 29988 820 29988 0 E6END[8]
rlabel metal2 3818 30481 3818 30481 0 E6END[9]
rlabel metal3 452 23460 452 23460 0 EE4END[0]
rlabel metal3 1372 26180 1372 26180 0 EE4END[10]
rlabel metal3 636 26452 636 26452 0 EE4END[11]
rlabel metal3 682 26724 682 26724 0 EE4END[12]
rlabel metal3 728 26996 728 26996 0 EE4END[13]
rlabel metal3 659 27268 659 27268 0 EE4END[14]
rlabel metal3 567 27540 567 27540 0 EE4END[15]
rlabel metal3 728 23732 728 23732 0 EE4END[1]
rlabel metal3 774 24004 774 24004 0 EE4END[2]
rlabel metal3 912 24276 912 24276 0 EE4END[3]
rlabel metal3 636 24548 636 24548 0 EE4END[4]
rlabel metal3 1142 24820 1142 24820 0 EE4END[5]
rlabel metal3 682 25092 682 25092 0 EE4END[6]
rlabel metal3 728 25364 728 25364 0 EE4END[7]
rlabel metal3 1441 25636 1441 25636 0 EE4END[8]
rlabel metal2 3542 26129 3542 26129 0 EE4END[9]
rlabel metal2 24150 15759 24150 15759 0 FAB2RAM_A0_O0
rlabel metal3 25572 16388 25572 16388 0 FAB2RAM_A0_O1
rlabel metal3 25020 16932 25020 16932 0 FAB2RAM_A0_O2
rlabel metal1 24380 17306 24380 17306 0 FAB2RAM_A0_O3
rlabel metal3 25158 13668 25158 13668 0 FAB2RAM_A1_O0
rlabel metal3 25526 14212 25526 14212 0 FAB2RAM_A1_O1
rlabel metal3 24974 14756 24974 14756 0 FAB2RAM_A1_O2
rlabel metal1 24748 14246 24748 14246 0 FAB2RAM_A1_O3
rlabel metal3 24882 11492 24882 11492 0 FAB2RAM_C_O0
rlabel metal3 25572 12036 25572 12036 0 FAB2RAM_C_O1
rlabel metal3 25066 12580 25066 12580 0 FAB2RAM_C_O2
rlabel metal3 25687 13124 25687 13124 0 FAB2RAM_C_O3
rlabel metal3 25158 24548 25158 24548 0 FAB2RAM_D0_O0
rlabel metal3 25526 25092 25526 25092 0 FAB2RAM_D0_O1
rlabel metal3 25158 25636 25158 25636 0 FAB2RAM_D0_O2
rlabel metal3 25526 26180 25526 26180 0 FAB2RAM_D0_O3
rlabel metal1 24472 21658 24472 21658 0 FAB2RAM_D1_O0
rlabel metal3 25526 22916 25526 22916 0 FAB2RAM_D1_O1
rlabel metal3 25158 23460 25158 23460 0 FAB2RAM_D1_O2
rlabel metal3 25526 24004 25526 24004 0 FAB2RAM_D1_O3
rlabel metal1 24012 20026 24012 20026 0 FAB2RAM_D2_O0
rlabel metal1 24794 19278 24794 19278 0 FAB2RAM_D2_O1
rlabel metal3 24882 21284 24882 21284 0 FAB2RAM_D2_O2
rlabel metal3 25526 21828 25526 21828 0 FAB2RAM_D2_O3
rlabel metal3 25158 18020 25158 18020 0 FAB2RAM_D3_O0
rlabel metal3 25526 18564 25526 18564 0 FAB2RAM_D3_O1
rlabel metal3 24882 19108 24882 19108 0 FAB2RAM_D3_O2
rlabel metal1 24748 18598 24748 18598 0 FAB2RAM_D3_O3
rlabel metal3 1464 31076 1464 31076 0 FrameData[0]
rlabel metal3 590 33796 590 33796 0 FrameData[10]
rlabel metal2 3450 34867 3450 34867 0 FrameData[11]
rlabel metal3 1441 34340 1441 34340 0 FrameData[12]
rlabel metal3 452 34612 452 34612 0 FrameData[13]
rlabel metal3 774 34884 774 34884 0 FrameData[14]
rlabel metal2 3818 35649 3818 35649 0 FrameData[15]
rlabel metal3 866 35428 866 35428 0 FrameData[16]
rlabel metal2 2898 36431 2898 36431 0 FrameData[17]
rlabel via2 3450 35989 3450 35989 0 FrameData[18]
rlabel metal3 728 36244 728 36244 0 FrameData[19]
rlabel metal3 774 31348 774 31348 0 FrameData[1]
rlabel metal3 590 36516 590 36516 0 FrameData[20]
rlabel metal2 3266 38369 3266 38369 0 FrameData[21]
rlabel metal2 3910 37247 3910 37247 0 FrameData[22]
rlabel metal3 4508 37400 4508 37400 0 FrameData[23]
rlabel metal3 774 37604 774 37604 0 FrameData[24]
rlabel metal3 452 37876 452 37876 0 FrameData[25]
rlabel metal3 682 38148 682 38148 0 FrameData[26]
rlabel metal2 3082 38675 3082 38675 0 FrameData[27]
rlabel metal3 1441 38692 1441 38692 0 FrameData[28]
rlabel metal2 2806 39695 2806 39695 0 FrameData[29]
rlabel metal3 1970 31620 1970 31620 0 FrameData[2]
rlabel metal3 774 39236 774 39236 0 FrameData[30]
rlabel metal3 475 39508 475 39508 0 FrameData[31]
rlabel metal3 1740 31892 1740 31892 0 FrameData[3]
rlabel metal3 682 32164 682 32164 0 FrameData[4]
rlabel metal3 728 32436 728 32436 0 FrameData[5]
rlabel metal2 2806 33337 2806 33337 0 FrameData[6]
rlabel metal3 820 32980 820 32980 0 FrameData[7]
rlabel metal2 2898 33660 2898 33660 0 FrameData[8]
rlabel metal3 728 33524 728 33524 0 FrameData[9]
rlabel metal3 25158 26724 25158 26724 0 FrameData_O[0]
rlabel metal3 25158 32164 25158 32164 0 FrameData_O[10]
rlabel metal3 25572 32708 25572 32708 0 FrameData_O[11]
rlabel metal3 25158 33252 25158 33252 0 FrameData_O[12]
rlabel metal3 25572 33796 25572 33796 0 FrameData_O[13]
rlabel metal3 25503 34340 25503 34340 0 FrameData_O[14]
rlabel metal3 25572 34884 25572 34884 0 FrameData_O[15]
rlabel metal3 25158 35428 25158 35428 0 FrameData_O[16]
rlabel metal3 25526 35972 25526 35972 0 FrameData_O[17]
rlabel metal3 25158 36516 25158 36516 0 FrameData_O[18]
rlabel metal3 25503 37060 25503 37060 0 FrameData_O[19]
rlabel metal3 25526 27268 25526 27268 0 FrameData_O[1]
rlabel metal3 25158 37604 25158 37604 0 FrameData_O[20]
rlabel metal3 25572 38148 25572 38148 0 FrameData_O[21]
rlabel metal3 25158 38692 25158 38692 0 FrameData_O[22]
rlabel metal3 25572 39236 25572 39236 0 FrameData_O[23]
rlabel metal3 25158 39780 25158 39780 0 FrameData_O[24]
rlabel metal3 25526 40324 25526 40324 0 FrameData_O[25]
rlabel metal3 24790 40868 24790 40868 0 FrameData_O[26]
rlabel metal3 25526 41412 25526 41412 0 FrameData_O[27]
rlabel metal3 25020 41956 25020 41956 0 FrameData_O[28]
rlabel metal3 25526 42500 25526 42500 0 FrameData_O[29]
rlabel metal3 25158 27812 25158 27812 0 FrameData_O[2]
rlabel metal1 24748 41786 24748 41786 0 FrameData_O[30]
rlabel metal1 23184 42330 23184 42330 0 FrameData_O[31]
rlabel metal3 25526 28356 25526 28356 0 FrameData_O[3]
rlabel metal3 25158 28900 25158 28900 0 FrameData_O[4]
rlabel metal3 25526 29444 25526 29444 0 FrameData_O[5]
rlabel metal3 25158 29988 25158 29988 0 FrameData_O[6]
rlabel metal3 25526 30532 25526 30532 0 FrameData_O[7]
rlabel metal3 25158 31076 25158 31076 0 FrameData_O[8]
rlabel metal1 24702 31790 24702 31790 0 FrameData_O[9]
rlabel metal1 19964 1938 19964 1938 0 FrameStrobe[0]
rlabel metal2 23138 1010 23138 1010 0 FrameStrobe[10]
rlabel metal2 23414 704 23414 704 0 FrameStrobe[11]
rlabel metal1 22011 1938 22011 1938 0 FrameStrobe[12]
rlabel metal2 23966 636 23966 636 0 FrameStrobe[13]
rlabel metal2 20010 3247 20010 3247 0 FrameStrobe[14]
rlabel metal2 24518 942 24518 942 0 FrameStrobe[15]
rlabel metal2 24695 68 24695 68 0 FrameStrobe[16]
rlabel metal1 19596 2958 19596 2958 0 FrameStrobe[17]
rlabel metal2 18814 1700 18814 1700 0 FrameStrobe[18]
rlabel metal2 21206 1122 21206 1122 0 FrameStrobe[19]
rlabel metal2 20654 704 20654 704 0 FrameStrobe[1]
rlabel metal2 20838 1003 20838 1003 0 FrameStrobe[2]
rlabel metal2 21206 279 21206 279 0 FrameStrobe[3]
rlabel metal2 21383 68 21383 68 0 FrameStrobe[4]
rlabel metal1 19504 2414 19504 2414 0 FrameStrobe[5]
rlabel metal2 22034 364 22034 364 0 FrameStrobe[6]
rlabel metal1 22264 5202 22264 5202 0 FrameStrobe[7]
rlabel metal2 22685 68 22685 68 0 FrameStrobe[8]
rlabel metal1 20930 2414 20930 2414 0 FrameStrobe[9]
rlabel metal1 20240 43418 20240 43418 0 FrameStrobe_O[0]
rlabel metal2 23138 43972 23138 43972 0 FrameStrobe_O[10]
rlabel metal1 23276 41242 23276 41242 0 FrameStrobe_O[11]
rlabel metal1 22402 41650 22402 41650 0 FrameStrobe_O[12]
rlabel metal1 23368 41786 23368 41786 0 FrameStrobe_O[13]
rlabel metal1 24196 42670 24196 42670 0 FrameStrobe_O[14]
rlabel metal1 24104 42330 24104 42330 0 FrameStrobe_O[15]
rlabel metal1 23000 42602 23000 42602 0 FrameStrobe_O[16]
rlabel metal1 24656 41242 24656 41242 0 FrameStrobe_O[17]
rlabel metal1 24426 41718 24426 41718 0 FrameStrobe_O[18]
rlabel metal1 22816 42330 22816 42330 0 FrameStrobe_O[19]
rlabel metal2 20654 43972 20654 43972 0 FrameStrobe_O[1]
rlabel metal1 21252 43146 21252 43146 0 FrameStrobe_O[2]
rlabel metal1 21620 43418 21620 43418 0 FrameStrobe_O[3]
rlabel metal2 21482 43938 21482 43938 0 FrameStrobe_O[4]
rlabel metal2 21758 44176 21758 44176 0 FrameStrobe_O[5]
rlabel metal2 21942 42721 21942 42721 0 FrameStrobe_O[6]
rlabel metal2 22310 43530 22310 43530 0 FrameStrobe_O[7]
rlabel metal1 20700 43146 20700 43146 0 FrameStrobe_O[8]
rlabel metal1 21666 42228 21666 42228 0 FrameStrobe_O[9]
rlabel metal1 24058 9554 24058 9554 0 Inst_Config_accessConfig_access.ConfigBits\[0\]
rlabel metal1 24518 8500 24518 8500 0 Inst_Config_accessConfig_access.ConfigBits\[1\]
rlabel metal1 22678 10540 22678 10540 0 Inst_Config_accessConfig_access.ConfigBits\[2\]
rlabel metal1 23644 11322 23644 11322 0 Inst_Config_accessConfig_access.ConfigBits\[3\]
rlabel metal2 19826 15164 19826 15164 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21942 17000 21942 17000 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal2 23782 18258 23782 18258 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 22494 19380 22494 19380 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel via1 18165 16150 18165 16150 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 20316 17578 20316 17578 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 14582 18360 14582 18360 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 20920 19822 20920 19822 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19826 16116 19826 16116 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 22678 17612 22678 17612 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23552 16558 23552 16558 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal2 22126 20230 22126 20230 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18860 15674 18860 15674 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 20010 15436 20010 15436 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 19550 15436 19550 15436 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19826 14926 19826 14926 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 22218 17476 22218 17476 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21666 17204 21666 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 22310 17136 22310 17136 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21574 16694 21574 16694 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 24334 17204 24334 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23138 16422 23138 16422 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 24288 16082 24288 16082 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23920 16014 23920 16014 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21850 19380 21850 19380 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal2 22678 19822 22678 19822 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 22080 19142 22080 19142 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 22494 19278 22494 19278 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 19090 13498 19090 13498 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 23920 14994 23920 14994 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal2 23782 21012 23782 21012 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20378 19346 20378 19346 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel via1 17429 14994 17429 14994 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\]
rlabel metal4 17204 17476 17204 17476 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 15318 25194 15318 25194 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18400 19822 18400 19822 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 18722 14382 18722 14382 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23322 14348 23322 14348 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23368 19346 23368 19346 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20424 18734 20424 18734 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18446 14348 18446 14348 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19642 13940 19642 13940 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18584 13498 18584 13498 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19182 13362 19182 13362 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23414 15028 23414 15028 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel viali 22949 13912 22949 13912 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23920 14858 23920 14858 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 22862 13804 22862 13804 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 22494 20740 22494 20740 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23368 19210 23368 19210 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 24242 20604 24242 20604 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23966 20366 23966 20366 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 19412 18734 19412 18734 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20240 18870 20240 18870 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 20010 18938 20010 18938 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20930 19278 20930 19278 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 22494 14688 22494 14688 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20746 31178 20746 31178 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23046 37706 23046 37706 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 21022 16422 21022 16422 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 20465 15062 20465 15062 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 19596 31790 19596 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 21344 38930 21344 38930 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 19258 17578 19258 17578 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 22352 14382 22352 14382 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20700 31790 20700 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23414 38318 23414 38318 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20700 17170 20700 17170 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21482 14348 21482 14348 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 22632 14382 22632 14382 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21758 14518 21758 14518 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22356 14450 22356 14450 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20102 31824 20102 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20700 31926 20700 31926 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 20332 31790 20332 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21114 30906 21114 30906 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 22126 38522 22126 38522 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 22954 38284 22954 38284 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 23138 37842 23138 37842 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23368 37910 23368 37910 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20102 17204 20102 17204 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20838 16116 20838 16116 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 20746 16762 20746 16762 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 21160 16218 21160 16218 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 22218 29716 22218 29716 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20976 28050 20976 28050 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18814 35666 18814 35666 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19780 28934 19780 28934 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 19862 30226 19862 30226 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 19627 28050 19627 28050 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 17618 36754 17618 36754 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18262 28526 18262 28526 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\]
rlabel metal2 22310 30362 22310 30362 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20976 27438 20976 27438 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 18676 36142 18676 36142 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 19228 28186 19228 28186 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21666 29580 21666 29580 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 22586 30090 22586 30090 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21942 29682 21942 29682 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22402 29682 22402 29682 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20010 27608 20010 27608 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21206 27642 21206 27642 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 21206 27914 21206 27914 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21574 27982 21574 27982 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18078 35054 18078 35054 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19550 35700 19550 35700 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18676 35258 18676 35258 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19366 35598 19366 35598 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 19274 28560 19274 28560 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19320 28730 19320 28730 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19550 28594 19550 28594 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 19918 28662 19918 28662 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 21666 22270 21666 22270 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 23460 25262 23460 25262 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18676 33490 18676 33490 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19826 25874 19826 25874 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 20822 23018 20822 23018 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\]
rlabel metal2 4186 24735 4186 24735 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 17424 33490 17424 33490 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18998 26758 18998 26758 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 22356 21998 22356 21998 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23414 25398 23414 25398 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19550 33558 19550 33558 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 19688 25262 19688 25262 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21436 22746 21436 22746 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 22448 22134 22448 22134 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 22172 22202 22172 22202 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21942 22406 21942 22406 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23046 25908 23046 25908 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23552 26010 23552 26010 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23322 25466 23322 25466 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23690 25398 23690 25398 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18170 34000 18170 34000 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 19458 33422 19458 33422 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18814 33524 18814 33524 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 18998 33388 18998 33388 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal2 19274 25738 19274 25738 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19918 25398 19918 25398 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19734 25466 19734 25466 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20378 25806 20378 25806 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20884 21658 20884 21658 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 22678 27404 22678 27404 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20838 33966 20838 33966 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19274 30634 19274 30634 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 19913 21998 19913 21998 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\]
rlabel metal2 9154 27914 9154 27914 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 18998 35054 18998 35054 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 17802 30906 17802 30906 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20792 21862 20792 21862 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 22724 27642 22724 27642 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 21022 34612 21022 34612 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20102 30804 20102 30804 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 20010 20910 20010 20910 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 20746 21488 20746 21488 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 20930 21114 20930 21114 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21482 21454 21482 21454 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 22908 27438 22908 27438 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal2 23506 27642 23506 27642 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22954 27574 22954 27574 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23184 27506 23184 27506 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20102 34578 20102 34578 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 21574 34034 21574 34034 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 21114 34340 21114 34340 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21390 34034 21390 34034 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18538 31280 18538 31280 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19872 30702 19872 30702 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18998 30906 18998 30906 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 19642 30770 19642 30770 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20010 23494 20010 23494 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 23184 21964 23184 21964 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23230 33490 23230 33490 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 21390 25670 21390 25670 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18068 23698 18068 23698 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\]
rlabel metal2 6118 24429 6118 24429 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 17250 33320 17250 33320 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 20138 24786 20138 24786 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19504 23834 19504 23834 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23874 23290 23874 23290 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23046 33626 23046 33626 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 22034 24718 22034 24718 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19274 23120 19274 23120 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20010 24140 20010 24140 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19550 23154 19550 23154 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19918 23222 19918 23222 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23506 23732 23506 23732 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23414 23664 23414 23664 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23414 22202 23414 22202 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23368 22066 23368 22066 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 22218 33082 22218 33082 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23874 33422 23874 33422 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 22862 33082 22862 33082 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23690 33422 23690 33422 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20930 24140 20930 24140 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21712 24922 21712 24922 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21252 24378 21252 24378 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 21574 24718 21574 24718 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 20378 7378 20378 7378 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20194 10778 20194 10778 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23414 7514 23414 7514 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 22172 9554 22172 9554 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 19550 8024 19550 8024 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
rlabel metal2 13846 11220 13846 11220 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
rlabel metal1 1978 17102 1978 17102 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
rlabel metal1 19734 9384 19734 9384 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
rlabel metal1 22034 7446 22034 7446 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\]
rlabel metal2 21114 10166 21114 10166 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 22494 7820 22494 7820 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 22586 9146 22586 9146 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 20516 6970 20516 6970 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 21206 6970 21206 6970 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 20332 7514 20332 7514 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 21114 7412 21114 7412 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20240 10030 20240 10030 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20884 10642 20884 10642 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 20240 10234 20240 10234 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 20746 10948 20746 10948 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 23920 7242 23920 7242 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 24150 6732 24150 6732 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 22862 8058 22862 8058 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal2 24058 7650 24058 7650 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21850 9520 21850 9520 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 22310 9622 22310 9622 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 22126 8976 22126 8976 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 22678 8500 22678 8500 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 19596 7854 19596 7854 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21942 11764 21942 11764 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23506 2550 23506 2550 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 23276 6290 23276 6290 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal2 16836 8058 16836 8058 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
rlabel metal2 2024 14382 2024 14382 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
rlabel metal2 2622 5355 2622 5355 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
rlabel metal1 21114 7208 21114 7208 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
rlabel metal1 19734 7514 19734 7514 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 23506 12308 23506 12308 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 24380 5338 24380 5338 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 21850 5882 21850 5882 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\]
rlabel metal2 18630 7412 18630 7412 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20056 8058 20056 8058 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19458 7888 19458 7888 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19918 7786 19918 7786 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 22770 12036 22770 12036 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23276 12206 23276 12206 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22402 11764 22402 11764 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 22862 11730 22862 11730 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 24196 3162 24196 3162 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 23552 2414 23552 2414 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 23690 5712 23690 5712 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23736 2482 23736 2482 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel viali 21206 6292 21206 6292 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 23414 6188 23414 6188 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21252 6086 21252 6086 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 23046 6426 23046 6426 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 19412 5202 19412 5202 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21022 5151 21022 5151 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18998 11186 18998 11186 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19274 12784 19274 12784 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 15226 11084 15226 11084 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\]
rlabel metal2 20194 4862 20194 4862 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\]
rlabel metal1 1702 17068 1702 17068 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\]
rlabel metal2 20194 13090 20194 13090 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\]
rlabel metal1 20746 3706 20746 3706 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 21574 4250 21574 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 19136 10030 19136 10030 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 21574 12886 21574 12886 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 19504 3978 19504 3978 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19734 4556 19734 4556 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19182 4726 19182 4726 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 19550 5032 19550 5032 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23920 3366 23920 3366 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21390 4522 21390 4522 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 21068 4726 21068 4726 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21436 4794 21436 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 17940 10030 17940 10030 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19182 9894 19182 9894 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18538 10234 18538 10234 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19228 11050 19228 11050 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20746 12614 20746 12614 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21482 12682 21482 12682 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19918 13328 19918 13328 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20286 13192 20286 13192 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 18262 6086 18262 6086 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 23598 13396 23598 13396 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 22632 3366 22632 3366 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20102 4216 20102 4216 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 17940 6426 17940 6426 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\]
rlabel metal1 1380 14382 1380 14382 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\]
rlabel metal1 1150 10030 1150 10030 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\]
rlabel metal3 21137 2516 21137 2516 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\]
rlabel metal2 18814 4964 18814 4964 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 22494 13260 22494 13260 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 22770 4522 22770 4522 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 24058 2890 24058 2890 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 17848 3978 17848 3978 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18538 5270 18538 5270 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 18170 5746 18170 5746 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 18446 5780 18446 5780 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23000 11526 23000 11526 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 22448 13498 22448 13498 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23092 13498 23092 13498 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23552 13974 23552 13974 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal3 18998 6868 18998 6868 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23000 1258 23000 1258 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 22402 5508 22402 5508 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23966 3978 23966 3978 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18538 3672 18538 3672 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20332 4590 20332 4590 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 23736 2414 23736 2414 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20976 1870 20976 1870 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 12880 20366 12880 20366 0 Inst_RAM_IO_ConfigMem.ConfigBits\[100\]
rlabel metal2 13570 20230 13570 20230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
rlabel metal2 5198 22236 5198 22236 0 Inst_RAM_IO_ConfigMem.ConfigBits\[102\]
rlabel metal1 5474 21658 5474 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
rlabel metal1 9200 18394 9200 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[104\]
rlabel metal1 9614 18734 9614 18734 0 Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
rlabel metal2 14490 18972 14490 18972 0 Inst_RAM_IO_ConfigMem.ConfigBits\[106\]
rlabel metal1 14950 18394 14950 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
rlabel metal1 13478 27880 13478 27880 0 Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
rlabel metal2 14030 28220 14030 28220 0 Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
rlabel metal1 15916 25874 15916 25874 0 Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
rlabel metal2 5842 24990 5842 24990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
rlabel metal2 6394 24684 6394 24684 0 Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
rlabel metal1 7912 23494 7912 23494 0 Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
rlabel metal1 11086 30362 11086 30362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
rlabel metal1 11914 30770 11914 30770 0 Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
rlabel metal1 13754 31314 13754 31314 0 Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
rlabel metal2 17342 22338 17342 22338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
rlabel metal1 17940 21114 17940 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
rlabel metal1 18952 20978 18952 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
rlabel metal1 11546 5882 11546 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
rlabel metal1 12190 5814 12190 5814 0 Inst_RAM_IO_ConfigMem.ConfigBits\[121\]
rlabel metal1 4462 17816 4462 17816 0 Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
rlabel metal2 5014 17850 5014 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[123\]
rlabel metal1 9614 11288 9614 11288 0 Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
rlabel metal1 10212 10778 10212 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[125\]
rlabel metal1 13524 4794 13524 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
rlabel metal1 14536 3706 14536 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[127\]
rlabel metal1 9338 6902 9338 6902 0 Inst_RAM_IO_ConfigMem.ConfigBits\[128\]
rlabel metal1 10258 6834 10258 6834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
rlabel metal2 5014 5338 5014 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[130\]
rlabel metal2 5566 4964 5566 4964 0 Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
rlabel metal1 4508 9690 4508 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[132\]
rlabel metal2 5014 10268 5014 10268 0 Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
rlabel metal2 7406 5542 7406 5542 0 Inst_RAM_IO_ConfigMem.ConfigBits\[134\]
rlabel metal1 7360 5882 7360 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
rlabel metal1 15962 5848 15962 5848 0 Inst_RAM_IO_ConfigMem.ConfigBits\[136\]
rlabel metal1 17434 5338 17434 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
rlabel metal2 2438 12070 2438 12070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[138\]
rlabel metal1 3174 12274 3174 12274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
rlabel metal2 2530 4488 2530 4488 0 Inst_RAM_IO_ConfigMem.ConfigBits\[140\]
rlabel metal2 3634 4556 3634 4556 0 Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
rlabel metal1 9062 3638 9062 3638 0 Inst_RAM_IO_ConfigMem.ConfigBits\[142\]
rlabel metal1 10350 3570 10350 3570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
rlabel metal1 9016 5882 9016 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[144\]
rlabel metal2 10258 5780 10258 5780 0 Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
rlabel metal2 5014 6834 5014 6834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[146\]
rlabel metal2 5566 7174 5566 7174 0 Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
rlabel metal1 2392 17102 2392 17102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[148\]
rlabel metal2 2898 17884 2898 17884 0 Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
rlabel metal1 6440 7990 6440 7990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[150\]
rlabel metal2 7498 7684 7498 7684 0 Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
rlabel metal1 15456 4250 15456 4250 0 Inst_RAM_IO_ConfigMem.ConfigBits\[152\]
rlabel metal2 16422 4964 16422 4964 0 Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
rlabel metal1 2438 14552 2438 14552 0 Inst_RAM_IO_ConfigMem.ConfigBits\[154\]
rlabel metal1 3128 14042 3128 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
rlabel metal1 2576 2074 2576 2074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[156\]
rlabel metal1 3128 2618 3128 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
rlabel metal1 8786 3944 8786 3944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[158\]
rlabel metal1 9246 2074 9246 2074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
rlabel metal1 18216 8058 18216 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[160\]
rlabel metal1 17526 8568 17526 8568 0 Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
rlabel metal1 5474 14518 5474 14518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[162\]
rlabel metal1 6026 14042 6026 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
rlabel metal1 2576 9690 2576 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[164\]
rlabel metal2 2990 10081 2990 10081 0 Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
rlabel metal1 8280 8602 8280 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[166\]
rlabel metal1 9062 9146 9062 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
rlabel metal1 15640 11254 15640 11254 0 Inst_RAM_IO_ConfigMem.ConfigBits\[168\]
rlabel metal1 16790 11186 16790 11186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
rlabel metal1 5750 11866 5750 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[170\]
rlabel metal1 6762 12614 6762 12614 0 Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
rlabel metal1 4416 12750 4416 12750 0 Inst_RAM_IO_ConfigMem.ConfigBits\[172\]
rlabel metal1 4738 11866 4738 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
rlabel metal1 10396 13430 10396 13430 0 Inst_RAM_IO_ConfigMem.ConfigBits\[174\]
rlabel metal1 11040 12954 11040 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
rlabel metal1 17388 11866 17388 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[176\]
rlabel metal2 17710 12308 17710 12308 0 Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
rlabel metal1 6164 9690 6164 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[178\]
rlabel metal1 7176 10098 7176 10098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
rlabel metal1 2438 17816 2438 17816 0 Inst_RAM_IO_ConfigMem.ConfigBits\[180\]
rlabel metal2 2990 17850 2990 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
rlabel metal1 8280 12682 8280 12682 0 Inst_RAM_IO_ConfigMem.ConfigBits\[182\]
rlabel metal2 9246 13260 9246 13260 0 Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
rlabel metal1 15962 8024 15962 8024 0 Inst_RAM_IO_ConfigMem.ConfigBits\[184\]
rlabel metal1 16836 7922 16836 7922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
rlabel metal1 7038 14824 7038 14824 0 Inst_RAM_IO_ConfigMem.ConfigBits\[186\]
rlabel metal1 7728 14586 7728 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
rlabel metal1 3036 7310 3036 7310 0 Inst_RAM_IO_ConfigMem.ConfigBits\[188\]
rlabel metal1 3496 6970 3496 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
rlabel metal1 10258 8602 10258 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[190\]
rlabel metal1 10718 9146 10718 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
rlabel metal1 14950 14518 14950 14518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[192\]
rlabel metal1 15594 14042 15594 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
rlabel metal1 6026 39542 6026 39542 0 Inst_RAM_IO_ConfigMem.ConfigBits\[194\]
rlabel metal2 6670 39882 6670 39882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
rlabel metal2 6026 39678 6026 39678 0 Inst_RAM_IO_ConfigMem.ConfigBits\[196\]
rlabel metal1 6992 37978 6992 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
rlabel metal2 13110 13889 13110 13889 0 Inst_RAM_IO_ConfigMem.ConfigBits\[198\]
rlabel metal2 13662 13702 13662 13702 0 Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
rlabel metal1 16698 13498 16698 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[200\]
rlabel metal1 17572 14042 17572 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
rlabel metal1 7590 11322 7590 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[202\]
rlabel metal1 8004 11866 8004 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
rlabel metal1 3680 15946 3680 15946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[204\]
rlabel metal1 4784 15674 4784 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
rlabel metal1 9660 15606 9660 15606 0 Inst_RAM_IO_ConfigMem.ConfigBits\[206\]
rlabel metal1 10212 15130 10212 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
rlabel metal1 16330 16694 16330 16694 0 Inst_RAM_IO_ConfigMem.ConfigBits\[208\]
rlabel metal1 17342 16626 17342 16626 0 Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
rlabel metal1 7728 15674 7728 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[210\]
rlabel metal1 8326 16218 8326 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
rlabel metal1 3450 20026 3450 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[212\]
rlabel metal2 4094 20604 4094 20604 0 Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
rlabel metal1 10488 17782 10488 17782 0 Inst_RAM_IO_ConfigMem.ConfigBits\[214\]
rlabel metal1 11040 17306 11040 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
rlabel metal1 12519 25330 12519 25330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[216\]
rlabel metal2 12466 26248 12466 26248 0 Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
rlabel metal2 3266 28458 3266 28458 0 Inst_RAM_IO_ConfigMem.ConfigBits\[218\]
rlabel metal1 3266 28118 3266 28118 0 Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
rlabel metal1 11040 36278 11040 36278 0 Inst_RAM_IO_ConfigMem.ConfigBits\[220\]
rlabel viali 11563 36142 11563 36142 0 Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
rlabel metal1 16468 28186 16468 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[222\]
rlabel metal1 17342 28594 17342 28594 0 Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
rlabel metal2 13478 28186 13478 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[224\]
rlabel metal1 14306 26894 14306 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
rlabel metal2 3542 24276 3542 24276 0 Inst_RAM_IO_ConfigMem.ConfigBits\[226\]
rlabel metal1 3312 23290 3312 23290 0 Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
rlabel metal1 10580 32946 10580 32946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[228\]
rlabel metal1 11132 32538 11132 32538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
rlabel metal1 17296 26894 17296 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[230\]
rlabel metal2 17894 27132 17894 27132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
rlabel metal2 11086 27132 11086 27132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[232\]
rlabel metal2 11914 27336 11914 27336 0 Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
rlabel metal2 4922 28186 4922 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[234\]
rlabel metal1 5566 26826 5566 26826 0 Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
rlabel metal1 10534 35190 10534 35190 0 Inst_RAM_IO_ConfigMem.ConfigBits\[236\]
rlabel metal2 11086 34714 11086 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
rlabel metal1 16284 30838 16284 30838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[238\]
rlabel metal1 17204 30770 17204 30770 0 Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
rlabel metal1 13248 23630 13248 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[240\]
rlabel metal2 13846 23868 13846 23868 0 Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
rlabel metal1 3588 25398 3588 25398 0 Inst_RAM_IO_ConfigMem.ConfigBits\[242\]
rlabel metal1 4416 25262 4416 25262 0 Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
rlabel metal2 12926 33184 12926 33184 0 Inst_RAM_IO_ConfigMem.ConfigBits\[244\]
rlabel metal1 13386 33422 13386 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
rlabel metal1 17526 24922 17526 24922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[246\]
rlabel metal1 18814 24582 18814 24582 0 Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
rlabel metal1 16698 18938 16698 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[248\]
rlabel metal1 17296 19482 17296 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
rlabel metal2 7682 19482 7682 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[250\]
rlabel metal1 7820 18938 7820 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
rlabel metal2 5842 20060 5842 20060 0 Inst_RAM_IO_ConfigMem.ConfigBits\[252\]
rlabel metal1 5888 19482 5888 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
rlabel metal2 15410 20774 15410 20774 0 Inst_RAM_IO_ConfigMem.ConfigBits\[254\]
rlabel metal1 16054 20978 16054 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
rlabel metal2 15686 24038 15686 24038 0 Inst_RAM_IO_ConfigMem.ConfigBits\[256\]
rlabel metal1 16607 24242 16607 24242 0 Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
rlabel metal1 7084 22406 7084 22406 0 Inst_RAM_IO_ConfigMem.ConfigBits\[258\]
rlabel metal1 7544 21862 7544 21862 0 Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
rlabel metal2 7590 26010 7590 26010 0 Inst_RAM_IO_ConfigMem.ConfigBits\[260\]
rlabel metal1 8050 25466 8050 25466 0 Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
rlabel metal1 14536 21658 14536 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[262\]
rlabel via1 15318 22073 15318 22073 0 Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
rlabel metal1 12926 16218 12926 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[264\]
rlabel metal1 13478 17306 13478 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
rlabel metal1 2645 33354 2645 33354 0 Inst_RAM_IO_ConfigMem.ConfigBits\[266\]
rlabel metal1 3404 33082 3404 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
rlabel metal2 12374 40154 12374 40154 0 Inst_RAM_IO_ConfigMem.ConfigBits\[268\]
rlabel metal2 13386 39780 13386 39780 0 Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
rlabel metal1 18032 17850 18032 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[270\]
rlabel metal2 18354 18428 18354 18428 0 Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
rlabel metal1 10994 10132 10994 10132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[272\]
rlabel metal1 12742 9690 12742 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
rlabel metal1 3358 35156 3358 35156 0 Inst_RAM_IO_ConfigMem.ConfigBits\[274\]
rlabel metal1 4462 34714 4462 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
rlabel metal2 9154 38250 9154 38250 0 Inst_RAM_IO_ConfigMem.ConfigBits\[276\]
rlabel metal1 9338 37944 9338 37944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
rlabel metal1 13754 8058 13754 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[278\]
rlabel metal1 14214 8568 14214 8568 0 Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
rlabel metal2 12558 12070 12558 12070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[280\]
rlabel metal1 12466 12201 12466 12201 0 Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
rlabel metal1 3082 36618 3082 36618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[282\]
rlabel metal1 3818 36856 3818 36856 0 Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
rlabel metal1 8464 36550 8464 36550 0 Inst_RAM_IO_ConfigMem.ConfigBits\[284\]
rlabel metal2 8602 35870 8602 35870 0 Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
rlabel metal2 13938 12070 13938 12070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[286\]
rlabel metal2 14674 12410 14674 12410 0 Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
rlabel metal2 11914 15130 11914 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[288\]
rlabel metal1 12190 14586 12190 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
rlabel metal2 4830 40052 4830 40052 0 Inst_RAM_IO_ConfigMem.ConfigBits\[290\]
rlabel metal1 4462 39406 4462 39406 0 Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
rlabel metal2 7958 40154 7958 40154 0 Inst_RAM_IO_ConfigMem.ConfigBits\[292\]
rlabel metal2 8418 39984 8418 39984 0 Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
rlabel metal1 13294 10506 13294 10506 0 Inst_RAM_IO_ConfigMem.ConfigBits\[294\]
rlabel metal1 14582 10234 14582 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
rlabel metal1 11040 8058 11040 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[296\]
rlabel metal1 12190 8058 12190 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
rlabel metal1 2990 37740 2990 37740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[298\]
rlabel metal1 3910 37944 3910 37944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
rlabel metal2 9614 40426 9614 40426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[300\]
rlabel metal1 10166 39610 10166 39610 0 Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
rlabel metal1 13524 6970 13524 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[302\]
rlabel metal1 14214 6426 14214 6426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
rlabel metal1 10856 2618 10856 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[304\]
rlabel metal2 10350 3502 10350 3502 0 Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
rlabel metal2 3358 31076 3358 31076 0 Inst_RAM_IO_ConfigMem.ConfigBits\[306\]
rlabel metal1 4968 30906 4968 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
rlabel metal2 5198 29852 5198 29852 0 Inst_RAM_IO_ConfigMem.ConfigBits\[308\]
rlabel metal1 5658 29274 5658 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
rlabel metal2 11086 22950 11086 22950 0 Inst_RAM_IO_ConfigMem.ConfigBits\[310\]
rlabel metal1 11592 23086 11592 23086 0 Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
rlabel metal2 6118 3162 6118 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[312\]
rlabel metal1 6900 2618 6900 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
rlabel metal1 6164 17034 6164 17034 0 Inst_RAM_IO_ConfigMem.ConfigBits\[314\]
rlabel metal2 6946 17238 6946 17238 0 Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
rlabel metal2 9108 31892 9108 31892 0 Inst_RAM_IO_ConfigMem.ConfigBits\[316\]
rlabel metal1 9522 30906 9522 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
rlabel metal2 12558 3740 12558 3740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[318\]
rlabel metal1 12834 3162 12834 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
rlabel metal2 12558 18666 12558 18666 0 Inst_RAM_IO_ConfigMem.ConfigBits\[320\]
rlabel metal1 12190 18326 12190 18326 0 Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
rlabel metal1 2714 38794 2714 38794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[322\]
rlabel metal2 2346 39576 2346 39576 0 Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
rlabel metal1 10626 41650 10626 41650 0 Inst_RAM_IO_ConfigMem.ConfigBits\[324\]
rlabel metal2 11086 40732 11086 40732 0 Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
rlabel metal1 13662 16660 13662 16660 0 Inst_RAM_IO_ConfigMem.ConfigBits\[326\]
rlabel metal1 15180 16218 15180 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
rlabel metal1 9200 27098 9200 27098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[48\]
rlabel metal1 10258 27506 10258 27506 0 Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
rlabel metal1 2300 34714 2300 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[50\]
rlabel metal2 2714 35836 2714 35836 0 Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
rlabel metal2 12558 38624 12558 38624 0 Inst_RAM_IO_ConfigMem.ConfigBits\[52\]
rlabel metal1 12880 37978 12880 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
rlabel metal1 14766 33048 14766 33048 0 Inst_RAM_IO_ConfigMem.ConfigBits\[54\]
rlabel metal2 15318 33796 15318 33796 0 Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
rlabel metal1 9989 23630 9989 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[56\]
rlabel metal2 9246 23494 9246 23494 0 Inst_RAM_IO_ConfigMem.ConfigBits\[57\]
rlabel metal2 2162 30634 2162 30634 0 Inst_RAM_IO_ConfigMem.ConfigBits\[58\]
rlabel metal2 2714 30022 2714 30022 0 Inst_RAM_IO_ConfigMem.ConfigBits\[59\]
rlabel metal1 1932 32334 1932 32334 0 Inst_RAM_IO_ConfigMem.ConfigBits\[60\]
rlabel metal1 2530 31994 2530 31994 0 Inst_RAM_IO_ConfigMem.ConfigBits\[61\]
rlabel metal1 7590 29784 7590 29784 0 Inst_RAM_IO_ConfigMem.ConfigBits\[62\]
rlabel metal1 8280 29274 8280 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[63\]
rlabel metal1 2392 21658 2392 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[64\]
rlabel metal1 2300 21998 2300 21998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[65\]
rlabel metal2 2622 23766 2622 23766 0 Inst_RAM_IO_ConfigMem.ConfigBits\[66\]
rlabel metal2 1978 24888 1978 24888 0 Inst_RAM_IO_ConfigMem.ConfigBits\[67\]
rlabel metal2 2530 27098 2530 27098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[68\]
rlabel metal1 2530 26554 2530 26554 0 Inst_RAM_IO_ConfigMem.ConfigBits\[69\]
rlabel metal2 8510 21284 8510 21284 0 Inst_RAM_IO_ConfigMem.ConfigBits\[70\]
rlabel metal1 9430 21114 9430 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[71\]
rlabel metal2 9706 25194 9706 25194 0 Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
rlabel metal1 10350 25806 10350 25806 0 Inst_RAM_IO_ConfigMem.ConfigBits\[73\]
rlabel metal1 10994 29138 10994 29138 0 Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
rlabel metal2 5750 36686 5750 36686 0 Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
rlabel metal2 6302 35700 6302 35700 0 Inst_RAM_IO_ConfigMem.ConfigBits\[76\]
rlabel metal1 7774 37230 7774 37230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
rlabel metal1 7452 34102 7452 34102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
rlabel metal2 8096 33490 8096 33490 0 Inst_RAM_IO_ConfigMem.ConfigBits\[79\]
rlabel metal1 9798 34442 9798 34442 0 Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
rlabel metal2 16238 31518 16238 31518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
rlabel metal1 16882 31858 16882 31858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[82\]
rlabel viali 16698 34600 16698 34600 0 Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
rlabel metal2 10994 20570 10994 20570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[84\]
rlabel metal1 10902 20026 10902 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
rlabel metal2 5566 33388 5566 33388 0 Inst_RAM_IO_ConfigMem.ConfigBits\[86\]
rlabel metal2 5382 33082 5382 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
rlabel metal2 12834 35428 12834 35428 0 Inst_RAM_IO_ConfigMem.ConfigBits\[88\]
rlabel metal1 12098 35768 12098 35768 0 Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
rlabel metal2 15134 32164 15134 32164 0 Inst_RAM_IO_ConfigMem.ConfigBits\[90\]
rlabel metal2 14490 33694 14490 33694 0 Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
rlabel metal1 11270 22202 11270 22202 0 Inst_RAM_IO_ConfigMem.ConfigBits\[92\]
rlabel metal2 12006 21794 12006 21794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[93\]
rlabel metal1 5842 27540 5842 27540 0 Inst_RAM_IO_ConfigMem.ConfigBits\[94\]
rlabel metal2 6762 27642 6762 27642 0 Inst_RAM_IO_ConfigMem.ConfigBits\[95\]
rlabel metal2 6854 31833 6854 31833 0 Inst_RAM_IO_ConfigMem.ConfigBits\[96\]
rlabel metal1 7268 30906 7268 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[97\]
rlabel metal2 14950 29546 14950 29546 0 Inst_RAM_IO_ConfigMem.ConfigBits\[98\]
rlabel metal1 14674 29240 14674 29240 0 Inst_RAM_IO_ConfigMem.ConfigBits\[99\]
rlabel metal1 12972 18122 12972 18122 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG0
rlabel metal1 4370 39270 4370 39270 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG1
rlabel metal1 12558 39882 12558 39882 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG2
rlabel metal1 18745 18190 18745 18190 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG3
rlabel metal1 16997 19890 16997 19890 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
rlabel metal1 6762 19482 6762 19482 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
rlabel metal1 5612 26214 5612 26214 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
rlabel metal2 16238 8449 16238 8449 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
rlabel metal2 2070 21267 2070 21267 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
rlabel metal1 5704 24242 5704 24242 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
rlabel metal1 2622 4658 2622 4658 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
rlabel metal1 14766 18734 14766 18734 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
rlabel metal1 12834 9928 12834 9928 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG0
rlabel metal1 3036 20366 3036 20366 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG1
rlabel metal3 9085 13668 9085 13668 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
rlabel metal1 16744 21386 16744 21386 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
rlabel metal2 8510 9146 8510 9146 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
rlabel metal1 4462 25194 4462 25194 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
rlabel metal2 12742 33558 12742 33558 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
rlabel via1 17779 21522 17779 21522 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
rlabel metal1 1012 34170 1012 34170 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG2
rlabel metal1 16836 32198 16836 32198 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG3
rlabel metal1 12834 12104 12834 12104 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
rlabel via1 2818 17646 2818 17646 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
rlabel metal1 1150 21998 1150 21998 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
rlabel metal2 16882 21114 16882 21114 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
rlabel metal1 13202 25806 13202 25806 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
rlabel metal1 5244 39270 5244 39270 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
rlabel metal3 1035 27132 1035 27132 0 Inst_RAM_IO_switch_matrix.N1BEG0
rlabel metal1 3450 35802 3450 35802 0 Inst_RAM_IO_switch_matrix.N1BEG1
rlabel metal2 13202 42636 13202 42636 0 Inst_RAM_IO_switch_matrix.N1BEG2
rlabel metal1 16054 33082 16054 33082 0 Inst_RAM_IO_switch_matrix.N1BEG3
rlabel metal1 1656 41446 1656 41446 0 Inst_RAM_IO_switch_matrix.N2BEG0
rlabel metal1 1150 43282 1150 43282 0 Inst_RAM_IO_switch_matrix.N2BEG1
rlabel metal1 3496 32470 3496 32470 0 Inst_RAM_IO_switch_matrix.N2BEG2
rlabel metal2 8694 41400 8694 41400 0 Inst_RAM_IO_switch_matrix.N2BEG3
rlabel metal3 3335 40052 3335 40052 0 Inst_RAM_IO_switch_matrix.N2BEG4
rlabel metal1 1150 36074 1150 36074 0 Inst_RAM_IO_switch_matrix.N2BEG5
rlabel metal1 1932 41650 1932 41650 0 Inst_RAM_IO_switch_matrix.N2BEG6
rlabel metal4 13892 30124 13892 30124 0 Inst_RAM_IO_switch_matrix.N2BEG7
rlabel metal4 1012 22712 1012 22712 0 Inst_RAM_IO_switch_matrix.N2BEGb0
rlabel metal2 3266 36550 3266 36550 0 Inst_RAM_IO_switch_matrix.N2BEGb1
rlabel metal4 2668 36380 2668 36380 0 Inst_RAM_IO_switch_matrix.N2BEGb2
rlabel metal1 2438 42194 2438 42194 0 Inst_RAM_IO_switch_matrix.N2BEGb3
rlabel metal4 828 22508 828 22508 0 Inst_RAM_IO_switch_matrix.N2BEGb4
rlabel metal2 1104 27676 1104 27676 0 Inst_RAM_IO_switch_matrix.N2BEGb5
rlabel metal1 4922 31994 4922 31994 0 Inst_RAM_IO_switch_matrix.N2BEGb6
rlabel metal4 644 22508 644 22508 0 Inst_RAM_IO_switch_matrix.N2BEGb7
rlabel metal2 10902 35337 10902 35337 0 Inst_RAM_IO_switch_matrix.N4BEG0
rlabel metal1 8188 37094 8188 37094 0 Inst_RAM_IO_switch_matrix.N4BEG1
rlabel metal2 9200 41684 9200 41684 0 Inst_RAM_IO_switch_matrix.N4BEG2
rlabel metal1 16192 34714 16192 34714 0 Inst_RAM_IO_switch_matrix.N4BEG3
rlabel metal2 782 16388 782 16388 0 Inst_RAM_IO_switch_matrix.S1BEG0
rlabel metal2 14030 32368 14030 32368 0 Inst_RAM_IO_switch_matrix.S1BEG1
rlabel metal1 13432 2618 13432 2618 0 Inst_RAM_IO_switch_matrix.S1BEG2
rlabel metal1 15548 2618 15548 2618 0 Inst_RAM_IO_switch_matrix.S1BEG3
rlabel metal2 13846 1887 13846 1887 0 Inst_RAM_IO_switch_matrix.S2BEG0
rlabel metal2 598 16252 598 16252 0 Inst_RAM_IO_switch_matrix.S2BEG1
rlabel metal1 13616 1938 13616 1938 0 Inst_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 16100 2414 16100 2414 0 Inst_RAM_IO_switch_matrix.S2BEG3
rlabel metal1 15226 1870 15226 1870 0 Inst_RAM_IO_switch_matrix.S2BEG4
rlabel metal3 14375 2380 14375 2380 0 Inst_RAM_IO_switch_matrix.S2BEG5
rlabel metal4 10948 17068 10948 17068 0 Inst_RAM_IO_switch_matrix.S2BEG6
rlabel via3 15571 18020 15571 18020 0 Inst_RAM_IO_switch_matrix.S2BEG7
rlabel metal2 13524 1394 13524 1394 0 Inst_RAM_IO_switch_matrix.S2BEGb0
rlabel metal3 11615 4012 11615 4012 0 Inst_RAM_IO_switch_matrix.S2BEGb1
rlabel via3 11845 4012 11845 4012 0 Inst_RAM_IO_switch_matrix.S2BEGb2
rlabel metal1 9108 1326 9108 1326 0 Inst_RAM_IO_switch_matrix.S2BEGb3
rlabel metal2 11868 2788 11868 2788 0 Inst_RAM_IO_switch_matrix.S2BEGb4
rlabel via3 12581 16660 12581 16660 0 Inst_RAM_IO_switch_matrix.S2BEGb5
rlabel metal3 13961 2652 13961 2652 0 Inst_RAM_IO_switch_matrix.S2BEGb6
rlabel metal2 13386 1873 13386 1873 0 Inst_RAM_IO_switch_matrix.S2BEGb7
rlabel metal3 17641 17204 17641 17204 0 Inst_RAM_IO_switch_matrix.S4BEG0
rlabel metal2 19458 22882 19458 22882 0 Inst_RAM_IO_switch_matrix.S4BEG1
rlabel metal1 17480 20230 17480 20230 0 Inst_RAM_IO_switch_matrix.S4BEG2
rlabel metal2 20240 17068 20240 17068 0 Inst_RAM_IO_switch_matrix.S4BEG3
rlabel metal1 2346 3400 2346 3400 0 Inst_RAM_IO_switch_matrix.W1BEG0
rlabel metal1 5750 5746 5750 5746 0 Inst_RAM_IO_switch_matrix.W1BEG1
rlabel metal1 8464 11050 8464 11050 0 Inst_RAM_IO_switch_matrix.W1BEG2
rlabel via2 8050 4539 8050 4539 0 Inst_RAM_IO_switch_matrix.W1BEG3
rlabel metal1 4278 6698 4278 6698 0 Inst_RAM_IO_switch_matrix.W2BEG0
rlabel metal1 6026 5338 6026 5338 0 Inst_RAM_IO_switch_matrix.W2BEG1
rlabel metal1 5612 6290 5612 6290 0 Inst_RAM_IO_switch_matrix.W2BEG2
rlabel metal1 8372 6290 8372 6290 0 Inst_RAM_IO_switch_matrix.W2BEG3
rlabel metal1 2346 4012 2346 4012 0 Inst_RAM_IO_switch_matrix.W2BEG4
rlabel metal2 4278 10064 4278 10064 0 Inst_RAM_IO_switch_matrix.W2BEG5
rlabel metal1 4416 4114 4416 4114 0 Inst_RAM_IO_switch_matrix.W2BEG6
rlabel metal1 2507 3026 2507 3026 0 Inst_RAM_IO_switch_matrix.W2BEG7
rlabel metal1 2254 6732 2254 6732 0 Inst_RAM_IO_switch_matrix.W2BEGb0
rlabel metal1 2208 7378 2208 7378 0 Inst_RAM_IO_switch_matrix.W2BEGb1
rlabel metal1 3496 17238 3496 17238 0 Inst_RAM_IO_switch_matrix.W2BEGb2
rlabel metal1 7728 8058 7728 8058 0 Inst_RAM_IO_switch_matrix.W2BEGb3
rlabel metal1 14490 5032 14490 5032 0 Inst_RAM_IO_switch_matrix.W2BEGb4
rlabel metal1 3588 14246 3588 14246 0 Inst_RAM_IO_switch_matrix.W2BEGb5
rlabel metal1 1702 4522 1702 4522 0 Inst_RAM_IO_switch_matrix.W2BEGb6
rlabel metal1 5014 3604 5014 3604 0 Inst_RAM_IO_switch_matrix.W2BEGb7
rlabel metal2 7406 14127 7406 14127 0 Inst_RAM_IO_switch_matrix.W6BEG0
rlabel metal1 1518 39032 1518 39032 0 Inst_RAM_IO_switch_matrix.W6BEG1
rlabel metal1 3266 19380 3266 19380 0 Inst_RAM_IO_switch_matrix.W6BEG10
rlabel metal1 11684 17646 11684 17646 0 Inst_RAM_IO_switch_matrix.W6BEG11
rlabel metal1 1610 36856 1610 36856 0 Inst_RAM_IO_switch_matrix.W6BEG2
rlabel metal2 7866 14467 7866 14467 0 Inst_RAM_IO_switch_matrix.W6BEG3
rlabel metal2 15318 14535 15318 14535 0 Inst_RAM_IO_switch_matrix.W6BEG4
rlabel metal2 1886 13464 1886 13464 0 Inst_RAM_IO_switch_matrix.W6BEG5
rlabel metal2 5382 16354 5382 16354 0 Inst_RAM_IO_switch_matrix.W6BEG6
rlabel metal1 10718 15674 10718 15674 0 Inst_RAM_IO_switch_matrix.W6BEG7
rlabel metal1 17664 16558 17664 16558 0 Inst_RAM_IO_switch_matrix.W6BEG8
rlabel metal1 6302 16762 6302 16762 0 Inst_RAM_IO_switch_matrix.W6BEG9
rlabel metal2 18446 7888 18446 7888 0 Inst_RAM_IO_switch_matrix.WW4BEG0
rlabel metal1 4646 13940 4646 13940 0 Inst_RAM_IO_switch_matrix.WW4BEG1
rlabel metal1 1610 17238 1610 17238 0 Inst_RAM_IO_switch_matrix.WW4BEG10
rlabel metal1 9706 12954 9706 12954 0 Inst_RAM_IO_switch_matrix.WW4BEG11
rlabel metal1 15962 7718 15962 7718 0 Inst_RAM_IO_switch_matrix.WW4BEG12
rlabel metal1 4002 14416 4002 14416 0 Inst_RAM_IO_switch_matrix.WW4BEG13
rlabel metal1 4232 7514 4232 7514 0 Inst_RAM_IO_switch_matrix.WW4BEG14
rlabel metal2 11270 10166 11270 10166 0 Inst_RAM_IO_switch_matrix.WW4BEG15
rlabel metal2 2162 10438 2162 10438 0 Inst_RAM_IO_switch_matrix.WW4BEG2
rlabel via2 1610 9571 1610 9571 0 Inst_RAM_IO_switch_matrix.WW4BEG3
rlabel via2 17066 11237 17066 11237 0 Inst_RAM_IO_switch_matrix.WW4BEG4
rlabel metal1 5658 11186 5658 11186 0 Inst_RAM_IO_switch_matrix.WW4BEG5
rlabel metal1 4692 12614 4692 12614 0 Inst_RAM_IO_switch_matrix.WW4BEG6
rlabel metal1 3818 13430 3818 13430 0 Inst_RAM_IO_switch_matrix.WW4BEG7
rlabel metal2 18262 11917 18262 11917 0 Inst_RAM_IO_switch_matrix.WW4BEG8
rlabel metal2 7590 10472 7590 10472 0 Inst_RAM_IO_switch_matrix.WW4BEG9
rlabel metal1 10810 26010 10810 26010 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0
rlabel metal1 11040 26554 11040 26554 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1
rlabel metal1 11086 28492 11086 28492 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 11546 28560 11546 28560 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 11178 28866 11178 28866 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_
rlabel metal1 11178 29070 11178 29070 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
rlabel metal1 6762 35802 6762 35802 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0
rlabel metal1 7176 36210 7176 36210 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1
rlabel metal1 6992 36346 6992 36346 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 7222 36856 7222 36856 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 7176 36754 7176 36754 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_
rlabel metal1 8326 37298 8326 37298 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
rlabel metal1 9338 33456 9338 33456 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0
rlabel metal1 8878 33490 8878 33490 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1
rlabel metal1 9384 33626 9384 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 8970 33626 8970 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 9292 34442 9292 34442 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_
rlabel metal1 8924 34510 8924 34510 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
rlabel metal1 17296 31858 17296 31858 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0
rlabel metal1 17480 29818 17480 29818 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1
rlabel metal1 16974 33592 16974 33592 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 17434 34170 17434 34170 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 16974 34442 16974 34442 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_
rlabel metal1 17204 34510 17204 34510 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
rlabel metal1 14950 27438 14950 27438 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0
rlabel metal1 15226 25874 15226 25874 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1
rlabel metal1 15594 25908 15594 25908 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 16054 25840 16054 25840 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 15686 26180 15686 26180 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_
rlabel metal2 16054 26146 16054 26146 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
rlabel metal1 7129 24174 7129 24174 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0
rlabel metal1 7958 24208 7958 24208 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1
rlabel metal1 7498 24140 7498 24140 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 8510 23732 8510 23732 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 7820 23086 7820 23086 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_
rlabel metal1 8464 23086 8464 23086 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
rlabel metal1 12558 30702 12558 30702 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0
rlabel metal1 13018 30634 13018 30634 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1
rlabel metal2 12558 31348 12558 31348 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 13248 30906 13248 30906 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 13524 31790 13524 31790 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_
rlabel metal1 14950 30736 14950 30736 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
rlabel metal1 18492 21998 18492 21998 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0
rlabel metal1 18676 21522 18676 21522 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1
rlabel metal1 18446 21862 18446 21862 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 19458 20944 19458 20944 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 18677 20910 18677 20910 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_
rlabel metal1 19228 20842 19228 20842 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
rlabel metal2 230 44193 230 44193 0 N1BEG[0]
rlabel metal2 506 43428 506 43428 0 N1BEG[1]
rlabel metal2 782 43156 782 43156 0 N1BEG[2]
rlabel metal2 1058 43309 1058 43309 0 N1BEG[3]
rlabel metal2 230 1214 230 1214 0 N1END[0]
rlabel metal2 506 1248 506 1248 0 N1END[1]
rlabel metal2 881 68 881 68 0 N1END[2]
rlabel metal1 1288 3026 1288 3026 0 N1END[3]
rlabel metal2 1334 43649 1334 43649 0 N2BEG[0]
rlabel metal2 1610 43156 1610 43156 0 N2BEG[1]
rlabel metal2 1886 43972 1886 43972 0 N2BEG[2]
rlabel metal2 2162 44057 2162 44057 0 N2BEG[3]
rlabel metal1 2576 41242 2576 41242 0 N2BEG[4]
rlabel metal2 2714 43649 2714 43649 0 N2BEG[5]
rlabel metal1 2898 43418 2898 43418 0 N2BEG[6]
rlabel metal2 3266 44057 3266 44057 0 N2BEG[7]
rlabel metal1 2990 42092 2990 42092 0 N2BEGb[0]
rlabel metal1 4186 42126 4186 42126 0 N2BEGb[1]
rlabel metal2 4094 44057 4094 44057 0 N2BEGb[2]
rlabel metal2 4370 43972 4370 43972 0 N2BEGb[3]
rlabel metal1 4692 42534 4692 42534 0 N2BEGb[4]
rlabel metal2 4922 43632 4922 43632 0 N2BEGb[5]
rlabel metal1 4968 42330 4968 42330 0 N2BEGb[6]
rlabel metal2 5474 44193 5474 44193 0 N2BEGb[7]
rlabel metal2 3489 68 3489 68 0 N2END[0]
rlabel metal2 3818 636 3818 636 0 N2END[1]
rlabel metal2 4094 755 4094 755 0 N2END[2]
rlabel metal2 4469 68 4469 68 0 N2END[3]
rlabel metal2 4646 1044 4646 1044 0 N2END[4]
rlabel metal2 4922 551 4922 551 0 N2END[5]
rlabel metal2 5251 68 5251 68 0 N2END[6]
rlabel metal2 5474 1180 5474 1180 0 N2END[7]
rlabel metal2 1334 1010 1334 1010 0 N2MID[0]
rlabel metal2 1663 68 1663 68 0 N2MID[1]
rlabel metal2 1985 68 1985 68 0 N2MID[2]
rlabel metal2 2261 68 2261 68 0 N2MID[3]
rlabel metal2 2438 398 2438 398 0 N2MID[4]
rlabel metal2 2714 1520 2714 1520 0 N2MID[5]
rlabel metal2 3043 68 3043 68 0 N2MID[6]
rlabel metal2 3266 1248 3266 1248 0 N2MID[7]
rlabel metal2 5750 43530 5750 43530 0 N4BEG[0]
rlabel metal1 8418 43418 8418 43418 0 N4BEG[10]
rlabel metal1 8740 42738 8740 42738 0 N4BEG[11]
rlabel metal1 8878 43418 8878 43418 0 N4BEG[12]
rlabel metal2 9338 43632 9338 43632 0 N4BEG[13]
rlabel metal1 9430 43418 9430 43418 0 N4BEG[14]
rlabel metal1 9844 43418 9844 43418 0 N4BEG[15]
rlabel metal2 6026 44057 6026 44057 0 N4BEG[1]
rlabel metal1 6210 43418 6210 43418 0 N4BEG[2]
rlabel metal2 6578 43921 6578 43921 0 N4BEG[3]
rlabel metal2 6854 44193 6854 44193 0 N4BEG[4]
rlabel metal2 7130 44193 7130 44193 0 N4BEG[5]
rlabel metal1 7728 42534 7728 42534 0 N4BEG[6]
rlabel metal1 7544 43418 7544 43418 0 N4BEG[7]
rlabel metal1 7866 43418 7866 43418 0 N4BEG[8]
rlabel metal2 8234 43428 8234 43428 0 N4BEG[9]
rlabel metal4 1196 22236 1196 22236 0 N4BEG_outbuf_0.A
rlabel metal2 4554 41786 4554 41786 0 N4BEG_outbuf_0.X
rlabel metal1 1656 2278 1656 2278 0 N4BEG_outbuf_1.A
rlabel metal1 5934 41616 5934 41616 0 N4BEG_outbuf_1.X
rlabel metal3 20355 13532 20355 13532 0 N4BEG_outbuf_10.A
rlabel metal1 9016 41582 9016 41582 0 N4BEG_outbuf_10.X
rlabel metal3 20447 13668 20447 13668 0 N4BEG_outbuf_11.A
rlabel metal1 10166 42160 10166 42160 0 N4BEG_outbuf_11.X
rlabel metal2 6210 2227 6210 2227 0 N4BEG_outbuf_2.A
rlabel metal1 5106 41548 5106 41548 0 N4BEG_outbuf_2.X
rlabel metal2 5842 2125 5842 2125 0 N4BEG_outbuf_3.A
rlabel metal1 5750 41582 5750 41582 0 N4BEG_outbuf_3.X
rlabel metal1 6808 2074 6808 2074 0 N4BEG_outbuf_4.A
rlabel metal1 6164 42330 6164 42330 0 N4BEG_outbuf_4.X
rlabel metal4 19780 24140 19780 24140 0 N4BEG_outbuf_5.A
rlabel metal1 7406 41616 7406 41616 0 N4BEG_outbuf_5.X
rlabel metal2 14628 16560 14628 16560 0 N4BEG_outbuf_6.A
rlabel metal1 7774 41616 7774 41616 0 N4BEG_outbuf_6.X
rlabel via3 7613 20740 7613 20740 0 N4BEG_outbuf_7.A
rlabel metal1 7958 41582 7958 41582 0 N4BEG_outbuf_7.X
rlabel metal2 13662 23324 13662 23324 0 N4BEG_outbuf_8.A
rlabel metal1 8326 41616 8326 41616 0 N4BEG_outbuf_8.X
rlabel metal1 8004 1938 8004 1938 0 N4BEG_outbuf_9.A
rlabel metal2 7958 41253 7958 41253 0 N4BEG_outbuf_9.X
rlabel metal2 5750 364 5750 364 0 N4END[0]
rlabel metal2 8510 1214 8510 1214 0 N4END[10]
rlabel metal2 8786 1248 8786 1248 0 N4END[11]
rlabel metal2 9115 68 9115 68 0 N4END[12]
rlabel metal2 9338 806 9338 806 0 N4END[13]
rlabel metal1 9062 2958 9062 2958 0 N4END[14]
rlabel metal2 9890 364 9890 364 0 N4END[15]
rlabel metal2 6026 551 6026 551 0 N4END[1]
rlabel metal2 6302 636 6302 636 0 N4END[2]
rlabel metal2 6578 670 6578 670 0 N4END[3]
rlabel metal2 6854 483 6854 483 0 N4END[4]
rlabel metal2 7130 483 7130 483 0 N4END[5]
rlabel metal2 7406 1231 7406 1231 0 N4END[6]
rlabel metal2 7682 1248 7682 1248 0 N4END[7]
rlabel metal2 7905 68 7905 68 0 N4END[8]
rlabel metal2 8181 68 8181 68 0 N4END[9]
rlabel metal3 24836 7140 24836 7140 0 RAM2FAB_D0_I0
rlabel metal2 21574 7293 21574 7293 0 RAM2FAB_D0_I1
rlabel metal3 25204 8228 25204 8228 0 RAM2FAB_D0_I2
rlabel metal3 25503 8772 25503 8772 0 RAM2FAB_D0_I3
rlabel metal2 20746 5389 20746 5389 0 RAM2FAB_D1_I0
rlabel metal3 25503 5508 25503 5508 0 RAM2FAB_D1_I1
rlabel metal2 20286 6239 20286 6239 0 RAM2FAB_D1_I2
rlabel metal2 20746 6528 20746 6528 0 RAM2FAB_D1_I3
rlabel metal2 20746 2975 20746 2975 0 RAM2FAB_D2_I0
rlabel metal2 20654 3332 20654 3332 0 RAM2FAB_D2_I1
rlabel metal2 21850 4301 21850 4301 0 RAM2FAB_D2_I2
rlabel metal3 25503 4420 25503 4420 0 RAM2FAB_D2_I3
rlabel metal1 19412 986 19412 986 0 RAM2FAB_D3_I0
rlabel metal3 25710 1156 25710 1156 0 RAM2FAB_D3_I1
rlabel metal2 20700 1836 20700 1836 0 RAM2FAB_D3_I2
rlabel metal1 19366 2550 19366 2550 0 RAM2FAB_D3_I3
rlabel metal2 10166 347 10166 347 0 S1BEG[0]
rlabel metal2 10495 68 10495 68 0 S1BEG[1]
rlabel metal2 10718 534 10718 534 0 S1BEG[2]
rlabel metal2 10994 908 10994 908 0 S1BEG[3]
rlabel metal2 10166 43904 10166 43904 0 S1END[0]
rlabel metal2 10442 43904 10442 43904 0 S1END[1]
rlabel metal2 10718 43904 10718 43904 0 S1END[2]
rlabel metal2 10994 43904 10994 43904 0 S1END[3]
rlabel metal2 13478 636 13478 636 0 S2BEG[0]
rlabel metal2 13754 738 13754 738 0 S2BEG[1]
rlabel metal2 14030 636 14030 636 0 S2BEG[2]
rlabel metal2 14306 908 14306 908 0 S2BEG[3]
rlabel metal2 14681 68 14681 68 0 S2BEG[4]
rlabel metal2 14858 347 14858 347 0 S2BEG[5]
rlabel metal2 15134 772 15134 772 0 S2BEG[6]
rlabel metal2 15410 942 15410 942 0 S2BEG[7]
rlabel metal2 11270 738 11270 738 0 S2BEGb[0]
rlabel metal2 11546 500 11546 500 0 S2BEGb[1]
rlabel metal2 11822 908 11822 908 0 S2BEGb[2]
rlabel metal2 12098 466 12098 466 0 S2BEGb[3]
rlabel metal2 12374 738 12374 738 0 S2BEGb[4]
rlabel metal2 12650 908 12650 908 0 S2BEGb[5]
rlabel metal2 12926 364 12926 364 0 S2BEGb[6]
rlabel metal2 13202 636 13202 636 0 S2BEGb[7]
rlabel metal2 11270 43904 11270 43904 0 S2END[0]
rlabel metal2 11546 44057 11546 44057 0 S2END[1]
rlabel metal2 11822 44329 11822 44329 0 S2END[2]
rlabel metal2 12098 43904 12098 43904 0 S2END[3]
rlabel metal2 12374 43938 12374 43938 0 S2END[4]
rlabel metal2 12650 43938 12650 43938 0 S2END[5]
rlabel metal2 12926 44125 12926 44125 0 S2END[6]
rlabel metal2 13202 44193 13202 44193 0 S2END[7]
rlabel metal2 13478 43904 13478 43904 0 S2MID[0]
rlabel metal2 13754 43632 13754 43632 0 S2MID[1]
rlabel metal2 14030 44057 14030 44057 0 S2MID[2]
rlabel metal2 14306 44057 14306 44057 0 S2MID[3]
rlabel metal2 14582 43938 14582 43938 0 S2MID[4]
rlabel metal2 14858 43938 14858 43938 0 S2MID[5]
rlabel metal2 15134 43632 15134 43632 0 S2MID[6]
rlabel metal2 15410 43904 15410 43904 0 S2MID[7]
rlabel metal2 15686 908 15686 908 0 S4BEG[0]
rlabel metal2 18446 1180 18446 1180 0 S4BEG[10]
rlabel metal2 18722 483 18722 483 0 S4BEG[11]
rlabel metal2 19097 68 19097 68 0 S4BEG[12]
rlabel metal1 19182 3366 19182 3366 0 S4BEG[13]
rlabel metal2 19649 68 19649 68 0 S4BEG[14]
rlabel metal2 19925 68 19925 68 0 S4BEG[15]
rlabel metal2 15962 347 15962 347 0 S4BEG[1]
rlabel metal2 16337 68 16337 68 0 S4BEG[2]
rlabel metal2 16514 143 16514 143 0 S4BEG[3]
rlabel metal2 16843 68 16843 68 0 S4BEG[4]
rlabel metal2 17066 619 17066 619 0 S4BEG[5]
rlabel metal2 17395 68 17395 68 0 S4BEG[6]
rlabel metal2 17618 908 17618 908 0 S4BEG[7]
rlabel metal2 17894 738 17894 738 0 S4BEG[8]
rlabel metal2 18223 68 18223 68 0 S4BEG[9]
rlabel metal1 16560 42194 16560 42194 0 S4BEG_outbuf_0.A
rlabel metal2 16422 20026 16422 20026 0 S4BEG_outbuf_0.X
rlabel metal1 16790 42296 16790 42296 0 S4BEG_outbuf_1.A
rlabel via2 17710 2397 17710 2397 0 S4BEG_outbuf_1.X
rlabel metal1 19228 40494 19228 40494 0 S4BEG_outbuf_10.A
rlabel metal3 18929 33116 18929 33116 0 S4BEG_outbuf_10.X
rlabel metal1 19458 40086 19458 40086 0 S4BEG_outbuf_11.A
rlabel metal2 19274 12580 19274 12580 0 S4BEG_outbuf_11.X
rlabel metal1 17250 42262 17250 42262 0 S4BEG_outbuf_2.A
rlabel metal1 17526 3026 17526 3026 0 S4BEG_outbuf_2.X
rlabel metal1 17664 42262 17664 42262 0 S4BEG_outbuf_3.A
rlabel metal3 17319 3876 17319 3876 0 S4BEG_outbuf_3.X
rlabel metal1 17986 42262 17986 42262 0 S4BEG_outbuf_4.A
rlabel metal1 17572 1870 17572 1870 0 S4BEG_outbuf_4.X
rlabel metal1 18308 42262 18308 42262 0 S4BEG_outbuf_5.A
rlabel metal3 21091 1292 21091 1292 0 S4BEG_outbuf_5.X
rlabel metal2 18630 42398 18630 42398 0 S4BEG_outbuf_6.A
rlabel metal2 18492 33116 18492 33116 0 S4BEG_outbuf_6.X
rlabel metal1 18998 42296 18998 42296 0 S4BEG_outbuf_7.A
rlabel via3 17733 3876 17733 3876 0 S4BEG_outbuf_7.X
rlabel metal1 18400 41582 18400 41582 0 S4BEG_outbuf_8.A
rlabel via3 18515 3876 18515 3876 0 S4BEG_outbuf_8.X
rlabel metal1 19458 42262 19458 42262 0 S4BEG_outbuf_9.A
rlabel metal3 19251 1292 19251 1292 0 S4BEG_outbuf_9.X
rlabel metal2 15686 43904 15686 43904 0 S4END[0]
rlabel metal2 18446 44125 18446 44125 0 S4END[10]
rlabel metal2 18722 44465 18722 44465 0 S4END[11]
rlabel metal2 19366 42126 19366 42126 0 S4END[12]
rlabel metal1 20102 40494 20102 40494 0 S4END[13]
rlabel metal2 19734 41253 19734 41253 0 S4END[14]
rlabel metal2 19826 43037 19826 43037 0 S4END[15]
rlabel metal2 15962 43938 15962 43938 0 S4END[1]
rlabel metal2 16238 43938 16238 43938 0 S4END[2]
rlabel metal2 16514 43649 16514 43649 0 S4END[3]
rlabel metal2 16790 43938 16790 43938 0 S4END[4]
rlabel metal2 17066 43972 17066 43972 0 S4END[5]
rlabel metal2 17342 43870 17342 43870 0 S4END[6]
rlabel metal2 17618 43921 17618 43921 0 S4END[7]
rlabel metal2 17894 43989 17894 43989 0 S4END[8]
rlabel metal2 18170 44176 18170 44176 0 S4END[9]
rlabel metal1 20746 17782 20746 17782 0 UserCLK
rlabel via1 20746 41803 20746 41803 0 UserCLKo
rlabel metal3 1142 4964 1142 4964 0 W1BEG[0]
rlabel metal2 2898 5389 2898 5389 0 W1BEG[1]
rlabel metal3 567 5508 567 5508 0 W1BEG[2]
rlabel metal3 728 5780 728 5780 0 W1BEG[3]
rlabel metal3 866 6052 866 6052 0 W2BEG[0]
rlabel metal3 728 6324 728 6324 0 W2BEG[1]
rlabel metal3 590 6596 590 6596 0 W2BEG[2]
rlabel metal3 682 6868 682 6868 0 W2BEG[3]
rlabel metal3 1142 7140 1142 7140 0 W2BEG[4]
rlabel metal3 958 7412 958 7412 0 W2BEG[5]
rlabel metal3 774 7684 774 7684 0 W2BEG[6]
rlabel metal2 3358 8143 3358 8143 0 W2BEG[7]
rlabel metal3 866 8228 866 8228 0 W2BEGb[0]
rlabel metal3 728 8500 728 8500 0 W2BEGb[1]
rlabel metal3 958 8772 958 8772 0 W2BEGb[2]
rlabel metal1 1978 8602 1978 8602 0 W2BEGb[3]
rlabel metal3 1234 9316 1234 9316 0 W2BEGb[4]
rlabel metal3 544 9588 544 9588 0 W2BEGb[5]
rlabel metal3 774 9860 774 9860 0 W2BEGb[6]
rlabel metal3 544 10132 544 10132 0 W2BEGb[7]
rlabel metal1 2438 13192 2438 13192 0 W6BEG[0]
rlabel metal3 958 17476 958 17476 0 W6BEG[10]
rlabel metal3 475 17748 475 17748 0 W6BEG[11]
rlabel metal3 1234 15028 1234 15028 0 W6BEG[1]
rlabel metal3 774 15300 774 15300 0 W6BEG[2]
rlabel metal2 3082 15351 3082 15351 0 W6BEG[3]
rlabel metal3 3404 15708 3404 15708 0 W6BEG[4]
rlabel metal2 3082 16269 3082 16269 0 W6BEG[5]
rlabel via2 4002 16405 4002 16405 0 W6BEG[6]
rlabel metal2 2898 16167 2898 16167 0 W6BEG[7]
rlabel metal3 567 16932 567 16932 0 W6BEG[8]
rlabel metal3 820 17204 820 17204 0 W6BEG[9]
rlabel metal3 912 10404 912 10404 0 WW4BEG[0]
rlabel metal3 682 13124 682 13124 0 WW4BEG[10]
rlabel metal2 4186 13396 4186 13396 0 WW4BEG[11]
rlabel metal3 728 13668 728 13668 0 WW4BEG[12]
rlabel metal3 912 13940 912 13940 0 WW4BEG[13]
rlabel metal3 1027 14212 1027 14212 0 WW4BEG[14]
rlabel metal3 1740 14484 1740 14484 0 WW4BEG[15]
rlabel metal2 4002 10829 4002 10829 0 WW4BEG[1]
rlabel metal3 1188 10948 1188 10948 0 WW4BEG[2]
rlabel metal2 3910 11271 3910 11271 0 WW4BEG[3]
rlabel metal3 1050 11492 1050 11492 0 WW4BEG[4]
rlabel metal2 3266 11509 3266 11509 0 WW4BEG[5]
rlabel metal3 774 12036 774 12036 0 WW4BEG[6]
rlabel metal2 3818 12189 3818 12189 0 WW4BEG[7]
rlabel metal3 866 12580 866 12580 0 WW4BEG[8]
rlabel metal3 1142 12852 1142 12852 0 WW4BEG[9]
rlabel metal1 23276 26554 23276 26554 0 data_inbuf_0.X
rlabel metal1 23782 27642 23782 27642 0 data_inbuf_1.X
rlabel metal1 21965 32266 21965 32266 0 data_inbuf_10.X
rlabel metal1 23598 32470 23598 32470 0 data_inbuf_11.X
rlabel metal1 23046 32946 23046 32946 0 data_inbuf_12.X
rlabel metal1 23552 33966 23552 33966 0 data_inbuf_13.X
rlabel metal1 22770 34646 22770 34646 0 data_inbuf_14.X
rlabel metal2 19458 34850 19458 34850 0 data_inbuf_15.X
rlabel metal1 21896 35666 21896 35666 0 data_inbuf_16.X
rlabel metal1 23322 35598 23322 35598 0 data_inbuf_17.X
rlabel metal1 21850 36176 21850 36176 0 data_inbuf_18.X
rlabel metal1 19826 36720 19826 36720 0 data_inbuf_19.X
rlabel metal1 23690 28016 23690 28016 0 data_inbuf_2.X
rlabel metal1 21114 36720 21114 36720 0 data_inbuf_20.X
rlabel metal1 23138 37128 23138 37128 0 data_inbuf_21.X
rlabel metal1 23138 37434 23138 37434 0 data_inbuf_22.X
rlabel metal2 23230 37842 23230 37842 0 data_inbuf_23.X
rlabel metal1 20286 38522 20286 38522 0 data_inbuf_24.X
rlabel metal1 23046 39372 23046 39372 0 data_inbuf_25.X
rlabel metal1 21206 40018 21206 40018 0 data_inbuf_26.X
rlabel metal1 20470 40528 20470 40528 0 data_inbuf_27.X
rlabel metal1 20194 41650 20194 41650 0 data_inbuf_28.X
rlabel metal2 21942 39984 21942 39984 0 data_inbuf_29.X
rlabel metal1 23690 28560 23690 28560 0 data_inbuf_3.X
rlabel metal1 23184 39270 23184 39270 0 data_inbuf_30.X
rlabel metal1 20654 40018 20654 40018 0 data_inbuf_31.X
rlabel metal1 23874 29172 23874 29172 0 data_inbuf_4.X
rlabel metal1 23736 29614 23736 29614 0 data_inbuf_5.X
rlabel metal1 23966 30192 23966 30192 0 data_inbuf_6.X
rlabel metal1 23690 30804 23690 30804 0 data_inbuf_7.X
rlabel metal1 23138 31280 23138 31280 0 data_inbuf_8.X
rlabel metal1 21390 31824 21390 31824 0 data_inbuf_9.X
rlabel metal1 24150 26928 24150 26928 0 data_outbuf_0.X
rlabel metal1 23506 26996 23506 26996 0 data_outbuf_1.X
rlabel metal1 23138 32402 23138 32402 0 data_outbuf_10.X
rlabel metal1 23874 32368 23874 32368 0 data_outbuf_11.X
rlabel metal1 23046 32742 23046 32742 0 data_outbuf_12.X
rlabel metal1 23230 33966 23230 33966 0 data_outbuf_13.X
rlabel metal1 23230 34476 23230 34476 0 data_outbuf_14.X
rlabel metal1 20746 35054 20746 35054 0 data_outbuf_15.X
rlabel metal1 22310 35734 22310 35734 0 data_outbuf_16.X
rlabel metal1 23092 35802 23092 35802 0 data_outbuf_17.X
rlabel metal1 21873 36006 21873 36006 0 data_outbuf_18.X
rlabel metal1 20792 36754 20792 36754 0 data_outbuf_19.X
rlabel metal1 23459 28050 23459 28050 0 data_outbuf_2.X
rlabel metal1 21390 36890 21390 36890 0 data_outbuf_20.X
rlabel metal1 23782 39066 23782 39066 0 data_outbuf_21.X
rlabel metal1 23644 38522 23644 38522 0 data_outbuf_22.X
rlabel metal1 23414 38454 23414 38454 0 data_outbuf_23.X
rlabel metal1 20470 39032 20470 39032 0 data_outbuf_24.X
rlabel metal1 22172 39270 22172 39270 0 data_outbuf_25.X
rlabel metal1 20286 40052 20286 40052 0 data_outbuf_26.X
rlabel metal2 20286 40477 20286 40477 0 data_outbuf_27.X
rlabel metal1 21298 41582 21298 41582 0 data_outbuf_28.X
rlabel metal2 22954 40086 22954 40086 0 data_outbuf_29.X
rlabel metal1 23506 28526 23506 28526 0 data_outbuf_3.X
rlabel metal1 23414 40086 23414 40086 0 data_outbuf_30.X
rlabel metal1 22586 39984 22586 39984 0 data_outbuf_31.X
rlabel metal1 23598 29070 23598 29070 0 data_outbuf_4.X
rlabel metal1 23556 29614 23556 29614 0 data_outbuf_5.X
rlabel metal1 23828 30362 23828 30362 0 data_outbuf_6.X
rlabel metal1 23046 30736 23046 30736 0 data_outbuf_7.X
rlabel metal1 23598 31314 23598 31314 0 data_outbuf_8.X
rlabel metal1 21850 31858 21850 31858 0 data_outbuf_9.X
rlabel metal1 12282 17612 12282 17612 0 net1
rlabel metal1 2070 31926 2070 31926 0 net10
rlabel via1 21850 17085 21850 17085 0 net100
rlabel metal1 2024 2550 2024 2550 0 net101
rlabel metal1 1196 2618 1196 2618 0 net102
rlabel metal2 21666 19805 21666 19805 0 net103
rlabel metal1 14582 7446 14582 7446 0 net104
rlabel metal1 3312 1734 3312 1734 0 net105
rlabel metal1 1288 1394 1288 1394 0 net106
rlabel metal3 3887 2244 3887 2244 0 net107
rlabel metal1 5198 2618 5198 2618 0 net108
rlabel metal1 4002 1734 4002 1734 0 net109
rlabel metal2 2622 28101 2622 28101 0 net11
rlabel metal1 4002 1836 4002 1836 0 net110
rlabel metal3 5313 1292 5313 1292 0 net111
rlabel metal1 12696 3434 12696 3434 0 net112
rlabel metal1 1978 2074 1978 2074 0 net113
rlabel metal2 1886 1241 1886 1241 0 net114
rlabel metal3 4531 9724 4531 9724 0 net115
rlabel via2 2530 1275 2530 1275 0 net116
rlabel metal2 1610 1054 1610 1054 0 net117
rlabel metal1 5566 18258 5566 18258 0 net118
rlabel metal3 16537 19380 16537 19380 0 net119
rlabel metal1 14122 21964 14122 21964 0 net12
rlabel metal1 3910 2618 3910 2618 0 net120
rlabel metal1 4876 1190 4876 1190 0 net121
rlabel metal1 7130 1972 7130 1972 0 net122
rlabel viali 7498 1943 7498 1943 0 net123
rlabel metal1 8464 2414 8464 2414 0 net124
rlabel metal1 7866 1904 7866 1904 0 net125
rlabel metal1 8924 2482 8924 2482 0 net126
rlabel metal1 7038 1326 7038 1326 0 net127
rlabel metal2 15226 17068 15226 17068 0 net128
rlabel via2 5106 1173 5106 1173 0 net129
rlabel metal1 7958 19380 7958 19380 0 net13
rlabel metal2 14398 1496 14398 1496 0 net130
rlabel metal1 4830 1972 4830 1972 0 net131
rlabel metal1 5198 1938 5198 1938 0 net132
rlabel metal1 6624 2074 6624 2074 0 net133
rlabel metal1 5658 2040 5658 2040 0 net134
rlabel metal1 6854 1938 6854 1938 0 net135
rlabel metal1 7452 1258 7452 1258 0 net136
rlabel metal1 20930 6698 20930 6698 0 net137
rlabel metal1 20562 9962 20562 9962 0 net138
rlabel metal1 24150 7378 24150 7378 0 net139
rlabel metal2 2254 18275 2254 18275 0 net14
rlabel metal1 22632 8806 22632 8806 0 net140
rlabel metal1 18998 6766 18998 6766 0 net141
rlabel metal1 21022 11730 21022 11730 0 net142
rlabel metal2 20102 5712 20102 5712 0 net143
rlabel metal1 21666 6324 21666 6324 0 net144
rlabel metal1 19729 3502 19729 3502 0 net145
rlabel metal1 20511 4114 20511 4114 0 net146
rlabel metal1 17710 10710 17710 10710 0 net147
rlabel metal1 21298 12852 21298 12852 0 net148
rlabel metal1 18032 4114 18032 4114 0 net149
rlabel metal2 5474 22338 5474 22338 0 net15
rlabel metal1 21344 5542 21344 5542 0 net150
rlabel metal1 18078 2482 18078 2482 0 net151
rlabel metal1 18814 3162 18814 3162 0 net152
rlabel metal1 11684 18394 11684 18394 0 net153
rlabel metal2 1978 39168 1978 39168 0 net154
rlabel metal1 13662 20774 13662 20774 0 net155
rlabel metal1 14168 16490 14168 16490 0 net156
rlabel metal3 17204 3536 17204 3536 0 net157
rlabel metal3 8763 32300 8763 32300 0 net158
rlabel metal3 11891 42092 11891 42092 0 net159
rlabel metal1 13938 20264 13938 20264 0 net16
rlabel metal2 14490 25636 14490 25636 0 net160
rlabel metal2 12558 42993 12558 42993 0 net161
rlabel metal3 17940 26860 17940 26860 0 net162
rlabel metal1 13202 42636 13202 42636 0 net163
rlabel metal3 13823 42908 13823 42908 0 net164
rlabel metal3 19389 21148 19389 21148 0 net165
rlabel metal1 13662 34408 13662 34408 0 net166
rlabel metal1 14628 42602 14628 42602 0 net167
rlabel metal2 14582 38573 14582 38573 0 net168
rlabel metal2 12466 18785 12466 18785 0 net169
rlabel metal1 15410 29172 15410 29172 0 net17
rlabel metal4 12604 19244 12604 19244 0 net170
rlabel metal1 15686 42534 15686 42534 0 net171
rlabel metal3 14145 9860 14145 9860 0 net172
rlabel metal2 14306 15130 14306 15130 0 net173
rlabel metal2 20838 42602 20838 42602 0 net174
rlabel metal1 18538 41786 18538 41786 0 net175
rlabel metal1 19550 41786 19550 41786 0 net176
rlabel metal1 20332 40358 20332 40358 0 net177
rlabel metal1 19412 41106 19412 41106 0 net178
rlabel metal1 19642 40494 19642 40494 0 net179
rlabel metal1 1748 20910 1748 20910 0 net18
rlabel metal1 5382 39474 5382 39474 0 net180
rlabel metal1 16882 42840 16882 42840 0 net181
rlabel metal1 14030 8466 14030 8466 0 net182
rlabel metal1 17158 42636 17158 42636 0 net183
rlabel metal1 17434 42704 17434 42704 0 net184
rlabel metal1 17802 42670 17802 42670 0 net185
rlabel metal1 17986 42704 17986 42704 0 net186
rlabel metal1 18308 42670 18308 42670 0 net187
rlabel metal1 18538 42704 18538 42704 0 net188
rlabel metal1 23920 8942 23920 8942 0 net189
rlabel metal2 2622 25840 2622 25840 0 net19
rlabel metal1 24104 7446 24104 7446 0 net190
rlabel metal1 22862 8874 22862 8874 0 net191
rlabel metal1 24150 11662 24150 11662 0 net192
rlabel metal1 20286 15130 20286 15130 0 net193
rlabel metal1 23690 16626 23690 16626 0 net194
rlabel metal1 24104 16218 24104 16218 0 net195
rlabel metal1 23138 17170 23138 17170 0 net196
rlabel metal1 18722 13464 18722 13464 0 net197
rlabel metal1 23460 14382 23460 14382 0 net198
rlabel metal1 24058 15062 24058 15062 0 net199
rlabel metal1 3910 18938 3910 18938 0 net2
rlabel metal1 13524 21862 13524 21862 0 net20
rlabel metal1 20976 19482 20976 19482 0 net200
rlabel metal1 23690 11696 23690 11696 0 net201
rlabel metal2 21160 19924 21160 19924 0 net202
rlabel metal1 24794 17510 24794 17510 0 net203
rlabel metal1 22310 16558 22310 16558 0 net204
rlabel metal1 24242 24786 24242 24786 0 net205
rlabel metal1 23230 25194 23230 25194 0 net206
rlabel metal2 21206 35292 21206 35292 0 net207
rlabel metal1 23874 26384 23874 26384 0 net208
rlabel metal1 23230 21590 23230 21590 0 net209
rlabel metal2 12190 18479 12190 18479 0 net21
rlabel metal1 23874 23086 23874 23086 0 net210
rlabel via2 18998 33541 18998 33541 0 net211
rlabel metal2 23966 24956 23966 24956 0 net212
rlabel metal2 23690 20604 23690 20604 0 net213
rlabel metal2 24150 20747 24150 20747 0 net214
rlabel metal1 21482 33830 21482 33830 0 net215
rlabel metal1 24656 22066 24656 22066 0 net216
rlabel metal2 21436 21658 21436 21658 0 net217
rlabel metal2 23414 20298 23414 20298 0 net218
rlabel metal1 24564 19346 24564 19346 0 net219
rlabel via1 7970 33422 7970 33422 0 net22
rlabel metal2 21574 21760 21574 21760 0 net220
rlabel metal1 24242 26996 24242 26996 0 net221
rlabel metal1 24242 32334 24242 32334 0 net222
rlabel metal1 23828 32538 23828 32538 0 net223
rlabel metal1 23920 33558 23920 33558 0 net224
rlabel metal1 23966 34000 23966 34000 0 net225
rlabel metal1 24150 34680 24150 34680 0 net226
rlabel metal1 23966 35122 23966 35122 0 net227
rlabel metal1 24150 35632 24150 35632 0 net228
rlabel metal1 23874 36176 23874 36176 0 net229
rlabel metal2 3726 30770 3726 30770 0 net23
rlabel metal2 22402 36516 22402 36516 0 net230
rlabel metal1 21367 36618 21367 36618 0 net231
rlabel metal1 23460 27098 23460 27098 0 net232
rlabel metal2 22954 37366 22954 37366 0 net233
rlabel metal2 23966 38794 23966 38794 0 net234
rlabel metal1 23782 38998 23782 38998 0 net235
rlabel metal2 23966 39610 23966 39610 0 net236
rlabel metal1 21114 39338 21114 39338 0 net237
rlabel metal2 19826 39491 19826 39491 0 net238
rlabel via2 20102 39899 20102 39899 0 net239
rlabel metal2 2714 34255 2714 34255 0 net24
rlabel metal1 23782 40698 23782 40698 0 net240
rlabel metal1 21390 41480 21390 41480 0 net241
rlabel metal1 21344 40358 21344 40358 0 net242
rlabel metal1 24150 27982 24150 27982 0 net243
rlabel metal1 23368 39882 23368 39882 0 net244
rlabel metal1 22632 39814 22632 39814 0 net245
rlabel metal1 23966 28628 23966 28628 0 net246
rlabel metal1 24150 29104 24150 29104 0 net247
rlabel metal1 23966 29580 23966 29580 0 net248
rlabel metal1 24150 30328 24150 30328 0 net249
rlabel metal1 11546 39950 11546 39950 0 net25
rlabel metal1 23368 30634 23368 30634 0 net250
rlabel metal1 24242 31280 24242 31280 0 net251
rlabel metal1 21873 31994 21873 31994 0 net252
rlabel metal1 20102 41990 20102 41990 0 net253
rlabel metal1 21344 40902 21344 40902 0 net254
rlabel metal1 21574 40358 21574 40358 0 net255
rlabel metal1 23828 37094 23828 37094 0 net256
rlabel metal2 21114 41242 21114 41242 0 net257
rlabel via2 21850 40171 21850 40171 0 net258
rlabel metal2 23690 34986 23690 34986 0 net259
rlabel metal1 17296 18258 17296 18258 0 net26
rlabel metal1 21068 41242 21068 41242 0 net260
rlabel metal1 22218 39814 22218 39814 0 net261
rlabel metal2 20654 41321 20654 41321 0 net262
rlabel metal1 23322 36618 23322 36618 0 net263
rlabel metal1 20608 42330 20608 42330 0 net264
rlabel metal2 20424 42364 20424 42364 0 net265
rlabel metal1 21758 42330 21758 42330 0 net266
rlabel metal1 22724 43350 22724 43350 0 net267
rlabel metal1 22310 41242 22310 41242 0 net268
rlabel metal1 20700 40698 20700 40698 0 net269
rlabel via1 13858 26962 13858 26962 0 net27
rlabel metal1 17434 43078 17434 43078 0 net270
rlabel metal1 22264 40902 22264 40902 0 net271
rlabel metal1 21390 41242 21390 41242 0 net272
rlabel metal1 10028 42534 10028 42534 0 net273
rlabel metal1 2162 42330 2162 42330 0 net274
rlabel metal1 2622 41548 2622 41548 0 net275
rlabel metal2 5842 42313 5842 42313 0 net276
rlabel metal1 2622 41752 2622 41752 0 net277
rlabel metal1 1932 41514 1932 41514 0 net278
rlabel metal1 1794 43248 1794 43248 0 net279
rlabel metal1 2944 24922 2944 24922 0 net28
rlabel metal2 8418 42296 8418 42296 0 net280
rlabel metal1 2645 41106 2645 41106 0 net281
rlabel metal1 3266 40698 3266 40698 0 net282
rlabel metal2 2530 42534 2530 42534 0 net283
rlabel metal1 3358 42330 3358 42330 0 net284
rlabel metal1 2990 41786 2990 41786 0 net285
rlabel metal2 3450 41939 3450 41939 0 net286
rlabel metal1 5106 41446 5106 41446 0 net287
rlabel metal2 3174 42432 3174 42432 0 net288
rlabel metal1 4186 41786 4186 41786 0 net289
rlabel metal1 5152 29614 5152 29614 0 net29
rlabel metal1 4922 42670 4922 42670 0 net290
rlabel metal1 4830 42228 4830 42228 0 net291
rlabel metal1 4830 41786 4830 41786 0 net292
rlabel metal1 4600 41718 4600 41718 0 net293
rlabel metal2 8970 42568 8970 42568 0 net294
rlabel metal1 9844 42330 9844 42330 0 net295
rlabel metal2 10626 43010 10626 43010 0 net296
rlabel metal1 9384 42670 9384 42670 0 net297
rlabel metal1 10028 42874 10028 42874 0 net298
rlabel metal1 10994 42840 10994 42840 0 net299
rlabel metal1 2162 16524 2162 16524 0 net3
rlabel metal1 13386 32878 13386 32878 0 net30
rlabel metal1 5888 41786 5888 41786 0 net300
rlabel metal1 5152 41718 5152 41718 0 net301
rlabel metal1 5796 41718 5796 41718 0 net302
rlabel metal1 6578 43350 6578 43350 0 net303
rlabel metal1 7268 41786 7268 41786 0 net304
rlabel metal1 7682 41786 7682 41786 0 net305
rlabel metal1 7544 41446 7544 41446 0 net306
rlabel metal2 8142 42500 8142 42500 0 net307
rlabel metal1 7820 41242 7820 41242 0 net308
rlabel metal2 9706 1802 9706 1802 0 net309
rlabel metal1 11454 21862 11454 21862 0 net31
rlabel metal1 10166 1326 10166 1326 0 net310
rlabel metal2 12466 1530 12466 1530 0 net311
rlabel metal1 14030 1972 14030 1972 0 net312
rlabel metal1 13478 1326 13478 1326 0 net313
rlabel metal1 14076 1258 14076 1258 0 net314
rlabel metal1 14352 1326 14352 1326 0 net315
rlabel metal1 14490 1972 14490 1972 0 net316
rlabel metal1 15042 1938 15042 1938 0 net317
rlabel metal1 15272 1326 15272 1326 0 net318
rlabel metal1 15686 1326 15686 1326 0 net319
rlabel metal1 5612 32878 5612 32878 0 net32
rlabel metal1 15870 2006 15870 2006 0 net320
rlabel metal1 12282 1428 12282 1428 0 net321
rlabel metal1 10902 1258 10902 1258 0 net322
rlabel metal1 11730 2006 11730 2006 0 net323
rlabel metal1 8740 1326 8740 1326 0 net324
rlabel metal1 12236 1258 12236 1258 0 net325
rlabel metal1 12144 2006 12144 2006 0 net326
rlabel metal2 13202 1904 13202 1904 0 net327
rlabel metal1 12926 1258 12926 1258 0 net328
rlabel metal2 16330 1700 16330 1700 0 net329
rlabel via1 2622 24667 2622 24667 0 net33
rlabel metal1 18308 2414 18308 2414 0 net330
rlabel metal1 18676 3094 18676 3094 0 net331
rlabel metal1 18032 4182 18032 4182 0 net332
rlabel metal1 20470 2278 20470 2278 0 net333
rlabel metal1 20792 3502 20792 3502 0 net334
rlabel metal1 21436 3094 21436 3094 0 net335
rlabel metal1 16928 1326 16928 1326 0 net336
rlabel metal1 17296 1326 17296 1326 0 net337
rlabel metal1 17710 1326 17710 1326 0 net338
rlabel metal1 17572 1938 17572 1938 0 net339
rlabel metal1 10074 36142 10074 36142 0 net34
rlabel metal1 19596 1190 19596 1190 0 net340
rlabel metal1 17572 2074 17572 2074 0 net341
rlabel metal1 17710 2006 17710 2006 0 net342
rlabel metal1 18400 1326 18400 1326 0 net343
rlabel metal1 18722 1462 18722 1462 0 net344
rlabel metal1 20562 41650 20562 41650 0 net345
rlabel metal1 1932 3162 1932 3162 0 net346
rlabel metal1 3082 5644 3082 5644 0 net347
rlabel metal1 1702 4216 1702 4216 0 net348
rlabel metal2 3818 5474 3818 5474 0 net349
rlabel metal1 15640 28526 15640 28526 0 net35
rlabel metal1 1518 3536 1518 3536 0 net350
rlabel metal1 5566 5882 5566 5882 0 net351
rlabel metal1 3542 5678 3542 5678 0 net352
rlabel metal1 2622 6358 2622 6358 0 net353
rlabel metal1 2116 3910 2116 3910 0 net354
rlabel metal1 1702 6256 1702 6256 0 net355
rlabel metal1 2162 5644 2162 5644 0 net356
rlabel metal1 1840 2822 1840 2822 0 net357
rlabel metal1 1794 6698 1794 6698 0 net358
rlabel metal1 2392 7514 2392 7514 0 net359
rlabel metal1 12880 26894 12880 26894 0 net36
rlabel metal1 2438 8908 2438 8908 0 net360
rlabel metal1 7130 8568 7130 8568 0 net361
rlabel metal1 3772 6630 3772 6630 0 net362
rlabel metal1 3174 9044 3174 9044 0 net363
rlabel metal2 1518 6290 1518 6290 0 net364
rlabel metal2 2714 5423 2714 5423 0 net365
rlabel metal2 3358 13498 3358 13498 0 net366
rlabel metal2 1978 17476 1978 17476 0 net367
rlabel metal2 1518 18207 1518 18207 0 net368
rlabel metal4 2484 18632 2484 18632 0 net369
rlabel metal1 3910 25126 3910 25126 0 net37
rlabel metal3 1909 13668 1909 13668 0 net370
rlabel metal1 3312 15062 3312 15062 0 net371
rlabel metal1 3956 14586 3956 14586 0 net372
rlabel metal1 1932 15130 1932 15130 0 net373
rlabel metal1 3680 16490 3680 16490 0 net374
rlabel metal1 7452 15470 7452 15470 0 net375
rlabel metal1 1702 16184 1702 16184 0 net376
rlabel metal1 1564 13974 1564 13974 0 net377
rlabel metal1 2852 8058 2852 8058 0 net378
rlabel metal2 2622 15096 2622 15096 0 net379
rlabel metal1 9890 32878 9890 32878 0 net38
rlabel metal1 3818 12206 3818 12206 0 net380
rlabel metal1 3680 9146 3680 9146 0 net381
rlabel metal1 2024 11118 2024 11118 0 net382
rlabel metal1 3312 7990 3312 7990 0 net383
rlabel metal2 8050 13872 8050 13872 0 net384
rlabel metal2 4416 13702 4416 13702 0 net385
rlabel metal1 2024 8942 2024 8942 0 net386
rlabel metal2 4416 10268 4416 10268 0 net387
rlabel metal2 3036 8908 3036 8908 0 net388
rlabel metal1 5244 11118 5244 11118 0 net389
rlabel via2 1610 29733 1610 29733 0 net39
rlabel metal1 1702 8874 1702 8874 0 net390
rlabel metal2 1978 12886 1978 12886 0 net391
rlabel metal2 1518 11118 1518 11118 0 net392
rlabel metal2 2070 10914 2070 10914 0 net393
rlabel metal1 14536 16558 14536 16558 0 net394
rlabel metal1 16468 19278 16468 19278 0 net395
rlabel metal2 7406 19584 7406 19584 0 net396
rlabel metal1 5198 19822 5198 19822 0 net397
rlabel metal1 15594 20978 15594 20978 0 net398
rlabel metal1 16100 23698 16100 23698 0 net399
rlabel via2 8694 16643 8694 16643 0 net4
rlabel via2 3910 28203 3910 28203 0 net40
rlabel metal1 6762 21590 6762 21590 0 net400
rlabel metal1 6854 25908 6854 25908 0 net401
rlabel metal1 14950 22066 14950 22066 0 net402
rlabel metal1 13662 17714 13662 17714 0 net403
rlabel metal2 4646 32946 4646 32946 0 net404
rlabel metal2 12742 40256 12742 40256 0 net405
rlabel metal1 11684 18258 11684 18258 0 net406
rlabel metal1 3450 39440 3450 39440 0 net407
rlabel metal1 10948 40018 10948 40018 0 net408
rlabel metal1 18400 17782 18400 17782 0 net409
rlabel metal1 1886 25398 1886 25398 0 net41
rlabel metal1 15548 31790 15548 31790 0 net42
rlabel metal2 2438 24208 2438 24208 0 net43
rlabel metal1 2369 25126 2369 25126 0 net44
rlabel metal1 9706 32946 9706 32946 0 net45
rlabel metal2 16882 26554 16882 26554 0 net46
rlabel metal2 12282 26146 12282 26146 0 net47
rlabel metal1 4416 28050 4416 28050 0 net48
rlabel metal1 20010 14892 20010 14892 0 net49
rlabel metal2 14306 19244 14306 19244 0 net5
rlabel metal1 2575 35054 2575 35054 0 net50
rlabel metal1 20102 32232 20102 32232 0 net51
rlabel metal1 2023 19346 2023 19346 0 net52
rlabel metal1 2115 18734 2115 18734 0 net53
rlabel metal1 19550 34646 19550 34646 0 net54
rlabel viali 5189 33520 5189 33520 0 net55
rlabel metal1 1702 40120 1702 40120 0 net56
rlabel metal1 14719 35666 14719 35666 0 net57
rlabel metal1 14351 31790 14351 31790 0 net58
rlabel metal1 2567 28496 2567 28496 0 net59
rlabel metal2 7866 19992 7866 19992 0 net6
rlabel metal1 19550 5168 19550 5168 0 net60
rlabel via1 1978 1987 1978 1987 0 net61
rlabel via2 2162 31773 2162 31773 0 net62
rlabel metal1 14627 20434 14627 20434 0 net63
rlabel via1 15409 21522 15409 21522 0 net64
rlabel metal1 2161 21522 2161 21522 0 net65
rlabel metal1 21758 17136 21758 17136 0 net66
rlabel metal2 21666 40239 21666 40239 0 net67
rlabel viali 2245 40048 2245 40048 0 net68
rlabel metal1 1702 9588 1702 9588 0 net69
rlabel metal1 2760 21658 2760 21658 0 net7
rlabel metal2 12650 19125 12650 19125 0 net70
rlabel metal1 1739 33490 1739 33490 0 net71
rlabel metal1 2507 40562 2507 40562 0 net72
rlabel via2 2254 41123 2254 41123 0 net73
rlabel metal1 3818 32334 3818 32334 0 net74
rlabel metal1 2438 16131 2438 16131 0 net75
rlabel metal1 14765 28526 14765 28526 0 net76
rlabel via3 21643 4012 21643 4012 0 net77
rlabel metal2 2254 35411 2254 35411 0 net78
rlabel metal1 15255 17170 15255 17170 0 net79
rlabel via1 13398 20434 13398 20434 0 net8
rlabel metal1 15447 33490 15447 33490 0 net80
rlabel metal1 1702 38828 1702 38828 0 net81
rlabel metal1 19274 10506 19274 10506 0 net82
rlabel metal2 23874 3026 23874 3026 0 net83
rlabel metal1 23690 1734 23690 1734 0 net84
rlabel via2 21206 5797 21206 5797 0 net85
rlabel metal1 18354 3706 18354 3706 0 net86
rlabel metal2 25392 21964 25392 21964 0 net87
rlabel metal2 24058 15572 24058 15572 0 net88
rlabel metal2 19504 17204 19504 17204 0 net89
rlabel metal1 1702 23562 1702 23562 0 net9
rlabel metal1 18538 1802 18538 1802 0 net90
rlabel metal2 21390 1207 21390 1207 0 net91
rlabel metal2 16422 40868 16422 40868 0 net92
rlabel metal1 16054 18836 16054 18836 0 net93
rlabel metal1 2254 19890 2254 19890 0 net94
rlabel metal1 1794 19346 1794 19346 0 net95
rlabel metal1 1518 18802 1518 18802 0 net96
rlabel metal2 20562 2057 20562 2057 0 net97
rlabel metal2 13340 19244 13340 19244 0 net98
rlabel metal1 18906 21080 18906 21080 0 net99
rlabel metal1 20194 42228 20194 42228 0 strobe_inbuf_0.X
rlabel metal1 20286 40970 20286 40970 0 strobe_inbuf_1.X
rlabel metal1 22356 12954 22356 12954 0 strobe_inbuf_10.X
rlabel metal1 25806 13940 25806 13940 0 strobe_inbuf_11.X
rlabel metal1 23552 35802 23552 35802 0 strobe_inbuf_12.X
rlabel metal2 23414 25092 23414 25092 0 strobe_inbuf_13.X
rlabel metal1 23920 21862 23920 21862 0 strobe_inbuf_14.X
rlabel metal1 23644 32878 23644 32878 0 strobe_inbuf_15.X
rlabel metal1 22632 37434 22632 37434 0 strobe_inbuf_16.X
rlabel metal1 22908 34170 22908 34170 0 strobe_inbuf_17.X
rlabel metal1 24012 36890 24012 36890 0 strobe_inbuf_18.X
rlabel metal1 23828 31994 23828 31994 0 strobe_inbuf_19.X
rlabel metal1 20562 36890 20562 36890 0 strobe_inbuf_2.X
rlabel metal1 20838 39066 20838 39066 0 strobe_inbuf_3.X
rlabel metal1 21942 41616 21942 41616 0 strobe_inbuf_4.X
rlabel metal1 21666 21658 21666 21658 0 strobe_inbuf_5.X
rlabel metal2 21528 41276 21528 41276 0 strobe_inbuf_6.X
rlabel metal1 20838 37706 20838 37706 0 strobe_inbuf_7.X
rlabel metal1 22494 39610 22494 39610 0 strobe_inbuf_8.X
rlabel metal2 22954 40885 22954 40885 0 strobe_inbuf_9.X
rlabel metal1 20470 42262 20470 42262 0 strobe_outbuf_0.X
rlabel metal2 20286 41786 20286 41786 0 strobe_outbuf_1.X
rlabel metal1 22310 39882 22310 39882 0 strobe_outbuf_10.X
rlabel metal1 21850 40460 21850 40460 0 strobe_outbuf_11.X
rlabel metal1 23506 36346 23506 36346 0 strobe_outbuf_12.X
rlabel metal2 21482 39746 21482 39746 0 strobe_outbuf_13.X
rlabel metal2 23828 38420 23828 38420 0 strobe_outbuf_14.X
rlabel metal1 23368 32742 23368 32742 0 strobe_outbuf_15.X
rlabel metal1 21850 38522 21850 38522 0 strobe_outbuf_16.X
rlabel metal1 22770 35258 22770 35258 0 strobe_outbuf_17.X
rlabel metal2 20746 39151 20746 39151 0 strobe_outbuf_18.X
rlabel metal1 24012 32198 24012 32198 0 strobe_outbuf_19.X
rlabel metal1 20562 37162 20562 37162 0 strobe_outbuf_2.X
rlabel metal1 20884 39610 20884 39610 0 strobe_outbuf_3.X
rlabel metal1 23276 40494 23276 40494 0 strobe_outbuf_4.X
rlabel metal1 22080 39610 22080 39610 0 strobe_outbuf_5.X
rlabel metal1 21344 39610 21344 39610 0 strobe_outbuf_6.X
rlabel metal1 20010 40392 20010 40392 0 strobe_outbuf_7.X
rlabel metal2 22218 40851 22218 40851 0 strobe_outbuf_8.X
rlabel metal2 22770 40868 22770 40868 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 44623
<< end >>
