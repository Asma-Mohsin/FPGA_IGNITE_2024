VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1432.120 2920.000 1432.720 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.790 3516.000 2229.070 3520.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.950 3516.000 1905.230 3520.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 3516.000 1581.390 3520.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 3516.000 1257.550 3520.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 3516.000 933.710 3520.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 3516.000 609.870 3520.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 3516.000 286.030 3520.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3453.080 4.000 3453.680 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3197.400 4.000 3198.000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2941.720 4.000 2942.320 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1693.240 2920.000 1693.840 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2686.040 4.000 2686.640 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2430.360 4.000 2430.960 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2174.680 4.000 2175.280 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1919.000 4.000 1919.600 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1663.320 4.000 1663.920 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1407.640 4.000 1408.240 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.280 4.000 896.880 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1954.360 2920.000 1954.960 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2215.480 2920.000 2216.080 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2476.600 2920.000 2477.200 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2737.720 2920.000 2738.320 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2998.840 2920.000 2999.440 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3259.960 2920.000 3260.560 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.470 3516.000 2876.750 3520.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2552.630 3516.000 2552.910 3520.000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 61.240 2920.000 61.840 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2280.760 2920.000 2281.360 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2541.880 2920.000 2542.480 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2803.000 2920.000 2803.600 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3064.120 2920.000 3064.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3325.240 2920.000 3325.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 2795.510 3516.000 2795.790 3520.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2471.670 3516.000 2471.950 3520.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 2147.830 3516.000 2148.110 3520.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1823.990 3516.000 1824.270 3520.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1500.150 3516.000 1500.430 3520.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 257.080 2920.000 257.680 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1176.310 3516.000 1176.590 3520.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 852.470 3516.000 852.750 3520.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 528.630 3516.000 528.910 3520.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 204.790 3516.000 205.070 3520.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3389.160 4.000 3389.760 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3133.480 4.000 3134.080 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2877.800 4.000 2878.400 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2622.120 4.000 2622.720 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2366.440 4.000 2367.040 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2110.760 4.000 2111.360 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 452.920 2920.000 453.520 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1855.080 4.000 1855.680 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1599.400 4.000 1600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.720 4.000 1344.320 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 648.760 2920.000 649.360 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 844.600 2920.000 845.200 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1040.440 2920.000 1041.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1236.280 2920.000 1236.880 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1497.400 2920.000 1498.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1758.520 2920.000 1759.120 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2019.640 2920.000 2020.240 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 191.800 2920.000 192.400 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2411.320 2920.000 2411.920 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2672.440 2920.000 2673.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2933.560 2920.000 2934.160 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3194.680 2920.000 3195.280 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3455.800 2920.000 3456.400 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2633.590 3516.000 2633.870 3520.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2309.750 3516.000 2310.030 3520.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1985.910 3516.000 1986.190 3520.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1662.070 3516.000 1662.350 3520.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1338.230 3516.000 1338.510 3520.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 387.640 2920.000 388.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1014.390 3516.000 1014.670 3520.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 690.550 3516.000 690.830 3520.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 366.710 3516.000 366.990 3520.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 42.870 3516.000 43.150 3520.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3261.320 4.000 3261.920 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3005.640 4.000 3006.240 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2749.960 4.000 2750.560 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2494.280 4.000 2494.880 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2238.600 4.000 2239.200 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1982.920 4.000 1983.520 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 583.480 2920.000 584.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1471.560 4.000 1472.160 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.880 4.000 1216.480 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 779.320 2920.000 779.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 975.160 2920.000 975.760 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1171.000 2920.000 1171.600 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1366.840 2920.000 1367.440 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1627.960 2920.000 1628.560 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1889.080 2920.000 1889.680 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2150.200 2920.000 2150.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 126.520 2920.000 127.120 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2346.040 2920.000 2346.640 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2607.160 2920.000 2607.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2868.280 2920.000 2868.880 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3129.400 2920.000 3130.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 2916.000 3390.520 2920.000 3391.120 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2714.550 3516.000 2714.830 3520.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2390.710 3516.000 2390.990 3520.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2066.870 3516.000 2067.150 3520.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1743.030 3516.000 1743.310 3520.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1419.190 3516.000 1419.470 3520.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 322.360 2920.000 322.960 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1095.350 3516.000 1095.630 3520.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 771.510 3516.000 771.790 3520.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 447.670 3516.000 447.950 3520.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 123.830 3516.000 124.110 3520.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3325.240 4.000 3325.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 3069.560 4.000 3070.160 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2813.880 4.000 2814.480 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2558.200 4.000 2558.800 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2302.520 4.000 2303.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2046.840 4.000 2047.440 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 518.200 2920.000 518.800 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1791.160 4.000 1791.760 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1535.480 4.000 1536.080 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.800 4.000 1280.400 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 714.040 2920.000 714.640 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 909.880 2920.000 910.480 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1105.720 2920.000 1106.320 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1301.560 2920.000 1302.160 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1562.680 2920.000 1563.280 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 1823.800 2920.000 1824.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2916.000 2084.920 2920.000 2085.520 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.110 0.000 2340.390 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.670 0.000 2356.950 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2373.230 0.000 2373.510 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2389.790 0.000 2390.070 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2406.350 0.000 2406.630 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2422.910 0.000 2423.190 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2439.470 0.000 2439.750 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2456.030 0.000 2456.310 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2472.590 0.000 2472.870 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.150 0.000 2489.430 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.710 0.000 2505.990 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.270 0.000 2522.550 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.830 0.000 2539.110 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.390 0.000 2555.670 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.950 0.000 2572.230 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.510 0.000 2588.790 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2605.070 0.000 2605.350 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.630 0.000 2621.910 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.190 0.000 2638.470 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.750 0.000 2655.030 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 0.000 866.550 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.310 0.000 2671.590 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.870 0.000 2688.150 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.430 0.000 2704.710 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.990 0.000 2721.270 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2737.550 0.000 2737.830 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2754.110 0.000 2754.390 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.670 0.000 2770.950 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2787.230 0.000 2787.510 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.390 0.000 899.670 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.310 0.000 1015.590 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.870 0.000 1032.150 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.550 0.000 1081.830 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.110 0.000 1098.390 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.670 0.000 1114.950 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 0.000 1131.510 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.910 0.000 1181.190 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.470 0.000 1197.750 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.030 0.000 1214.310 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 0.000 1230.870 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.710 0.000 1263.990 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.270 0.000 1280.550 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.390 0.000 1313.670 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1346.510 0.000 1346.790 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1379.630 0.000 1379.910 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1396.190 0.000 1396.470 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1429.310 0.000 1429.590 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1445.870 0.000 1446.150 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1462.430 0.000 1462.710 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1478.990 0.000 1479.270 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1495.550 0.000 1495.830 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1512.110 0.000 1512.390 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1528.670 0.000 1528.950 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1545.230 0.000 1545.510 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1561.790 0.000 1562.070 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1578.350 0.000 1578.630 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1594.910 0.000 1595.190 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1628.030 0.000 1628.310 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1644.590 0.000 1644.870 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1661.150 0.000 1661.430 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 0.000 767.190 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1694.270 0.000 1694.550 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1710.830 0.000 1711.110 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1727.390 0.000 1727.670 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1743.950 0.000 1744.230 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1760.510 0.000 1760.790 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1777.070 0.000 1777.350 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1793.630 0.000 1793.910 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1810.190 0.000 1810.470 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1826.750 0.000 1827.030 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1843.310 0.000 1843.590 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1859.870 0.000 1860.150 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1876.430 0.000 1876.710 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1892.990 0.000 1893.270 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1926.110 0.000 1926.390 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1942.670 0.000 1942.950 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1959.230 0.000 1959.510 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 1975.790 0.000 1976.070 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 1992.350 0.000 1992.630 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2008.910 0.000 2009.190 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2025.470 0.000 2025.750 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2042.030 0.000 2042.310 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 2058.590 0.000 2058.870 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.150 0.000 2075.430 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.710 0.000 2091.990 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.270 0.000 2108.550 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.830 0.000 2125.110 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 0.000 2141.670 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2157.950 0.000 2158.230 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 816.590 0.000 816.870 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2174.510 0.000 2174.790 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2191.070 0.000 2191.350 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.630 0.000 2207.910 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.190 0.000 2224.470 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.750 0.000 2241.030 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.310 0.000 2257.590 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.870 0.000 2274.150 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.430 0.000 2290.710 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.990 0.000 2307.270 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.550 0.000 2323.830 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.630 0.000 2345.910 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.190 0.000 2362.470 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.750 0.000 2379.030 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.310 0.000 2395.590 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.870 0.000 2412.150 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.430 0.000 2428.710 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.990 0.000 2445.270 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.550 0.000 2461.830 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2478.110 0.000 2478.390 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.670 0.000 2494.950 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.230 0.000 2511.510 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.790 0.000 2528.070 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.350 0.000 2544.630 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.910 0.000 2561.190 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.470 0.000 2577.750 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2594.030 0.000 2594.310 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2610.590 0.000 2610.870 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.150 0.000 2627.430 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.710 0.000 2643.990 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.270 0.000 2660.550 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.830 0.000 2677.110 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.390 0.000 2693.670 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.950 0.000 2710.230 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.510 0.000 2726.790 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2743.070 0.000 2743.350 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.630 0.000 2759.910 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2776.190 0.000 2776.470 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 2792.750 0.000 2793.030 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 888.350 0.000 888.630 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 904.910 0.000 905.190 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 954.590 0.000 954.870 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.150 0.000 971.430 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.270 0.000 1004.550 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 0.000 1037.670 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.950 0.000 1054.230 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.070 0.000 1087.350 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 0.000 1103.910 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.750 0.000 1137.030 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 0.000 1170.150 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 722.750 0.000 723.030 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.430 0.000 1186.710 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.990 0.000 1203.270 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.550 0.000 1219.830 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1236.110 0.000 1236.390 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.670 0.000 1252.950 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1269.230 0.000 1269.510 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1285.790 0.000 1286.070 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1335.470 0.000 1335.750 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.030 0.000 1352.310 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.710 0.000 1401.990 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 0.000 1418.550 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 0.000 1435.110 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 0.000 1451.670 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.950 0.000 1468.230 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 0.000 1484.790 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.070 0.000 1501.350 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.630 0.000 1517.910 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.190 0.000 1534.470 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.750 0.000 1551.030 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.310 0.000 1567.590 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 0.000 1584.150 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.430 0.000 1600.710 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.990 0.000 1617.270 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.550 0.000 1633.830 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 0.000 1650.390 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.670 0.000 1666.950 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.230 0.000 1683.510 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.790 0.000 1700.070 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.350 0.000 1716.630 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.910 0.000 1733.190 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.470 0.000 1749.750 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.590 0.000 1782.870 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.150 0.000 1799.430 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.710 0.000 1815.990 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 0.000 1832.550 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.830 0.000 1849.110 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.390 0.000 1865.670 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.950 0.000 1882.230 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.510 0.000 1898.790 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.070 0.000 1915.350 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.630 0.000 1931.910 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.190 0.000 1948.470 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.310 0.000 1981.590 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.870 0.000 1998.150 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.430 0.000 2014.710 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.990 0.000 2031.270 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.550 0.000 2047.830 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.670 0.000 2080.950 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.230 0.000 2097.510 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.790 0.000 2114.070 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.350 0.000 2130.630 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.910 0.000 2147.190 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.470 0.000 2163.750 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.030 0.000 2180.310 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.590 0.000 2196.870 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.150 0.000 2213.430 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.710 0.000 2229.990 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.270 0.000 2246.550 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.830 0.000 2263.110 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.390 0.000 2279.670 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.950 0.000 2296.230 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.510 0.000 2312.790 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2329.070 0.000 2329.350 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.150 0.000 2351.430 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.710 0.000 2367.990 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.270 0.000 2384.550 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2400.830 0.000 2401.110 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.390 0.000 2417.670 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.950 0.000 2434.230 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.510 0.000 2450.790 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.070 0.000 2467.350 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.630 0.000 2483.910 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.190 0.000 2500.470 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.750 0.000 861.030 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.750 0.000 2517.030 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.310 0.000 2533.590 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.870 0.000 2550.150 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.430 0.000 2566.710 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.990 0.000 2583.270 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.550 0.000 2599.830 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2616.110 0.000 2616.390 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.670 0.000 2632.950 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.230 0.000 2649.510 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.790 0.000 2666.070 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.310 0.000 877.590 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.350 0.000 2682.630 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.910 0.000 2699.190 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.470 0.000 2715.750 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.030 0.000 2732.310 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.590 0.000 2748.870 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.150 0.000 2765.430 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.710 0.000 2781.990 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.270 0.000 2798.550 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 0.000 894.150 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.110 0.000 960.390 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 0.000 976.950 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.910 0.000 1043.190 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.030 0.000 1076.310 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 0.000 1092.870 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.150 0.000 1109.430 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.710 0.000 1125.990 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 0.000 1159.110 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 0.000 1208.790 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.070 0.000 1225.350 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.630 0.000 1241.910 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.190 0.000 1258.470 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.750 0.000 1275.030 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.310 0.000 1291.590 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 0.000 1308.150 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.430 0.000 1324.710 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 0.000 1341.270 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.670 0.000 1390.950 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 0.000 1407.510 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.790 0.000 1424.070 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.350 0.000 1440.630 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.470 0.000 1473.750 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.030 0.000 1490.310 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.590 0.000 1506.870 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 0.000 1523.430 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.710 0.000 1539.990 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.270 0.000 1556.550 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.830 0.000 1573.110 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.390 0.000 1589.670 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 0.000 1606.230 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 0.000 1622.790 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.070 0.000 1639.350 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.630 0.000 1655.910 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.750 0.000 1689.030 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.310 0.000 1705.590 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 0.000 1722.150 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.430 0.000 1738.710 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.990 0.000 1755.270 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.550 0.000 1771.830 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1788.110 0.000 1788.390 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.670 0.000 1804.950 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.230 0.000 1821.510 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.790 0.000 1838.070 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.350 0.000 1854.630 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.910 0.000 1871.190 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 0.000 1887.750 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.030 0.000 1904.310 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.590 0.000 1920.870 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.150 0.000 1937.430 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.710 0.000 1953.990 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.270 0.000 1970.550 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.390 0.000 2003.670 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.950 0.000 2020.230 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.510 0.000 2036.790 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.070 0.000 2053.350 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.190 0.000 2086.470 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.750 0.000 2103.030 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.310 0.000 2119.590 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.870 0.000 2136.150 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.430 0.000 2152.710 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.990 0.000 2169.270 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.550 0.000 2185.830 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.110 0.000 2202.390 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.230 0.000 2235.510 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.790 0.000 2252.070 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.350 0.000 2268.630 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.910 0.000 2285.190 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.470 0.000 2301.750 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2318.030 0.000 2318.310 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.590 0.000 2334.870 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 0.000 844.470 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2803.790 0.000 2804.070 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.310 0.000 2809.590 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2814.830 0.000 2815.110 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2820.350 0.000 2820.630 4.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 3525.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 -6.220 2931.200 -3.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 3522.800 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.100 -6.220 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 4.020 -11.020 7.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.020 -11.020 57.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.020 2619.480 57.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.020 -11.020 107.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.020 2619.480 107.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.020 -11.020 157.020 404.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.020 1938.440 157.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.020 2619.480 157.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.020 -11.020 207.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.020 2619.480 207.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 -11.020 257.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 1940.065 257.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.020 2620.100 257.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.020 -11.020 307.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.020 1995.920 307.020 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.020 2619.480 307.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.020 -11.020 357.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.020 1979.185 357.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.020 2620.100 357.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 -11.020 407.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 1940.065 407.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.020 2619.480 407.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.020 -11.020 457.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.020 2619.480 457.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.020 -11.020 507.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.020 1940.065 507.020 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.020 2619.480 507.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.020 -11.020 557.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.020 1995.920 557.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.020 -11.020 607.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.020 1979.185 607.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.020 -11.020 657.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 654.020 1940.065 657.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 704.020 -11.020 707.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 754.020 -11.020 757.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 754.020 1940.065 757.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 804.020 -11.020 807.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 804.020 1995.920 807.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.020 -11.020 857.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.020 1979.185 857.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.020 -11.020 907.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 904.020 1940.065 907.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.020 -11.020 957.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 954.020 1940.065 957.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1004.020 -11.020 1007.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1004.020 1995.920 1007.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.020 -11.020 1057.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1054.020 1979.185 1057.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.020 -11.020 1107.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1104.020 1979.185 1107.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1154.020 -11.020 1157.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1154.020 1940.065 1157.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1204.020 -11.020 1207.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1204.020 1940.065 1207.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.020 -11.020 1257.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1254.020 1940.065 1257.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.020 -11.020 1307.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1304.020 1995.920 1307.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1354.020 -11.020 1357.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1354.020 1995.920 1357.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1404.020 -11.020 1407.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1404.020 1940.065 1407.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.020 -11.020 1457.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.020 1940.065 1457.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.020 -11.020 1507.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1504.020 1940.065 1507.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.020 -11.020 1557.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.020 1979.185 1557.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.020 -11.020 1607.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.020 1940.065 1607.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.020 -11.020 1657.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1654.020 1995.920 1657.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.020 -11.020 1707.020 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1704.020 1995.920 1707.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.020 -11.020 1757.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1754.020 1979.185 1757.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.020 -11.020 1807.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1804.020 1979.185 1807.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.020 -11.020 1857.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1854.020 1940.065 1857.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.020 -11.020 1907.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.020 1940.065 1907.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.020 -11.020 1957.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.020 1940.065 1957.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.020 -11.020 2007.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2004.020 1940.065 2007.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.020 -11.020 2057.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2054.020 1979.185 2057.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.020 -11.020 2107.020 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 2104.020 1940.065 2107.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.020 -11.020 2157.020 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.020 1940.065 2157.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2204.020 -11.020 2207.020 339.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2204.020 1995.480 2207.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.020 -11.020 2257.020 405.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.020 1994.385 2257.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.020 -11.020 2307.020 339.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2304.020 1995.480 2307.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2354.020 -11.020 2357.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 -11.020 2407.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 859.380 2407.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 1379.480 2407.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2404.020 1899.480 2407.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 -11.020 2457.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 859.380 2457.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 1379.480 2457.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2454.020 1899.480 2457.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 -11.020 2507.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 859.380 2507.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 1379.480 2507.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.020 1899.480 2507.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 -11.020 2557.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 860.100 2557.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 1380.100 2557.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2554.020 1900.100 2557.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 -11.020 2607.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 860.100 2607.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 1380.100 2607.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.020 1900.100 2607.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 -11.020 2657.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 860.100 2657.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 1380.100 2657.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2654.020 1900.100 2657.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 -11.020 2707.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 860.100 2707.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 1380.100 2707.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2704.020 1900.100 2707.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 -11.020 2757.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 859.380 2757.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 1379.480 2757.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2754.020 1899.480 2757.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 -11.020 2807.020 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 859.380 2807.020 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 1379.480 2807.020 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2804.020 1899.480 2807.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 -11.020 2857.020 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 859.380 2857.020 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 1379.480 2857.020 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2854.020 1899.480 2857.020 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2904.020 -11.020 2907.020 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 9.380 2936.000 12.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 59.380 2936.000 62.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 109.380 2936.000 112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 159.380 2936.000 162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 209.380 2936.000 212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 259.380 2936.000 262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 309.380 2936.000 312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 359.380 2936.000 362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 409.380 2936.000 412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 459.380 2936.000 462.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 509.380 2936.000 512.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 559.380 2936.000 562.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 609.380 2936.000 612.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 659.380 2936.000 662.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 709.380 2936.000 712.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 759.380 2936.000 762.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 809.380 2936.000 812.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 859.380 2936.000 862.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 909.380 2936.000 912.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 959.380 2936.000 962.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1009.380 2936.000 1012.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1059.380 2936.000 1062.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1109.380 2936.000 1112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1159.380 2936.000 1162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1209.380 2936.000 1212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1259.380 2936.000 1262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1309.380 2936.000 1312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1359.380 2936.000 1362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1409.380 2936.000 1412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1459.380 2936.000 1462.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1509.380 2936.000 1512.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1559.380 2936.000 1562.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1609.380 2936.000 1612.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1659.380 2936.000 1662.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1709.380 2936.000 1712.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1759.380 2936.000 1762.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1809.380 2936.000 1812.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1859.380 2936.000 1862.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1909.380 2936.000 1912.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1959.380 2936.000 1962.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2009.380 2936.000 2012.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2059.380 2936.000 2062.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2109.380 2936.000 2112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2159.380 2936.000 2162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2209.380 2936.000 2212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2259.380 2936.000 2262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2309.380 2936.000 2312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2359.380 2936.000 2362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2409.380 2936.000 2412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2459.380 2936.000 2462.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2509.380 2936.000 2512.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2559.380 2936.000 2562.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2609.380 2936.000 2612.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2659.380 2936.000 2662.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2709.380 2936.000 2712.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2759.380 2936.000 2762.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2809.380 2936.000 2812.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2859.380 2936.000 2862.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2909.380 2936.000 2912.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2959.380 2936.000 2962.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3009.380 2936.000 3012.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3059.380 2936.000 3062.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3109.380 2936.000 3112.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3159.380 2936.000 3162.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3209.380 2936.000 3212.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3259.380 2936.000 3262.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3309.380 2936.000 3312.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3359.380 2936.000 3362.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3409.380 2936.000 3412.380 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3459.380 2936.000 3462.380 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 -11.020 2936.000 -7.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3527.600 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2932.900 -11.020 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.720 -11.020 11.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.720 -11.020 61.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.720 2619.480 61.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.720 -11.020 111.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.720 2619.480 111.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 -11.020 161.720 408.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 1931.225 161.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 158.720 2619.480 161.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 -11.020 211.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 1940.065 211.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 208.720 2620.100 211.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.720 -11.020 261.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.720 1940.065 261.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 258.720 2620.100 261.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.720 -11.020 311.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.720 1979.185 311.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 308.720 2620.100 311.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.720 -11.020 361.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.720 1995.920 361.720 2201.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 358.720 2620.100 361.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.720 -11.020 411.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.720 1940.065 411.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 408.720 2619.480 411.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.720 -11.020 461.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.720 1940.065 461.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.720 2619.480 461.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.720 -11.020 511.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.720 1940.065 511.720 2202.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 508.720 2619.480 511.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.720 -11.020 561.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.720 1979.185 561.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.720 -11.020 611.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 608.720 1995.920 611.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.720 -11.020 661.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 658.720 1940.065 661.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.720 -11.020 711.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 708.720 1940.065 711.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.720 -11.020 761.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 758.720 1940.065 761.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.720 -11.020 811.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 808.720 1979.185 811.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 -11.020 861.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 858.720 1995.920 861.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 -11.020 911.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.720 1940.065 911.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 958.720 -11.020 961.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 958.720 1940.065 961.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.720 -11.020 1011.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1008.720 1940.065 1011.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.720 -11.020 1061.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1058.720 1995.920 1061.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.720 -11.020 1111.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1108.720 1979.185 1111.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.720 -11.020 1161.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1158.720 1940.065 1161.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.720 -11.020 1211.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1208.720 1940.065 1211.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.720 -11.020 1261.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1258.720 1940.065 1261.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.720 -11.020 1311.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1308.720 1979.185 1311.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.720 -11.020 1361.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.720 1995.920 1361.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.720 -11.020 1411.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1408.720 1995.920 1411.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.720 -11.020 1461.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1458.720 1940.065 1461.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.720 -11.020 1511.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1508.720 1940.065 1511.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.720 -11.020 1561.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1558.720 1979.185 1561.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.720 -11.020 1611.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.720 1940.065 1611.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.720 -11.020 1661.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1658.720 1940.065 1661.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1708.720 -11.020 1711.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1708.720 1940.065 1711.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.720 -11.020 1761.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1758.720 1995.920 1761.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.720 -11.020 1811.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.720 1979.185 1811.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.720 -11.020 1861.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 1858.720 1940.065 1861.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1908.720 -11.020 1911.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.720 -11.020 1961.720 345.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.720 1995.920 1961.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.720 -11.020 2011.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2008.720 1979.185 2011.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.720 -11.020 2061.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2058.720 1979.185 2061.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.720 -11.020 2111.720 353.615 ;
    END
    PORT
      LAYER met4 ;
        RECT 2108.720 1940.065 2111.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.720 -11.020 2161.720 400.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 2158.720 1940.065 2161.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.720 -11.020 2211.720 405.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2208.720 1935.305 2211.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.720 -11.020 2261.720 405.015 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.720 1994.385 2261.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.720 -11.020 2311.720 339.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2308.720 1995.480 2311.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2358.720 -11.020 2361.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 -11.020 2411.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 859.480 2411.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 1379.480 2411.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2408.720 1899.480 2411.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 -11.020 2461.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 859.480 2461.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 1379.480 2461.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2458.720 1899.480 2461.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 -11.020 2511.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 859.480 2511.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 1379.480 2511.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2508.720 1899.480 2511.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 -11.020 2561.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 860.100 2561.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 1380.100 2561.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2558.720 1900.100 2561.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 -11.020 2611.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 860.100 2611.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 1380.100 2611.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2608.720 1900.100 2611.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 -11.020 2661.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 860.100 2661.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 1380.100 2661.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2658.720 1900.100 2661.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 -11.020 2711.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 860.100 2711.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 1380.100 2711.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.720 1900.100 2711.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 -11.020 2761.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 859.480 2761.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 1379.480 2761.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2758.720 1899.480 2761.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 -11.020 2811.720 441.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 859.480 2811.720 961.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 1379.480 2811.720 1481.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2808.720 1899.480 2811.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 -11.020 2861.720 442.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 859.480 2861.720 962.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 1379.480 2861.720 1482.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2858.720 1899.480 2861.720 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2908.720 -11.020 2911.720 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 14.080 2936.000 17.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 64.080 2936.000 67.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 114.080 2936.000 117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 164.080 2936.000 167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 214.080 2936.000 217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 264.080 2936.000 267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 314.080 2936.000 317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 364.080 2936.000 367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 414.080 2936.000 417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 464.080 2936.000 467.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 514.080 2936.000 517.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 564.080 2936.000 567.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 614.080 2936.000 617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 664.080 2936.000 667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 714.080 2936.000 717.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 764.080 2936.000 767.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 814.080 2936.000 817.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 864.080 2936.000 867.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 914.080 2936.000 917.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 964.080 2936.000 967.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1014.080 2936.000 1017.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1064.080 2936.000 1067.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1114.080 2936.000 1117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1164.080 2936.000 1167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1214.080 2936.000 1217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1264.080 2936.000 1267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1314.080 2936.000 1317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1364.080 2936.000 1367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1414.080 2936.000 1417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1464.080 2936.000 1467.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1514.080 2936.000 1517.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1564.080 2936.000 1567.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1614.080 2936.000 1617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1664.080 2936.000 1667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1714.080 2936.000 1717.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1764.080 2936.000 1767.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1814.080 2936.000 1817.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1864.080 2936.000 1867.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1914.080 2936.000 1917.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 1964.080 2936.000 1967.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2014.080 2936.000 2017.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2064.080 2936.000 2067.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2114.080 2936.000 2117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2164.080 2936.000 2167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2214.080 2936.000 2217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2264.080 2936.000 2267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2314.080 2936.000 2317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2364.080 2936.000 2367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2414.080 2936.000 2417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2464.080 2936.000 2467.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2514.080 2936.000 2517.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2564.080 2936.000 2567.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2614.080 2936.000 2617.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2664.080 2936.000 2667.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2714.080 2936.000 2717.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2764.080 2936.000 2767.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2814.080 2936.000 2817.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2864.080 2936.000 2867.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2914.080 2936.000 2917.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 2964.080 2936.000 2967.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3014.080 2936.000 3017.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3064.080 2936.000 3067.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3114.080 2936.000 3117.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3164.080 2936.000 3167.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3214.080 2936.000 3217.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3264.080 2936.000 3267.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3314.080 2936.000 3317.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3364.080 2936.000 3367.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3414.080 2936.000 3417.080 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3464.080 2936.000 3467.080 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 336.350 0.000 336.630 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 667.550 0.000 667.830 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 590.270 0.000 590.550 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 0.000 331.110 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 0.000 513.270 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 0.000 612.630 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 0.000 645.750 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 0.990 0.380 2917.250 3509.040 ;
      LAYER met2 ;
        RECT 1.020 3515.720 42.590 3516.690 ;
        RECT 43.430 3515.720 123.550 3516.690 ;
        RECT 124.390 3515.720 204.510 3516.690 ;
        RECT 205.350 3515.720 285.470 3516.690 ;
        RECT 286.310 3515.720 366.430 3516.690 ;
        RECT 367.270 3515.720 447.390 3516.690 ;
        RECT 448.230 3515.720 528.350 3516.690 ;
        RECT 529.190 3515.720 609.310 3516.690 ;
        RECT 610.150 3515.720 690.270 3516.690 ;
        RECT 691.110 3515.720 771.230 3516.690 ;
        RECT 772.070 3515.720 852.190 3516.690 ;
        RECT 853.030 3515.720 933.150 3516.690 ;
        RECT 933.990 3515.720 1014.110 3516.690 ;
        RECT 1014.950 3515.720 1095.070 3516.690 ;
        RECT 1095.910 3515.720 1176.030 3516.690 ;
        RECT 1176.870 3515.720 1256.990 3516.690 ;
        RECT 1257.830 3515.720 1337.950 3516.690 ;
        RECT 1338.790 3515.720 1418.910 3516.690 ;
        RECT 1419.750 3515.720 1499.870 3516.690 ;
        RECT 1500.710 3515.720 1580.830 3516.690 ;
        RECT 1581.670 3515.720 1661.790 3516.690 ;
        RECT 1662.630 3515.720 1742.750 3516.690 ;
        RECT 1743.590 3515.720 1823.710 3516.690 ;
        RECT 1824.550 3515.720 1904.670 3516.690 ;
        RECT 1905.510 3515.720 1985.630 3516.690 ;
        RECT 1986.470 3515.720 2066.590 3516.690 ;
        RECT 2067.430 3515.720 2147.550 3516.690 ;
        RECT 2148.390 3515.720 2228.510 3516.690 ;
        RECT 2229.350 3515.720 2309.470 3516.690 ;
        RECT 2310.310 3515.720 2390.430 3516.690 ;
        RECT 2391.270 3515.720 2471.390 3516.690 ;
        RECT 2472.230 3515.720 2552.350 3516.690 ;
        RECT 2553.190 3515.720 2633.310 3516.690 ;
        RECT 2634.150 3515.720 2714.270 3516.690 ;
        RECT 2715.110 3515.720 2795.230 3516.690 ;
        RECT 2796.070 3515.720 2876.190 3516.690 ;
        RECT 2877.030 3515.720 2917.220 3516.690 ;
        RECT 1.020 4.280 2917.220 3515.720 ;
        RECT 1.020 0.350 98.710 4.280 ;
        RECT 99.550 0.350 104.230 4.280 ;
        RECT 105.070 0.350 109.750 4.280 ;
        RECT 110.590 0.350 115.270 4.280 ;
        RECT 116.110 0.350 120.790 4.280 ;
        RECT 121.630 0.350 126.310 4.280 ;
        RECT 127.150 0.350 131.830 4.280 ;
        RECT 132.670 0.350 137.350 4.280 ;
        RECT 138.190 0.350 142.870 4.280 ;
        RECT 143.710 0.350 148.390 4.280 ;
        RECT 149.230 0.350 153.910 4.280 ;
        RECT 154.750 0.350 159.430 4.280 ;
        RECT 160.270 0.350 164.950 4.280 ;
        RECT 165.790 0.350 170.470 4.280 ;
        RECT 171.310 0.350 175.990 4.280 ;
        RECT 176.830 0.350 181.510 4.280 ;
        RECT 182.350 0.350 187.030 4.280 ;
        RECT 187.870 0.350 192.550 4.280 ;
        RECT 193.390 0.350 198.070 4.280 ;
        RECT 198.910 0.350 203.590 4.280 ;
        RECT 204.430 0.350 209.110 4.280 ;
        RECT 209.950 0.350 214.630 4.280 ;
        RECT 215.470 0.350 220.150 4.280 ;
        RECT 220.990 0.350 225.670 4.280 ;
        RECT 226.510 0.350 231.190 4.280 ;
        RECT 232.030 0.350 236.710 4.280 ;
        RECT 237.550 0.350 242.230 4.280 ;
        RECT 243.070 0.350 247.750 4.280 ;
        RECT 248.590 0.350 253.270 4.280 ;
        RECT 254.110 0.350 258.790 4.280 ;
        RECT 259.630 0.350 264.310 4.280 ;
        RECT 265.150 0.350 269.830 4.280 ;
        RECT 270.670 0.350 275.350 4.280 ;
        RECT 276.190 0.350 280.870 4.280 ;
        RECT 281.710 0.350 286.390 4.280 ;
        RECT 287.230 0.350 291.910 4.280 ;
        RECT 292.750 0.350 297.430 4.280 ;
        RECT 298.270 0.350 302.950 4.280 ;
        RECT 303.790 0.350 308.470 4.280 ;
        RECT 309.310 0.350 313.990 4.280 ;
        RECT 314.830 0.350 319.510 4.280 ;
        RECT 320.350 0.350 325.030 4.280 ;
        RECT 325.870 0.350 330.550 4.280 ;
        RECT 331.390 0.350 336.070 4.280 ;
        RECT 336.910 0.350 341.590 4.280 ;
        RECT 342.430 0.350 347.110 4.280 ;
        RECT 347.950 0.350 352.630 4.280 ;
        RECT 353.470 0.350 358.150 4.280 ;
        RECT 358.990 0.350 363.670 4.280 ;
        RECT 364.510 0.350 369.190 4.280 ;
        RECT 370.030 0.350 374.710 4.280 ;
        RECT 375.550 0.350 380.230 4.280 ;
        RECT 381.070 0.350 385.750 4.280 ;
        RECT 386.590 0.350 391.270 4.280 ;
        RECT 392.110 0.350 396.790 4.280 ;
        RECT 397.630 0.350 402.310 4.280 ;
        RECT 403.150 0.350 407.830 4.280 ;
        RECT 408.670 0.350 413.350 4.280 ;
        RECT 414.190 0.350 418.870 4.280 ;
        RECT 419.710 0.350 424.390 4.280 ;
        RECT 425.230 0.350 429.910 4.280 ;
        RECT 430.750 0.350 435.430 4.280 ;
        RECT 436.270 0.350 440.950 4.280 ;
        RECT 441.790 0.350 446.470 4.280 ;
        RECT 447.310 0.350 451.990 4.280 ;
        RECT 452.830 0.350 457.510 4.280 ;
        RECT 458.350 0.350 463.030 4.280 ;
        RECT 463.870 0.350 468.550 4.280 ;
        RECT 469.390 0.350 474.070 4.280 ;
        RECT 474.910 0.350 479.590 4.280 ;
        RECT 480.430 0.350 485.110 4.280 ;
        RECT 485.950 0.350 490.630 4.280 ;
        RECT 491.470 0.350 496.150 4.280 ;
        RECT 496.990 0.350 501.670 4.280 ;
        RECT 502.510 0.350 507.190 4.280 ;
        RECT 508.030 0.350 512.710 4.280 ;
        RECT 513.550 0.350 518.230 4.280 ;
        RECT 519.070 0.350 523.750 4.280 ;
        RECT 524.590 0.350 529.270 4.280 ;
        RECT 530.110 0.350 534.790 4.280 ;
        RECT 535.630 0.350 540.310 4.280 ;
        RECT 541.150 0.350 545.830 4.280 ;
        RECT 546.670 0.350 551.350 4.280 ;
        RECT 552.190 0.350 556.870 4.280 ;
        RECT 557.710 0.350 562.390 4.280 ;
        RECT 563.230 0.350 567.910 4.280 ;
        RECT 568.750 0.350 573.430 4.280 ;
        RECT 574.270 0.350 578.950 4.280 ;
        RECT 579.790 0.350 584.470 4.280 ;
        RECT 585.310 0.350 589.990 4.280 ;
        RECT 590.830 0.350 595.510 4.280 ;
        RECT 596.350 0.350 601.030 4.280 ;
        RECT 601.870 0.350 606.550 4.280 ;
        RECT 607.390 0.350 612.070 4.280 ;
        RECT 612.910 0.350 617.590 4.280 ;
        RECT 618.430 0.350 623.110 4.280 ;
        RECT 623.950 0.350 628.630 4.280 ;
        RECT 629.470 0.350 634.150 4.280 ;
        RECT 634.990 0.350 639.670 4.280 ;
        RECT 640.510 0.350 645.190 4.280 ;
        RECT 646.030 0.350 650.710 4.280 ;
        RECT 651.550 0.350 656.230 4.280 ;
        RECT 657.070 0.350 661.750 4.280 ;
        RECT 662.590 0.350 667.270 4.280 ;
        RECT 668.110 0.350 672.790 4.280 ;
        RECT 673.630 0.350 678.310 4.280 ;
        RECT 679.150 0.350 683.830 4.280 ;
        RECT 684.670 0.350 689.350 4.280 ;
        RECT 690.190 0.350 694.870 4.280 ;
        RECT 695.710 0.350 700.390 4.280 ;
        RECT 701.230 0.350 705.910 4.280 ;
        RECT 706.750 0.350 711.430 4.280 ;
        RECT 712.270 0.350 716.950 4.280 ;
        RECT 717.790 0.350 722.470 4.280 ;
        RECT 723.310 0.350 727.990 4.280 ;
        RECT 728.830 0.350 733.510 4.280 ;
        RECT 734.350 0.350 739.030 4.280 ;
        RECT 739.870 0.350 744.550 4.280 ;
        RECT 745.390 0.350 750.070 4.280 ;
        RECT 750.910 0.350 755.590 4.280 ;
        RECT 756.430 0.350 761.110 4.280 ;
        RECT 761.950 0.350 766.630 4.280 ;
        RECT 767.470 0.350 772.150 4.280 ;
        RECT 772.990 0.350 777.670 4.280 ;
        RECT 778.510 0.350 783.190 4.280 ;
        RECT 784.030 0.350 788.710 4.280 ;
        RECT 789.550 0.350 794.230 4.280 ;
        RECT 795.070 0.350 799.750 4.280 ;
        RECT 800.590 0.350 805.270 4.280 ;
        RECT 806.110 0.350 810.790 4.280 ;
        RECT 811.630 0.350 816.310 4.280 ;
        RECT 817.150 0.350 821.830 4.280 ;
        RECT 822.670 0.350 827.350 4.280 ;
        RECT 828.190 0.350 832.870 4.280 ;
        RECT 833.710 0.350 838.390 4.280 ;
        RECT 839.230 0.350 843.910 4.280 ;
        RECT 844.750 0.350 849.430 4.280 ;
        RECT 850.270 0.350 854.950 4.280 ;
        RECT 855.790 0.350 860.470 4.280 ;
        RECT 861.310 0.350 865.990 4.280 ;
        RECT 866.830 0.350 871.510 4.280 ;
        RECT 872.350 0.350 877.030 4.280 ;
        RECT 877.870 0.350 882.550 4.280 ;
        RECT 883.390 0.350 888.070 4.280 ;
        RECT 888.910 0.350 893.590 4.280 ;
        RECT 894.430 0.350 899.110 4.280 ;
        RECT 899.950 0.350 904.630 4.280 ;
        RECT 905.470 0.350 910.150 4.280 ;
        RECT 910.990 0.350 915.670 4.280 ;
        RECT 916.510 0.350 921.190 4.280 ;
        RECT 922.030 0.350 926.710 4.280 ;
        RECT 927.550 0.350 932.230 4.280 ;
        RECT 933.070 0.350 937.750 4.280 ;
        RECT 938.590 0.350 943.270 4.280 ;
        RECT 944.110 0.350 948.790 4.280 ;
        RECT 949.630 0.350 954.310 4.280 ;
        RECT 955.150 0.350 959.830 4.280 ;
        RECT 960.670 0.350 965.350 4.280 ;
        RECT 966.190 0.350 970.870 4.280 ;
        RECT 971.710 0.350 976.390 4.280 ;
        RECT 977.230 0.350 981.910 4.280 ;
        RECT 982.750 0.350 987.430 4.280 ;
        RECT 988.270 0.350 992.950 4.280 ;
        RECT 993.790 0.350 998.470 4.280 ;
        RECT 999.310 0.350 1003.990 4.280 ;
        RECT 1004.830 0.350 1009.510 4.280 ;
        RECT 1010.350 0.350 1015.030 4.280 ;
        RECT 1015.870 0.350 1020.550 4.280 ;
        RECT 1021.390 0.350 1026.070 4.280 ;
        RECT 1026.910 0.350 1031.590 4.280 ;
        RECT 1032.430 0.350 1037.110 4.280 ;
        RECT 1037.950 0.350 1042.630 4.280 ;
        RECT 1043.470 0.350 1048.150 4.280 ;
        RECT 1048.990 0.350 1053.670 4.280 ;
        RECT 1054.510 0.350 1059.190 4.280 ;
        RECT 1060.030 0.350 1064.710 4.280 ;
        RECT 1065.550 0.350 1070.230 4.280 ;
        RECT 1071.070 0.350 1075.750 4.280 ;
        RECT 1076.590 0.350 1081.270 4.280 ;
        RECT 1082.110 0.350 1086.790 4.280 ;
        RECT 1087.630 0.350 1092.310 4.280 ;
        RECT 1093.150 0.350 1097.830 4.280 ;
        RECT 1098.670 0.350 1103.350 4.280 ;
        RECT 1104.190 0.350 1108.870 4.280 ;
        RECT 1109.710 0.350 1114.390 4.280 ;
        RECT 1115.230 0.350 1119.910 4.280 ;
        RECT 1120.750 0.350 1125.430 4.280 ;
        RECT 1126.270 0.350 1130.950 4.280 ;
        RECT 1131.790 0.350 1136.470 4.280 ;
        RECT 1137.310 0.350 1141.990 4.280 ;
        RECT 1142.830 0.350 1147.510 4.280 ;
        RECT 1148.350 0.350 1153.030 4.280 ;
        RECT 1153.870 0.350 1158.550 4.280 ;
        RECT 1159.390 0.350 1164.070 4.280 ;
        RECT 1164.910 0.350 1169.590 4.280 ;
        RECT 1170.430 0.350 1175.110 4.280 ;
        RECT 1175.950 0.350 1180.630 4.280 ;
        RECT 1181.470 0.350 1186.150 4.280 ;
        RECT 1186.990 0.350 1191.670 4.280 ;
        RECT 1192.510 0.350 1197.190 4.280 ;
        RECT 1198.030 0.350 1202.710 4.280 ;
        RECT 1203.550 0.350 1208.230 4.280 ;
        RECT 1209.070 0.350 1213.750 4.280 ;
        RECT 1214.590 0.350 1219.270 4.280 ;
        RECT 1220.110 0.350 1224.790 4.280 ;
        RECT 1225.630 0.350 1230.310 4.280 ;
        RECT 1231.150 0.350 1235.830 4.280 ;
        RECT 1236.670 0.350 1241.350 4.280 ;
        RECT 1242.190 0.350 1246.870 4.280 ;
        RECT 1247.710 0.350 1252.390 4.280 ;
        RECT 1253.230 0.350 1257.910 4.280 ;
        RECT 1258.750 0.350 1263.430 4.280 ;
        RECT 1264.270 0.350 1268.950 4.280 ;
        RECT 1269.790 0.350 1274.470 4.280 ;
        RECT 1275.310 0.350 1279.990 4.280 ;
        RECT 1280.830 0.350 1285.510 4.280 ;
        RECT 1286.350 0.350 1291.030 4.280 ;
        RECT 1291.870 0.350 1296.550 4.280 ;
        RECT 1297.390 0.350 1302.070 4.280 ;
        RECT 1302.910 0.350 1307.590 4.280 ;
        RECT 1308.430 0.350 1313.110 4.280 ;
        RECT 1313.950 0.350 1318.630 4.280 ;
        RECT 1319.470 0.350 1324.150 4.280 ;
        RECT 1324.990 0.350 1329.670 4.280 ;
        RECT 1330.510 0.350 1335.190 4.280 ;
        RECT 1336.030 0.350 1340.710 4.280 ;
        RECT 1341.550 0.350 1346.230 4.280 ;
        RECT 1347.070 0.350 1351.750 4.280 ;
        RECT 1352.590 0.350 1357.270 4.280 ;
        RECT 1358.110 0.350 1362.790 4.280 ;
        RECT 1363.630 0.350 1368.310 4.280 ;
        RECT 1369.150 0.350 1373.830 4.280 ;
        RECT 1374.670 0.350 1379.350 4.280 ;
        RECT 1380.190 0.350 1384.870 4.280 ;
        RECT 1385.710 0.350 1390.390 4.280 ;
        RECT 1391.230 0.350 1395.910 4.280 ;
        RECT 1396.750 0.350 1401.430 4.280 ;
        RECT 1402.270 0.350 1406.950 4.280 ;
        RECT 1407.790 0.350 1412.470 4.280 ;
        RECT 1413.310 0.350 1417.990 4.280 ;
        RECT 1418.830 0.350 1423.510 4.280 ;
        RECT 1424.350 0.350 1429.030 4.280 ;
        RECT 1429.870 0.350 1434.550 4.280 ;
        RECT 1435.390 0.350 1440.070 4.280 ;
        RECT 1440.910 0.350 1445.590 4.280 ;
        RECT 1446.430 0.350 1451.110 4.280 ;
        RECT 1451.950 0.350 1456.630 4.280 ;
        RECT 1457.470 0.350 1462.150 4.280 ;
        RECT 1462.990 0.350 1467.670 4.280 ;
        RECT 1468.510 0.350 1473.190 4.280 ;
        RECT 1474.030 0.350 1478.710 4.280 ;
        RECT 1479.550 0.350 1484.230 4.280 ;
        RECT 1485.070 0.350 1489.750 4.280 ;
        RECT 1490.590 0.350 1495.270 4.280 ;
        RECT 1496.110 0.350 1500.790 4.280 ;
        RECT 1501.630 0.350 1506.310 4.280 ;
        RECT 1507.150 0.350 1511.830 4.280 ;
        RECT 1512.670 0.350 1517.350 4.280 ;
        RECT 1518.190 0.350 1522.870 4.280 ;
        RECT 1523.710 0.350 1528.390 4.280 ;
        RECT 1529.230 0.350 1533.910 4.280 ;
        RECT 1534.750 0.350 1539.430 4.280 ;
        RECT 1540.270 0.350 1544.950 4.280 ;
        RECT 1545.790 0.350 1550.470 4.280 ;
        RECT 1551.310 0.350 1555.990 4.280 ;
        RECT 1556.830 0.350 1561.510 4.280 ;
        RECT 1562.350 0.350 1567.030 4.280 ;
        RECT 1567.870 0.350 1572.550 4.280 ;
        RECT 1573.390 0.350 1578.070 4.280 ;
        RECT 1578.910 0.350 1583.590 4.280 ;
        RECT 1584.430 0.350 1589.110 4.280 ;
        RECT 1589.950 0.350 1594.630 4.280 ;
        RECT 1595.470 0.350 1600.150 4.280 ;
        RECT 1600.990 0.350 1605.670 4.280 ;
        RECT 1606.510 0.350 1611.190 4.280 ;
        RECT 1612.030 0.350 1616.710 4.280 ;
        RECT 1617.550 0.350 1622.230 4.280 ;
        RECT 1623.070 0.350 1627.750 4.280 ;
        RECT 1628.590 0.350 1633.270 4.280 ;
        RECT 1634.110 0.350 1638.790 4.280 ;
        RECT 1639.630 0.350 1644.310 4.280 ;
        RECT 1645.150 0.350 1649.830 4.280 ;
        RECT 1650.670 0.350 1655.350 4.280 ;
        RECT 1656.190 0.350 1660.870 4.280 ;
        RECT 1661.710 0.350 1666.390 4.280 ;
        RECT 1667.230 0.350 1671.910 4.280 ;
        RECT 1672.750 0.350 1677.430 4.280 ;
        RECT 1678.270 0.350 1682.950 4.280 ;
        RECT 1683.790 0.350 1688.470 4.280 ;
        RECT 1689.310 0.350 1693.990 4.280 ;
        RECT 1694.830 0.350 1699.510 4.280 ;
        RECT 1700.350 0.350 1705.030 4.280 ;
        RECT 1705.870 0.350 1710.550 4.280 ;
        RECT 1711.390 0.350 1716.070 4.280 ;
        RECT 1716.910 0.350 1721.590 4.280 ;
        RECT 1722.430 0.350 1727.110 4.280 ;
        RECT 1727.950 0.350 1732.630 4.280 ;
        RECT 1733.470 0.350 1738.150 4.280 ;
        RECT 1738.990 0.350 1743.670 4.280 ;
        RECT 1744.510 0.350 1749.190 4.280 ;
        RECT 1750.030 0.350 1754.710 4.280 ;
        RECT 1755.550 0.350 1760.230 4.280 ;
        RECT 1761.070 0.350 1765.750 4.280 ;
        RECT 1766.590 0.350 1771.270 4.280 ;
        RECT 1772.110 0.350 1776.790 4.280 ;
        RECT 1777.630 0.350 1782.310 4.280 ;
        RECT 1783.150 0.350 1787.830 4.280 ;
        RECT 1788.670 0.350 1793.350 4.280 ;
        RECT 1794.190 0.350 1798.870 4.280 ;
        RECT 1799.710 0.350 1804.390 4.280 ;
        RECT 1805.230 0.350 1809.910 4.280 ;
        RECT 1810.750 0.350 1815.430 4.280 ;
        RECT 1816.270 0.350 1820.950 4.280 ;
        RECT 1821.790 0.350 1826.470 4.280 ;
        RECT 1827.310 0.350 1831.990 4.280 ;
        RECT 1832.830 0.350 1837.510 4.280 ;
        RECT 1838.350 0.350 1843.030 4.280 ;
        RECT 1843.870 0.350 1848.550 4.280 ;
        RECT 1849.390 0.350 1854.070 4.280 ;
        RECT 1854.910 0.350 1859.590 4.280 ;
        RECT 1860.430 0.350 1865.110 4.280 ;
        RECT 1865.950 0.350 1870.630 4.280 ;
        RECT 1871.470 0.350 1876.150 4.280 ;
        RECT 1876.990 0.350 1881.670 4.280 ;
        RECT 1882.510 0.350 1887.190 4.280 ;
        RECT 1888.030 0.350 1892.710 4.280 ;
        RECT 1893.550 0.350 1898.230 4.280 ;
        RECT 1899.070 0.350 1903.750 4.280 ;
        RECT 1904.590 0.350 1909.270 4.280 ;
        RECT 1910.110 0.350 1914.790 4.280 ;
        RECT 1915.630 0.350 1920.310 4.280 ;
        RECT 1921.150 0.350 1925.830 4.280 ;
        RECT 1926.670 0.350 1931.350 4.280 ;
        RECT 1932.190 0.350 1936.870 4.280 ;
        RECT 1937.710 0.350 1942.390 4.280 ;
        RECT 1943.230 0.350 1947.910 4.280 ;
        RECT 1948.750 0.350 1953.430 4.280 ;
        RECT 1954.270 0.350 1958.950 4.280 ;
        RECT 1959.790 0.350 1964.470 4.280 ;
        RECT 1965.310 0.350 1969.990 4.280 ;
        RECT 1970.830 0.350 1975.510 4.280 ;
        RECT 1976.350 0.350 1981.030 4.280 ;
        RECT 1981.870 0.350 1986.550 4.280 ;
        RECT 1987.390 0.350 1992.070 4.280 ;
        RECT 1992.910 0.350 1997.590 4.280 ;
        RECT 1998.430 0.350 2003.110 4.280 ;
        RECT 2003.950 0.350 2008.630 4.280 ;
        RECT 2009.470 0.350 2014.150 4.280 ;
        RECT 2014.990 0.350 2019.670 4.280 ;
        RECT 2020.510 0.350 2025.190 4.280 ;
        RECT 2026.030 0.350 2030.710 4.280 ;
        RECT 2031.550 0.350 2036.230 4.280 ;
        RECT 2037.070 0.350 2041.750 4.280 ;
        RECT 2042.590 0.350 2047.270 4.280 ;
        RECT 2048.110 0.350 2052.790 4.280 ;
        RECT 2053.630 0.350 2058.310 4.280 ;
        RECT 2059.150 0.350 2063.830 4.280 ;
        RECT 2064.670 0.350 2069.350 4.280 ;
        RECT 2070.190 0.350 2074.870 4.280 ;
        RECT 2075.710 0.350 2080.390 4.280 ;
        RECT 2081.230 0.350 2085.910 4.280 ;
        RECT 2086.750 0.350 2091.430 4.280 ;
        RECT 2092.270 0.350 2096.950 4.280 ;
        RECT 2097.790 0.350 2102.470 4.280 ;
        RECT 2103.310 0.350 2107.990 4.280 ;
        RECT 2108.830 0.350 2113.510 4.280 ;
        RECT 2114.350 0.350 2119.030 4.280 ;
        RECT 2119.870 0.350 2124.550 4.280 ;
        RECT 2125.390 0.350 2130.070 4.280 ;
        RECT 2130.910 0.350 2135.590 4.280 ;
        RECT 2136.430 0.350 2141.110 4.280 ;
        RECT 2141.950 0.350 2146.630 4.280 ;
        RECT 2147.470 0.350 2152.150 4.280 ;
        RECT 2152.990 0.350 2157.670 4.280 ;
        RECT 2158.510 0.350 2163.190 4.280 ;
        RECT 2164.030 0.350 2168.710 4.280 ;
        RECT 2169.550 0.350 2174.230 4.280 ;
        RECT 2175.070 0.350 2179.750 4.280 ;
        RECT 2180.590 0.350 2185.270 4.280 ;
        RECT 2186.110 0.350 2190.790 4.280 ;
        RECT 2191.630 0.350 2196.310 4.280 ;
        RECT 2197.150 0.350 2201.830 4.280 ;
        RECT 2202.670 0.350 2207.350 4.280 ;
        RECT 2208.190 0.350 2212.870 4.280 ;
        RECT 2213.710 0.350 2218.390 4.280 ;
        RECT 2219.230 0.350 2223.910 4.280 ;
        RECT 2224.750 0.350 2229.430 4.280 ;
        RECT 2230.270 0.350 2234.950 4.280 ;
        RECT 2235.790 0.350 2240.470 4.280 ;
        RECT 2241.310 0.350 2245.990 4.280 ;
        RECT 2246.830 0.350 2251.510 4.280 ;
        RECT 2252.350 0.350 2257.030 4.280 ;
        RECT 2257.870 0.350 2262.550 4.280 ;
        RECT 2263.390 0.350 2268.070 4.280 ;
        RECT 2268.910 0.350 2273.590 4.280 ;
        RECT 2274.430 0.350 2279.110 4.280 ;
        RECT 2279.950 0.350 2284.630 4.280 ;
        RECT 2285.470 0.350 2290.150 4.280 ;
        RECT 2290.990 0.350 2295.670 4.280 ;
        RECT 2296.510 0.350 2301.190 4.280 ;
        RECT 2302.030 0.350 2306.710 4.280 ;
        RECT 2307.550 0.350 2312.230 4.280 ;
        RECT 2313.070 0.350 2317.750 4.280 ;
        RECT 2318.590 0.350 2323.270 4.280 ;
        RECT 2324.110 0.350 2328.790 4.280 ;
        RECT 2329.630 0.350 2334.310 4.280 ;
        RECT 2335.150 0.350 2339.830 4.280 ;
        RECT 2340.670 0.350 2345.350 4.280 ;
        RECT 2346.190 0.350 2350.870 4.280 ;
        RECT 2351.710 0.350 2356.390 4.280 ;
        RECT 2357.230 0.350 2361.910 4.280 ;
        RECT 2362.750 0.350 2367.430 4.280 ;
        RECT 2368.270 0.350 2372.950 4.280 ;
        RECT 2373.790 0.350 2378.470 4.280 ;
        RECT 2379.310 0.350 2383.990 4.280 ;
        RECT 2384.830 0.350 2389.510 4.280 ;
        RECT 2390.350 0.350 2395.030 4.280 ;
        RECT 2395.870 0.350 2400.550 4.280 ;
        RECT 2401.390 0.350 2406.070 4.280 ;
        RECT 2406.910 0.350 2411.590 4.280 ;
        RECT 2412.430 0.350 2417.110 4.280 ;
        RECT 2417.950 0.350 2422.630 4.280 ;
        RECT 2423.470 0.350 2428.150 4.280 ;
        RECT 2428.990 0.350 2433.670 4.280 ;
        RECT 2434.510 0.350 2439.190 4.280 ;
        RECT 2440.030 0.350 2444.710 4.280 ;
        RECT 2445.550 0.350 2450.230 4.280 ;
        RECT 2451.070 0.350 2455.750 4.280 ;
        RECT 2456.590 0.350 2461.270 4.280 ;
        RECT 2462.110 0.350 2466.790 4.280 ;
        RECT 2467.630 0.350 2472.310 4.280 ;
        RECT 2473.150 0.350 2477.830 4.280 ;
        RECT 2478.670 0.350 2483.350 4.280 ;
        RECT 2484.190 0.350 2488.870 4.280 ;
        RECT 2489.710 0.350 2494.390 4.280 ;
        RECT 2495.230 0.350 2499.910 4.280 ;
        RECT 2500.750 0.350 2505.430 4.280 ;
        RECT 2506.270 0.350 2510.950 4.280 ;
        RECT 2511.790 0.350 2516.470 4.280 ;
        RECT 2517.310 0.350 2521.990 4.280 ;
        RECT 2522.830 0.350 2527.510 4.280 ;
        RECT 2528.350 0.350 2533.030 4.280 ;
        RECT 2533.870 0.350 2538.550 4.280 ;
        RECT 2539.390 0.350 2544.070 4.280 ;
        RECT 2544.910 0.350 2549.590 4.280 ;
        RECT 2550.430 0.350 2555.110 4.280 ;
        RECT 2555.950 0.350 2560.630 4.280 ;
        RECT 2561.470 0.350 2566.150 4.280 ;
        RECT 2566.990 0.350 2571.670 4.280 ;
        RECT 2572.510 0.350 2577.190 4.280 ;
        RECT 2578.030 0.350 2582.710 4.280 ;
        RECT 2583.550 0.350 2588.230 4.280 ;
        RECT 2589.070 0.350 2593.750 4.280 ;
        RECT 2594.590 0.350 2599.270 4.280 ;
        RECT 2600.110 0.350 2604.790 4.280 ;
        RECT 2605.630 0.350 2610.310 4.280 ;
        RECT 2611.150 0.350 2615.830 4.280 ;
        RECT 2616.670 0.350 2621.350 4.280 ;
        RECT 2622.190 0.350 2626.870 4.280 ;
        RECT 2627.710 0.350 2632.390 4.280 ;
        RECT 2633.230 0.350 2637.910 4.280 ;
        RECT 2638.750 0.350 2643.430 4.280 ;
        RECT 2644.270 0.350 2648.950 4.280 ;
        RECT 2649.790 0.350 2654.470 4.280 ;
        RECT 2655.310 0.350 2659.990 4.280 ;
        RECT 2660.830 0.350 2665.510 4.280 ;
        RECT 2666.350 0.350 2671.030 4.280 ;
        RECT 2671.870 0.350 2676.550 4.280 ;
        RECT 2677.390 0.350 2682.070 4.280 ;
        RECT 2682.910 0.350 2687.590 4.280 ;
        RECT 2688.430 0.350 2693.110 4.280 ;
        RECT 2693.950 0.350 2698.630 4.280 ;
        RECT 2699.470 0.350 2704.150 4.280 ;
        RECT 2704.990 0.350 2709.670 4.280 ;
        RECT 2710.510 0.350 2715.190 4.280 ;
        RECT 2716.030 0.350 2720.710 4.280 ;
        RECT 2721.550 0.350 2726.230 4.280 ;
        RECT 2727.070 0.350 2731.750 4.280 ;
        RECT 2732.590 0.350 2737.270 4.280 ;
        RECT 2738.110 0.350 2742.790 4.280 ;
        RECT 2743.630 0.350 2748.310 4.280 ;
        RECT 2749.150 0.350 2753.830 4.280 ;
        RECT 2754.670 0.350 2759.350 4.280 ;
        RECT 2760.190 0.350 2764.870 4.280 ;
        RECT 2765.710 0.350 2770.390 4.280 ;
        RECT 2771.230 0.350 2775.910 4.280 ;
        RECT 2776.750 0.350 2781.430 4.280 ;
        RECT 2782.270 0.350 2786.950 4.280 ;
        RECT 2787.790 0.350 2792.470 4.280 ;
        RECT 2793.310 0.350 2797.990 4.280 ;
        RECT 2798.830 0.350 2803.510 4.280 ;
        RECT 2804.350 0.350 2809.030 4.280 ;
        RECT 2809.870 0.350 2814.550 4.280 ;
        RECT 2815.390 0.350 2820.070 4.280 ;
        RECT 2820.910 0.350 2917.220 4.280 ;
      LAYER met3 ;
        RECT 2.150 3456.800 2916.000 3508.965 ;
        RECT 2.150 3455.400 2915.600 3456.800 ;
        RECT 2.150 3454.080 2916.000 3455.400 ;
        RECT 4.400 3452.680 2916.000 3454.080 ;
        RECT 2.150 3391.520 2916.000 3452.680 ;
        RECT 2.150 3390.160 2915.600 3391.520 ;
        RECT 4.400 3390.120 2915.600 3390.160 ;
        RECT 4.400 3388.760 2916.000 3390.120 ;
        RECT 2.150 3326.240 2916.000 3388.760 ;
        RECT 4.400 3324.840 2915.600 3326.240 ;
        RECT 2.150 3262.320 2916.000 3324.840 ;
        RECT 4.400 3260.960 2916.000 3262.320 ;
        RECT 4.400 3260.920 2915.600 3260.960 ;
        RECT 2.150 3259.560 2915.600 3260.920 ;
        RECT 2.150 3198.400 2916.000 3259.560 ;
        RECT 4.400 3197.000 2916.000 3198.400 ;
        RECT 2.150 3195.680 2916.000 3197.000 ;
        RECT 2.150 3194.280 2915.600 3195.680 ;
        RECT 2.150 3134.480 2916.000 3194.280 ;
        RECT 4.400 3133.080 2916.000 3134.480 ;
        RECT 2.150 3130.400 2916.000 3133.080 ;
        RECT 2.150 3129.000 2915.600 3130.400 ;
        RECT 2.150 3070.560 2916.000 3129.000 ;
        RECT 4.400 3069.160 2916.000 3070.560 ;
        RECT 2.150 3065.120 2916.000 3069.160 ;
        RECT 2.150 3063.720 2915.600 3065.120 ;
        RECT 2.150 3006.640 2916.000 3063.720 ;
        RECT 4.400 3005.240 2916.000 3006.640 ;
        RECT 2.150 2999.840 2916.000 3005.240 ;
        RECT 2.150 2998.440 2915.600 2999.840 ;
        RECT 2.150 2942.720 2916.000 2998.440 ;
        RECT 4.400 2941.320 2916.000 2942.720 ;
        RECT 2.150 2934.560 2916.000 2941.320 ;
        RECT 2.150 2933.160 2915.600 2934.560 ;
        RECT 2.150 2878.800 2916.000 2933.160 ;
        RECT 4.400 2877.400 2916.000 2878.800 ;
        RECT 2.150 2869.280 2916.000 2877.400 ;
        RECT 2.150 2867.880 2915.600 2869.280 ;
        RECT 2.150 2814.880 2916.000 2867.880 ;
        RECT 4.400 2813.480 2916.000 2814.880 ;
        RECT 2.150 2804.000 2916.000 2813.480 ;
        RECT 2.150 2802.600 2915.600 2804.000 ;
        RECT 2.150 2750.960 2916.000 2802.600 ;
        RECT 4.400 2749.560 2916.000 2750.960 ;
        RECT 2.150 2738.720 2916.000 2749.560 ;
        RECT 2.150 2737.320 2915.600 2738.720 ;
        RECT 2.150 2687.040 2916.000 2737.320 ;
        RECT 4.400 2685.640 2916.000 2687.040 ;
        RECT 2.150 2673.440 2916.000 2685.640 ;
        RECT 2.150 2672.040 2915.600 2673.440 ;
        RECT 2.150 2623.120 2916.000 2672.040 ;
        RECT 4.400 2621.720 2916.000 2623.120 ;
        RECT 2.150 2608.160 2916.000 2621.720 ;
        RECT 2.150 2606.760 2915.600 2608.160 ;
        RECT 2.150 2559.200 2916.000 2606.760 ;
        RECT 4.400 2557.800 2916.000 2559.200 ;
        RECT 2.150 2542.880 2916.000 2557.800 ;
        RECT 2.150 2541.480 2915.600 2542.880 ;
        RECT 2.150 2495.280 2916.000 2541.480 ;
        RECT 4.400 2493.880 2916.000 2495.280 ;
        RECT 2.150 2477.600 2916.000 2493.880 ;
        RECT 2.150 2476.200 2915.600 2477.600 ;
        RECT 2.150 2431.360 2916.000 2476.200 ;
        RECT 4.400 2429.960 2916.000 2431.360 ;
        RECT 2.150 2412.320 2916.000 2429.960 ;
        RECT 2.150 2410.920 2915.600 2412.320 ;
        RECT 2.150 2367.440 2916.000 2410.920 ;
        RECT 4.400 2366.040 2916.000 2367.440 ;
        RECT 2.150 2347.040 2916.000 2366.040 ;
        RECT 2.150 2345.640 2915.600 2347.040 ;
        RECT 2.150 2303.520 2916.000 2345.640 ;
        RECT 4.400 2302.120 2916.000 2303.520 ;
        RECT 2.150 2281.760 2916.000 2302.120 ;
        RECT 2.150 2280.360 2915.600 2281.760 ;
        RECT 2.150 2239.600 2916.000 2280.360 ;
        RECT 4.400 2238.200 2916.000 2239.600 ;
        RECT 2.150 2216.480 2916.000 2238.200 ;
        RECT 2.150 2215.080 2915.600 2216.480 ;
        RECT 2.150 2175.680 2916.000 2215.080 ;
        RECT 4.400 2174.280 2916.000 2175.680 ;
        RECT 2.150 2151.200 2916.000 2174.280 ;
        RECT 2.150 2149.800 2915.600 2151.200 ;
        RECT 2.150 2111.760 2916.000 2149.800 ;
        RECT 4.400 2110.360 2916.000 2111.760 ;
        RECT 2.150 2085.920 2916.000 2110.360 ;
        RECT 2.150 2084.520 2915.600 2085.920 ;
        RECT 2.150 2047.840 2916.000 2084.520 ;
        RECT 4.400 2046.440 2916.000 2047.840 ;
        RECT 2.150 2020.640 2916.000 2046.440 ;
        RECT 2.150 2019.240 2915.600 2020.640 ;
        RECT 2.150 1983.920 2916.000 2019.240 ;
        RECT 4.400 1982.520 2916.000 1983.920 ;
        RECT 2.150 1955.360 2916.000 1982.520 ;
        RECT 2.150 1953.960 2915.600 1955.360 ;
        RECT 2.150 1920.000 2916.000 1953.960 ;
        RECT 4.400 1918.600 2916.000 1920.000 ;
        RECT 2.150 1890.080 2916.000 1918.600 ;
        RECT 2.150 1888.680 2915.600 1890.080 ;
        RECT 2.150 1856.080 2916.000 1888.680 ;
        RECT 4.400 1854.680 2916.000 1856.080 ;
        RECT 2.150 1824.800 2916.000 1854.680 ;
        RECT 2.150 1823.400 2915.600 1824.800 ;
        RECT 2.150 1792.160 2916.000 1823.400 ;
        RECT 4.400 1790.760 2916.000 1792.160 ;
        RECT 2.150 1759.520 2916.000 1790.760 ;
        RECT 2.150 1758.120 2915.600 1759.520 ;
        RECT 2.150 1728.240 2916.000 1758.120 ;
        RECT 4.400 1726.840 2916.000 1728.240 ;
        RECT 2.150 1694.240 2916.000 1726.840 ;
        RECT 2.150 1692.840 2915.600 1694.240 ;
        RECT 2.150 1664.320 2916.000 1692.840 ;
        RECT 4.400 1662.920 2916.000 1664.320 ;
        RECT 2.150 1628.960 2916.000 1662.920 ;
        RECT 2.150 1627.560 2915.600 1628.960 ;
        RECT 2.150 1600.400 2916.000 1627.560 ;
        RECT 4.400 1599.000 2916.000 1600.400 ;
        RECT 2.150 1563.680 2916.000 1599.000 ;
        RECT 2.150 1562.280 2915.600 1563.680 ;
        RECT 2.150 1536.480 2916.000 1562.280 ;
        RECT 4.400 1535.080 2916.000 1536.480 ;
        RECT 2.150 1498.400 2916.000 1535.080 ;
        RECT 2.150 1497.000 2915.600 1498.400 ;
        RECT 2.150 1472.560 2916.000 1497.000 ;
        RECT 4.400 1471.160 2916.000 1472.560 ;
        RECT 2.150 1433.120 2916.000 1471.160 ;
        RECT 2.150 1431.720 2915.600 1433.120 ;
        RECT 2.150 1408.640 2916.000 1431.720 ;
        RECT 4.400 1407.240 2916.000 1408.640 ;
        RECT 2.150 1367.840 2916.000 1407.240 ;
        RECT 2.150 1366.440 2915.600 1367.840 ;
        RECT 2.150 1344.720 2916.000 1366.440 ;
        RECT 4.400 1343.320 2916.000 1344.720 ;
        RECT 2.150 1302.560 2916.000 1343.320 ;
        RECT 2.150 1301.160 2915.600 1302.560 ;
        RECT 2.150 1280.800 2916.000 1301.160 ;
        RECT 4.400 1279.400 2916.000 1280.800 ;
        RECT 2.150 1237.280 2916.000 1279.400 ;
        RECT 2.150 1235.880 2915.600 1237.280 ;
        RECT 2.150 1216.880 2916.000 1235.880 ;
        RECT 4.400 1215.480 2916.000 1216.880 ;
        RECT 2.150 1172.000 2916.000 1215.480 ;
        RECT 2.150 1170.600 2915.600 1172.000 ;
        RECT 2.150 1152.960 2916.000 1170.600 ;
        RECT 4.400 1151.560 2916.000 1152.960 ;
        RECT 2.150 1106.720 2916.000 1151.560 ;
        RECT 2.150 1105.320 2915.600 1106.720 ;
        RECT 2.150 1089.040 2916.000 1105.320 ;
        RECT 4.400 1087.640 2916.000 1089.040 ;
        RECT 2.150 1041.440 2916.000 1087.640 ;
        RECT 2.150 1040.040 2915.600 1041.440 ;
        RECT 2.150 1025.120 2916.000 1040.040 ;
        RECT 4.400 1023.720 2916.000 1025.120 ;
        RECT 2.150 976.160 2916.000 1023.720 ;
        RECT 2.150 974.760 2915.600 976.160 ;
        RECT 2.150 961.200 2916.000 974.760 ;
        RECT 4.400 959.800 2916.000 961.200 ;
        RECT 2.150 910.880 2916.000 959.800 ;
        RECT 2.150 909.480 2915.600 910.880 ;
        RECT 2.150 897.280 2916.000 909.480 ;
        RECT 4.400 895.880 2916.000 897.280 ;
        RECT 2.150 845.600 2916.000 895.880 ;
        RECT 2.150 844.200 2915.600 845.600 ;
        RECT 2.150 833.360 2916.000 844.200 ;
        RECT 4.400 831.960 2916.000 833.360 ;
        RECT 2.150 780.320 2916.000 831.960 ;
        RECT 2.150 778.920 2915.600 780.320 ;
        RECT 2.150 769.440 2916.000 778.920 ;
        RECT 4.400 768.040 2916.000 769.440 ;
        RECT 2.150 715.040 2916.000 768.040 ;
        RECT 2.150 713.640 2915.600 715.040 ;
        RECT 2.150 705.520 2916.000 713.640 ;
        RECT 4.400 704.120 2916.000 705.520 ;
        RECT 2.150 649.760 2916.000 704.120 ;
        RECT 2.150 648.360 2915.600 649.760 ;
        RECT 2.150 641.600 2916.000 648.360 ;
        RECT 4.400 640.200 2916.000 641.600 ;
        RECT 2.150 584.480 2916.000 640.200 ;
        RECT 2.150 583.080 2915.600 584.480 ;
        RECT 2.150 577.680 2916.000 583.080 ;
        RECT 4.400 576.280 2916.000 577.680 ;
        RECT 2.150 519.200 2916.000 576.280 ;
        RECT 2.150 517.800 2915.600 519.200 ;
        RECT 2.150 513.760 2916.000 517.800 ;
        RECT 4.400 512.360 2916.000 513.760 ;
        RECT 2.150 453.920 2916.000 512.360 ;
        RECT 2.150 452.520 2915.600 453.920 ;
        RECT 2.150 449.840 2916.000 452.520 ;
        RECT 4.400 448.440 2916.000 449.840 ;
        RECT 2.150 388.640 2916.000 448.440 ;
        RECT 2.150 387.240 2915.600 388.640 ;
        RECT 2.150 385.920 2916.000 387.240 ;
        RECT 4.400 384.520 2916.000 385.920 ;
        RECT 2.150 323.360 2916.000 384.520 ;
        RECT 2.150 322.000 2915.600 323.360 ;
        RECT 4.400 321.960 2915.600 322.000 ;
        RECT 4.400 320.600 2916.000 321.960 ;
        RECT 2.150 258.080 2916.000 320.600 ;
        RECT 4.400 256.680 2915.600 258.080 ;
        RECT 2.150 194.160 2916.000 256.680 ;
        RECT 4.400 192.800 2916.000 194.160 ;
        RECT 4.400 192.760 2915.600 192.800 ;
        RECT 2.150 191.400 2915.600 192.760 ;
        RECT 2.150 130.240 2916.000 191.400 ;
        RECT 4.400 128.840 2916.000 130.240 ;
        RECT 2.150 127.520 2916.000 128.840 ;
        RECT 2.150 126.120 2915.600 127.520 ;
        RECT 2.150 66.320 2916.000 126.120 ;
        RECT 4.400 64.920 2916.000 66.320 ;
        RECT 2.150 62.240 2916.000 64.920 ;
        RECT 2.150 60.840 2915.600 62.240 ;
        RECT 2.150 7.655 2916.000 60.840 ;
      LAYER met4 ;
        RECT 7.655 19.215 8.320 3507.945 ;
        RECT 12.120 2619.080 53.620 3507.945 ;
        RECT 57.420 2619.080 58.320 3507.945 ;
        RECT 62.120 2619.080 103.620 3507.945 ;
        RECT 107.420 2619.080 108.320 3507.945 ;
        RECT 112.120 2619.080 153.620 3507.945 ;
        RECT 157.420 2619.080 158.320 3507.945 ;
        RECT 162.120 2619.080 203.620 3507.945 ;
        RECT 207.420 2619.700 208.320 3507.945 ;
        RECT 212.120 2619.700 253.620 3507.945 ;
        RECT 257.420 2619.700 258.320 3507.945 ;
        RECT 262.120 2619.700 303.620 3507.945 ;
        RECT 207.420 2619.080 303.620 2619.700 ;
        RECT 307.420 2619.700 308.320 3507.945 ;
        RECT 312.120 2619.700 353.620 3507.945 ;
        RECT 357.420 2619.700 358.320 3507.945 ;
        RECT 362.120 2619.700 403.620 3507.945 ;
        RECT 307.420 2619.080 403.620 2619.700 ;
        RECT 407.420 2619.080 408.320 3507.945 ;
        RECT 412.120 2619.080 453.620 3507.945 ;
        RECT 457.420 2619.080 458.320 3507.945 ;
        RECT 462.120 2619.080 503.620 3507.945 ;
        RECT 507.420 2619.080 508.320 3507.945 ;
        RECT 512.120 2619.080 553.620 3507.945 ;
        RECT 12.120 2202.420 553.620 2619.080 ;
        RECT 12.120 19.215 53.620 2202.420 ;
        RECT 57.420 19.215 58.320 2202.420 ;
        RECT 62.120 19.215 103.620 2202.420 ;
        RECT 107.420 19.215 108.320 2202.420 ;
        RECT 112.120 2201.800 158.320 2202.420 ;
        RECT 112.120 1938.040 153.620 2201.800 ;
        RECT 157.420 1938.040 158.320 2201.800 ;
        RECT 112.120 1930.825 158.320 1938.040 ;
        RECT 162.120 2201.800 353.620 2202.420 ;
        RECT 162.120 1930.825 203.620 2201.800 ;
        RECT 112.120 408.815 203.620 1930.825 ;
        RECT 112.120 405.000 158.320 408.815 ;
        RECT 112.120 19.215 153.620 405.000 ;
        RECT 157.420 19.215 158.320 405.000 ;
        RECT 162.120 19.215 203.620 408.815 ;
        RECT 207.420 1939.665 208.320 2201.800 ;
        RECT 212.120 1939.665 253.620 2201.800 ;
        RECT 257.420 1939.665 258.320 2201.800 ;
        RECT 262.120 1995.520 303.620 2201.800 ;
        RECT 307.420 1995.520 308.320 2201.800 ;
        RECT 262.120 1978.785 308.320 1995.520 ;
        RECT 312.120 1978.785 353.620 2201.800 ;
        RECT 357.420 2201.800 403.620 2202.420 ;
        RECT 357.420 1995.520 358.320 2201.800 ;
        RECT 362.120 1995.520 403.620 2201.800 ;
        RECT 357.420 1978.785 403.620 1995.520 ;
        RECT 262.120 1939.665 403.620 1978.785 ;
        RECT 407.420 1939.665 408.320 2202.420 ;
        RECT 412.120 1939.665 453.620 2202.420 ;
        RECT 207.420 401.335 453.620 1939.665 ;
        RECT 207.420 19.215 208.320 401.335 ;
        RECT 212.120 19.215 253.620 401.335 ;
        RECT 257.420 19.215 258.320 401.335 ;
        RECT 262.120 345.440 308.320 401.335 ;
        RECT 262.120 19.215 303.620 345.440 ;
        RECT 307.420 19.215 308.320 345.440 ;
        RECT 312.120 19.215 353.620 401.335 ;
        RECT 357.420 354.015 453.620 401.335 ;
        RECT 357.420 345.440 403.620 354.015 ;
        RECT 357.420 19.215 358.320 345.440 ;
        RECT 362.120 19.215 403.620 345.440 ;
        RECT 407.420 19.215 408.320 354.015 ;
        RECT 412.120 19.215 453.620 354.015 ;
        RECT 457.420 1939.665 458.320 2202.420 ;
        RECT 462.120 1939.665 503.620 2202.420 ;
        RECT 507.420 1939.665 508.320 2202.420 ;
        RECT 512.120 1995.520 553.620 2202.420 ;
        RECT 557.420 1995.520 558.320 3507.945 ;
        RECT 512.120 1978.785 558.320 1995.520 ;
        RECT 562.120 1978.785 603.620 3507.945 ;
        RECT 607.420 1995.520 608.320 3507.945 ;
        RECT 612.120 1995.520 653.620 3507.945 ;
        RECT 607.420 1978.785 653.620 1995.520 ;
        RECT 512.120 1939.665 653.620 1978.785 ;
        RECT 657.420 1939.665 658.320 3507.945 ;
        RECT 662.120 1939.665 703.620 3507.945 ;
        RECT 457.420 401.335 703.620 1939.665 ;
        RECT 457.420 19.215 458.320 401.335 ;
        RECT 462.120 19.215 503.620 401.335 ;
        RECT 507.420 19.215 508.320 401.335 ;
        RECT 512.120 345.440 558.320 401.335 ;
        RECT 512.120 19.215 553.620 345.440 ;
        RECT 557.420 19.215 558.320 345.440 ;
        RECT 562.120 19.215 603.620 401.335 ;
        RECT 607.420 354.015 703.620 401.335 ;
        RECT 607.420 345.440 653.620 354.015 ;
        RECT 607.420 19.215 608.320 345.440 ;
        RECT 612.120 19.215 653.620 345.440 ;
        RECT 657.420 19.215 658.320 354.015 ;
        RECT 662.120 19.215 703.620 354.015 ;
        RECT 707.420 1939.665 708.320 3507.945 ;
        RECT 712.120 1939.665 753.620 3507.945 ;
        RECT 757.420 1939.665 758.320 3507.945 ;
        RECT 762.120 1995.520 803.620 3507.945 ;
        RECT 807.420 1995.520 808.320 3507.945 ;
        RECT 762.120 1978.785 808.320 1995.520 ;
        RECT 812.120 1978.785 853.620 3507.945 ;
        RECT 857.420 1995.520 858.320 3507.945 ;
        RECT 862.120 1995.520 903.620 3507.945 ;
        RECT 857.420 1978.785 903.620 1995.520 ;
        RECT 762.120 1939.665 903.620 1978.785 ;
        RECT 907.420 1939.665 908.320 3507.945 ;
        RECT 912.120 1939.665 953.620 3507.945 ;
        RECT 957.420 1939.665 958.320 3507.945 ;
        RECT 962.120 1995.520 1003.620 3507.945 ;
        RECT 1007.420 1995.520 1008.320 3507.945 ;
        RECT 962.120 1939.665 1008.320 1995.520 ;
        RECT 1012.120 1978.785 1053.620 3507.945 ;
        RECT 1057.420 1995.520 1058.320 3507.945 ;
        RECT 1062.120 1995.520 1103.620 3507.945 ;
        RECT 1057.420 1978.785 1103.620 1995.520 ;
        RECT 1107.420 1978.785 1108.320 3507.945 ;
        RECT 1112.120 1978.785 1153.620 3507.945 ;
        RECT 1012.120 1939.665 1153.620 1978.785 ;
        RECT 1157.420 1939.665 1158.320 3507.945 ;
        RECT 1162.120 1939.665 1203.620 3507.945 ;
        RECT 1207.420 1939.665 1208.320 3507.945 ;
        RECT 1212.120 1939.665 1253.620 3507.945 ;
        RECT 1257.420 1939.665 1258.320 3507.945 ;
        RECT 1262.120 1995.520 1303.620 3507.945 ;
        RECT 1307.420 1995.520 1308.320 3507.945 ;
        RECT 1262.120 1978.785 1308.320 1995.520 ;
        RECT 1312.120 1995.520 1353.620 3507.945 ;
        RECT 1357.420 1995.520 1358.320 3507.945 ;
        RECT 1362.120 1995.520 1403.620 3507.945 ;
        RECT 1312.120 1978.785 1403.620 1995.520 ;
        RECT 1262.120 1939.665 1403.620 1978.785 ;
        RECT 1407.420 1995.520 1408.320 3507.945 ;
        RECT 1412.120 1995.520 1453.620 3507.945 ;
        RECT 1407.420 1939.665 1453.620 1995.520 ;
        RECT 1457.420 1939.665 1458.320 3507.945 ;
        RECT 1462.120 1939.665 1503.620 3507.945 ;
        RECT 1507.420 1939.665 1508.320 3507.945 ;
        RECT 1512.120 1978.785 1553.620 3507.945 ;
        RECT 1557.420 1978.785 1558.320 3507.945 ;
        RECT 1562.120 1978.785 1603.620 3507.945 ;
        RECT 1512.120 1939.665 1603.620 1978.785 ;
        RECT 1607.420 1939.665 1608.320 3507.945 ;
        RECT 1612.120 1995.520 1653.620 3507.945 ;
        RECT 1657.420 1995.520 1658.320 3507.945 ;
        RECT 1612.120 1939.665 1658.320 1995.520 ;
        RECT 1662.120 1995.520 1703.620 3507.945 ;
        RECT 1707.420 1995.520 1708.320 3507.945 ;
        RECT 1662.120 1939.665 1708.320 1995.520 ;
        RECT 1712.120 1978.785 1753.620 3507.945 ;
        RECT 1757.420 1995.520 1758.320 3507.945 ;
        RECT 1762.120 1995.520 1803.620 3507.945 ;
        RECT 1757.420 1978.785 1803.620 1995.520 ;
        RECT 1807.420 1978.785 1808.320 3507.945 ;
        RECT 1812.120 1978.785 1853.620 3507.945 ;
        RECT 1712.120 1939.665 1853.620 1978.785 ;
        RECT 1857.420 1939.665 1858.320 3507.945 ;
        RECT 1862.120 1939.665 1903.620 3507.945 ;
        RECT 1907.420 1939.665 1908.320 3507.945 ;
        RECT 707.420 401.335 1908.320 1939.665 ;
        RECT 707.420 19.215 708.320 401.335 ;
        RECT 712.120 19.215 753.620 401.335 ;
        RECT 757.420 19.215 758.320 401.335 ;
        RECT 762.120 345.440 808.320 401.335 ;
        RECT 762.120 19.215 803.620 345.440 ;
        RECT 807.420 19.215 808.320 345.440 ;
        RECT 812.120 19.215 853.620 401.335 ;
        RECT 857.420 354.015 953.620 401.335 ;
        RECT 857.420 345.440 903.620 354.015 ;
        RECT 857.420 19.215 858.320 345.440 ;
        RECT 862.120 19.215 903.620 345.440 ;
        RECT 907.420 19.215 908.320 354.015 ;
        RECT 912.120 19.215 953.620 354.015 ;
        RECT 957.420 19.215 958.320 401.335 ;
        RECT 962.120 345.440 1008.320 401.335 ;
        RECT 962.120 19.215 1003.620 345.440 ;
        RECT 1007.420 19.215 1008.320 345.440 ;
        RECT 1012.120 19.215 1053.620 401.335 ;
        RECT 1057.420 345.440 1103.620 401.335 ;
        RECT 1057.420 19.215 1058.320 345.440 ;
        RECT 1062.120 19.215 1103.620 345.440 ;
        RECT 1107.420 19.215 1108.320 401.335 ;
        RECT 1112.120 19.215 1153.620 401.335 ;
        RECT 1157.420 19.215 1158.320 401.335 ;
        RECT 1162.120 19.215 1203.620 401.335 ;
        RECT 1207.420 19.215 1208.320 401.335 ;
        RECT 1212.120 19.215 1253.620 401.335 ;
        RECT 1257.420 19.215 1258.320 401.335 ;
        RECT 1262.120 345.440 1308.320 401.335 ;
        RECT 1262.120 19.215 1303.620 345.440 ;
        RECT 1307.420 19.215 1308.320 345.440 ;
        RECT 1312.120 345.440 1403.620 401.335 ;
        RECT 1312.120 19.215 1353.620 345.440 ;
        RECT 1357.420 19.215 1358.320 345.440 ;
        RECT 1362.120 19.215 1403.620 345.440 ;
        RECT 1407.420 345.440 1453.620 401.335 ;
        RECT 1407.420 19.215 1408.320 345.440 ;
        RECT 1412.120 19.215 1453.620 345.440 ;
        RECT 1457.420 19.215 1458.320 401.335 ;
        RECT 1462.120 19.215 1503.620 401.335 ;
        RECT 1507.420 19.215 1508.320 401.335 ;
        RECT 1512.120 19.215 1553.620 401.335 ;
        RECT 1557.420 19.215 1558.320 401.335 ;
        RECT 1562.120 354.015 1658.320 401.335 ;
        RECT 1562.120 19.215 1603.620 354.015 ;
        RECT 1607.420 19.215 1608.320 354.015 ;
        RECT 1612.120 345.440 1658.320 354.015 ;
        RECT 1612.120 19.215 1653.620 345.440 ;
        RECT 1657.420 19.215 1658.320 345.440 ;
        RECT 1662.120 345.440 1708.320 401.335 ;
        RECT 1662.120 19.215 1703.620 345.440 ;
        RECT 1707.420 19.215 1708.320 345.440 ;
        RECT 1712.120 19.215 1753.620 401.335 ;
        RECT 1757.420 345.440 1803.620 401.335 ;
        RECT 1757.420 19.215 1758.320 345.440 ;
        RECT 1762.120 19.215 1803.620 345.440 ;
        RECT 1807.420 19.215 1808.320 401.335 ;
        RECT 1812.120 354.015 1903.620 401.335 ;
        RECT 1812.120 19.215 1853.620 354.015 ;
        RECT 1857.420 19.215 1858.320 354.015 ;
        RECT 1862.120 19.215 1903.620 354.015 ;
        RECT 1907.420 19.215 1908.320 401.335 ;
        RECT 1912.120 1939.665 1953.620 3507.945 ;
        RECT 1957.420 1995.520 1958.320 3507.945 ;
        RECT 1962.120 1995.520 2003.620 3507.945 ;
        RECT 1957.420 1939.665 2003.620 1995.520 ;
        RECT 2007.420 1978.785 2008.320 3507.945 ;
        RECT 2012.120 1978.785 2053.620 3507.945 ;
        RECT 2057.420 1978.785 2058.320 3507.945 ;
        RECT 2062.120 1978.785 2103.620 3507.945 ;
        RECT 2007.420 1939.665 2103.620 1978.785 ;
        RECT 2107.420 1939.665 2108.320 3507.945 ;
        RECT 2112.120 1939.665 2153.620 3507.945 ;
        RECT 2157.420 1939.665 2158.320 3507.945 ;
        RECT 2162.120 1995.080 2203.620 3507.945 ;
        RECT 2207.420 1995.080 2208.320 3507.945 ;
        RECT 2162.120 1939.665 2208.320 1995.080 ;
        RECT 1912.120 1934.905 2208.320 1939.665 ;
        RECT 2212.120 1993.985 2253.620 3507.945 ;
        RECT 2257.420 1993.985 2258.320 3507.945 ;
        RECT 2262.120 1995.080 2303.620 3507.945 ;
        RECT 2307.420 1995.080 2308.320 3507.945 ;
        RECT 2312.120 1995.080 2353.620 3507.945 ;
        RECT 2262.120 1993.985 2353.620 1995.080 ;
        RECT 2212.120 1934.905 2353.620 1993.985 ;
        RECT 1912.120 405.415 2353.620 1934.905 ;
        RECT 1912.120 401.335 2208.320 405.415 ;
        RECT 1912.120 19.215 1953.620 401.335 ;
        RECT 1957.420 345.440 2003.620 401.335 ;
        RECT 1957.420 19.215 1958.320 345.440 ;
        RECT 1962.120 19.215 2003.620 345.440 ;
        RECT 2007.420 19.215 2008.320 401.335 ;
        RECT 2012.120 19.215 2053.620 401.335 ;
        RECT 2057.420 19.215 2058.320 401.335 ;
        RECT 2062.120 354.015 2153.620 401.335 ;
        RECT 2062.120 19.215 2103.620 354.015 ;
        RECT 2107.420 19.215 2108.320 354.015 ;
        RECT 2112.120 19.215 2153.620 354.015 ;
        RECT 2157.420 19.215 2158.320 401.335 ;
        RECT 2162.120 340.000 2208.320 401.335 ;
        RECT 2162.120 19.215 2203.620 340.000 ;
        RECT 2207.420 19.215 2208.320 340.000 ;
        RECT 2212.120 19.215 2253.620 405.415 ;
        RECT 2257.420 19.215 2258.320 405.415 ;
        RECT 2262.120 340.000 2353.620 405.415 ;
        RECT 2262.120 19.215 2303.620 340.000 ;
        RECT 2307.420 19.215 2308.320 340.000 ;
        RECT 2312.120 19.215 2353.620 340.000 ;
        RECT 2357.420 19.215 2358.320 3507.945 ;
        RECT 2362.120 1899.080 2403.620 3507.945 ;
        RECT 2407.420 1899.080 2408.320 3507.945 ;
        RECT 2412.120 1899.080 2453.620 3507.945 ;
        RECT 2457.420 1899.080 2458.320 3507.945 ;
        RECT 2462.120 1899.080 2503.620 3507.945 ;
        RECT 2507.420 1899.080 2508.320 3507.945 ;
        RECT 2512.120 1899.700 2553.620 3507.945 ;
        RECT 2557.420 1899.700 2558.320 3507.945 ;
        RECT 2562.120 1899.700 2603.620 3507.945 ;
        RECT 2607.420 1899.700 2608.320 3507.945 ;
        RECT 2612.120 1899.700 2653.620 3507.945 ;
        RECT 2657.420 1899.700 2658.320 3507.945 ;
        RECT 2662.120 1899.700 2703.620 3507.945 ;
        RECT 2707.420 1899.700 2708.320 3507.945 ;
        RECT 2712.120 1899.700 2753.620 3507.945 ;
        RECT 2512.120 1899.080 2753.620 1899.700 ;
        RECT 2757.420 1899.080 2758.320 3507.945 ;
        RECT 2762.120 1899.080 2803.620 3507.945 ;
        RECT 2807.420 1899.080 2808.320 3507.945 ;
        RECT 2812.120 1899.080 2853.620 3507.945 ;
        RECT 2857.420 1899.080 2858.320 3507.945 ;
        RECT 2862.120 1899.080 2873.160 3507.945 ;
        RECT 2362.120 1482.420 2873.160 1899.080 ;
        RECT 2362.120 1379.080 2403.620 1482.420 ;
        RECT 2407.420 1379.080 2408.320 1482.420 ;
        RECT 2412.120 1379.080 2453.620 1482.420 ;
        RECT 2457.420 1379.080 2458.320 1482.420 ;
        RECT 2462.120 1481.800 2753.620 1482.420 ;
        RECT 2462.120 1379.080 2503.620 1481.800 ;
        RECT 2507.420 1379.080 2508.320 1481.800 ;
        RECT 2512.120 1379.700 2553.620 1481.800 ;
        RECT 2557.420 1379.700 2558.320 1481.800 ;
        RECT 2562.120 1379.700 2603.620 1481.800 ;
        RECT 2607.420 1379.700 2608.320 1481.800 ;
        RECT 2612.120 1379.700 2653.620 1481.800 ;
        RECT 2657.420 1379.700 2658.320 1481.800 ;
        RECT 2662.120 1379.700 2703.620 1481.800 ;
        RECT 2707.420 1379.700 2708.320 1481.800 ;
        RECT 2712.120 1379.700 2753.620 1481.800 ;
        RECT 2512.120 1379.080 2753.620 1379.700 ;
        RECT 2757.420 1379.080 2758.320 1482.420 ;
        RECT 2762.120 1481.800 2853.620 1482.420 ;
        RECT 2762.120 1379.080 2803.620 1481.800 ;
        RECT 2807.420 1379.080 2808.320 1481.800 ;
        RECT 2812.120 1379.080 2853.620 1481.800 ;
        RECT 2857.420 1379.080 2858.320 1482.420 ;
        RECT 2862.120 1379.080 2873.160 1482.420 ;
        RECT 2362.120 962.420 2873.160 1379.080 ;
        RECT 2362.120 858.980 2403.620 962.420 ;
        RECT 2407.420 859.080 2408.320 962.420 ;
        RECT 2412.120 859.080 2453.620 962.420 ;
        RECT 2407.420 858.980 2453.620 859.080 ;
        RECT 2457.420 859.080 2458.320 962.420 ;
        RECT 2462.120 961.800 2753.620 962.420 ;
        RECT 2462.120 859.080 2503.620 961.800 ;
        RECT 2457.420 858.980 2503.620 859.080 ;
        RECT 2507.420 859.080 2508.320 961.800 ;
        RECT 2512.120 859.700 2553.620 961.800 ;
        RECT 2557.420 859.700 2558.320 961.800 ;
        RECT 2562.120 859.700 2603.620 961.800 ;
        RECT 2607.420 859.700 2608.320 961.800 ;
        RECT 2612.120 859.700 2653.620 961.800 ;
        RECT 2657.420 859.700 2658.320 961.800 ;
        RECT 2662.120 859.700 2703.620 961.800 ;
        RECT 2707.420 859.700 2708.320 961.800 ;
        RECT 2712.120 859.700 2753.620 961.800 ;
        RECT 2512.120 859.080 2753.620 859.700 ;
        RECT 2507.420 858.980 2753.620 859.080 ;
        RECT 2757.420 859.080 2758.320 962.420 ;
        RECT 2762.120 961.800 2853.620 962.420 ;
        RECT 2762.120 859.080 2803.620 961.800 ;
        RECT 2757.420 858.980 2803.620 859.080 ;
        RECT 2807.420 859.080 2808.320 961.800 ;
        RECT 2812.120 859.080 2853.620 961.800 ;
        RECT 2807.420 858.980 2853.620 859.080 ;
        RECT 2857.420 859.080 2858.320 962.420 ;
        RECT 2862.120 859.080 2873.160 962.420 ;
        RECT 2857.420 858.980 2873.160 859.080 ;
        RECT 2362.120 442.420 2873.160 858.980 ;
        RECT 2362.120 19.215 2403.620 442.420 ;
        RECT 2407.420 19.215 2408.320 442.420 ;
        RECT 2412.120 19.215 2453.620 442.420 ;
        RECT 2457.420 19.215 2458.320 442.420 ;
        RECT 2462.120 441.800 2753.620 442.420 ;
        RECT 2462.120 19.215 2503.620 441.800 ;
        RECT 2507.420 19.215 2508.320 441.800 ;
        RECT 2512.120 19.215 2553.620 441.800 ;
        RECT 2557.420 19.215 2558.320 441.800 ;
        RECT 2562.120 19.215 2603.620 441.800 ;
        RECT 2607.420 19.215 2608.320 441.800 ;
        RECT 2612.120 19.215 2653.620 441.800 ;
        RECT 2657.420 19.215 2658.320 441.800 ;
        RECT 2662.120 19.215 2703.620 441.800 ;
        RECT 2707.420 19.215 2708.320 441.800 ;
        RECT 2712.120 19.215 2753.620 441.800 ;
        RECT 2757.420 19.215 2758.320 442.420 ;
        RECT 2762.120 441.800 2853.620 442.420 ;
        RECT 2762.120 19.215 2803.620 441.800 ;
        RECT 2807.420 19.215 2808.320 441.800 ;
        RECT 2812.120 19.215 2853.620 441.800 ;
        RECT 2857.420 19.215 2858.320 442.420 ;
        RECT 2862.120 19.215 2873.160 442.420 ;
      LAYER met5 ;
        RECT 72.340 2568.680 890.900 2579.700 ;
        RECT 72.340 2518.680 890.900 2557.780 ;
        RECT 72.340 2468.680 890.900 2507.780 ;
        RECT 72.340 2418.680 890.900 2457.780 ;
        RECT 72.340 2368.680 890.900 2407.780 ;
        RECT 72.340 2318.680 890.900 2357.780 ;
        RECT 72.340 2268.680 890.900 2307.780 ;
        RECT 72.340 2218.680 890.900 2257.780 ;
        RECT 72.340 2168.680 890.900 2207.780 ;
        RECT 72.340 2118.680 890.900 2157.780 ;
        RECT 72.340 2068.680 890.900 2107.780 ;
        RECT 72.340 2018.680 890.900 2057.780 ;
        RECT 72.340 1968.680 890.900 2007.780 ;
        RECT 72.340 1918.680 890.900 1957.780 ;
        RECT 72.340 1868.680 890.900 1907.780 ;
        RECT 72.340 1818.680 890.900 1857.780 ;
        RECT 72.340 1768.680 890.900 1807.780 ;
        RECT 72.340 1718.680 890.900 1757.780 ;
        RECT 72.340 1668.680 890.900 1707.780 ;
        RECT 72.340 1618.680 890.900 1657.780 ;
        RECT 72.340 1568.680 890.900 1607.780 ;
        RECT 72.340 1518.680 890.900 1557.780 ;
        RECT 72.340 1468.680 890.900 1507.780 ;
        RECT 72.340 1418.680 890.900 1457.780 ;
        RECT 72.340 1368.680 890.900 1407.780 ;
        RECT 72.340 1318.680 890.900 1357.780 ;
        RECT 72.340 1268.680 890.900 1307.780 ;
        RECT 72.340 1218.680 890.900 1257.780 ;
        RECT 72.340 1168.680 890.900 1207.780 ;
        RECT 72.340 1118.680 890.900 1157.780 ;
        RECT 72.340 1068.680 890.900 1107.780 ;
        RECT 72.340 1018.680 890.900 1057.780 ;
        RECT 72.340 968.680 890.900 1007.780 ;
        RECT 72.340 918.680 890.900 957.780 ;
        RECT 72.340 868.680 890.900 907.780 ;
        RECT 72.340 818.680 890.900 857.780 ;
        RECT 72.340 768.680 890.900 807.780 ;
        RECT 72.340 718.680 890.900 757.780 ;
        RECT 72.340 668.680 890.900 707.780 ;
        RECT 72.340 618.680 890.900 657.780 ;
        RECT 72.340 568.680 890.900 607.780 ;
        RECT 72.340 518.680 890.900 557.780 ;
        RECT 72.340 468.680 890.900 507.780 ;
        RECT 72.340 418.680 890.900 457.780 ;
        RECT 72.340 368.680 890.900 407.780 ;
        RECT 72.340 318.680 890.900 357.780 ;
        RECT 72.340 279.700 890.900 307.780 ;
  END
END user_project_wrapper
END LIBRARY

