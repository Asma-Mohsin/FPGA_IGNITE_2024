module eFPGA
    #(
        parameter MaxFramesPerCol=20,
        parameter FrameBitsPerRow=32,
        parameter NoConfigBits=0
    )
    (
        input Tile_X1Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X1Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X1Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X2Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X2Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X3Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X3Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X4Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X4Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X5Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X5Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X6Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X6Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN0, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN1, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN10, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN11, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN12, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN13, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN14, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN15, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN16, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN17, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN18, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN19, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN2, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN3, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN4, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN5, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN6, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN7, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN8, //EXTERNAL
        input Tile_X7Y0_UIO_TOP_UIN9, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT0, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT1, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT10, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT11, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT12, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT13, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT14, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT15, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT16, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT17, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT18, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT19, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT2, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT3, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT4, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT5, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT6, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT7, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT8, //EXTERNAL
        output Tile_X7Y0_UIO_TOP_UOUT9, //EXTERNAL
        input Tile_X0Y1_A_O_top, //EXTERNAL
        output Tile_X0Y1_A_I_top, //EXTERNAL
        output Tile_X0Y1_A_T_top, //EXTERNAL
        input Tile_X0Y1_B_O_top, //EXTERNAL
        output Tile_X0Y1_B_I_top, //EXTERNAL
        output Tile_X0Y1_B_T_top, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y1_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y1_B_config_C_bit3, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D0_I0, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D0_I1, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D0_I2, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D0_I3, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D1_I0, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D1_I1, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D1_I2, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D1_I3, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D2_I0, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D2_I1, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D2_I2, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D2_I3, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D3_I0, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D3_I1, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D3_I2, //EXTERNAL
        input Tile_X8Y1_RAM2FAB_D3_I3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D0_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D0_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D0_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D0_O3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D1_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D1_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D1_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D1_O3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D2_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D2_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D2_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D2_O3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D3_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D3_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D3_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_D3_O3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A0_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A0_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A0_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A0_O3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A1_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A1_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A1_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_A1_O3, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_C_O0, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_C_O1, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_C_O2, //EXTERNAL
        output Tile_X8Y1_FAB2RAM_C_O3, //EXTERNAL
        output Tile_X8Y1_Config_accessC_bit0, //EXTERNAL
        output Tile_X8Y1_Config_accessC_bit1, //EXTERNAL
        output Tile_X8Y1_Config_accessC_bit2, //EXTERNAL
        output Tile_X8Y1_Config_accessC_bit3, //EXTERNAL
        input Tile_X0Y2_A_O_top, //EXTERNAL
        output Tile_X0Y2_A_I_top, //EXTERNAL
        output Tile_X0Y2_A_T_top, //EXTERNAL
        input Tile_X0Y2_B_O_top, //EXTERNAL
        output Tile_X0Y2_B_I_top, //EXTERNAL
        output Tile_X0Y2_B_T_top, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y2_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y2_B_config_C_bit3, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D0_I0, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D0_I1, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D0_I2, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D0_I3, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D1_I0, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D1_I1, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D1_I2, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D1_I3, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D2_I0, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D2_I1, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D2_I2, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D2_I3, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D3_I0, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D3_I1, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D3_I2, //EXTERNAL
        input Tile_X8Y2_RAM2FAB_D3_I3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D0_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D0_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D0_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D0_O3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D1_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D1_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D1_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D1_O3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D2_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D2_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D2_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D2_O3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D3_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D3_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D3_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_D3_O3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A0_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A0_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A0_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A0_O3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A1_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A1_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A1_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_A1_O3, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_C_O0, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_C_O1, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_C_O2, //EXTERNAL
        output Tile_X8Y2_FAB2RAM_C_O3, //EXTERNAL
        output Tile_X8Y2_Config_accessC_bit0, //EXTERNAL
        output Tile_X8Y2_Config_accessC_bit1, //EXTERNAL
        output Tile_X8Y2_Config_accessC_bit2, //EXTERNAL
        output Tile_X8Y2_Config_accessC_bit3, //EXTERNAL
        input Tile_X0Y3_A_O_top, //EXTERNAL
        output Tile_X0Y3_A_I_top, //EXTERNAL
        output Tile_X0Y3_A_T_top, //EXTERNAL
        input Tile_X0Y3_B_O_top, //EXTERNAL
        output Tile_X0Y3_B_I_top, //EXTERNAL
        output Tile_X0Y3_B_T_top, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y3_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y3_B_config_C_bit3, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D0_I0, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D0_I1, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D0_I2, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D0_I3, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D1_I0, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D1_I1, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D1_I2, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D1_I3, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D2_I0, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D2_I1, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D2_I2, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D2_I3, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D3_I0, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D3_I1, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D3_I2, //EXTERNAL
        input Tile_X8Y3_RAM2FAB_D3_I3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D0_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D0_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D0_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D0_O3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D1_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D1_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D1_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D1_O3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D2_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D2_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D2_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D2_O3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D3_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D3_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D3_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_D3_O3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A0_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A0_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A0_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A0_O3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A1_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A1_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A1_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_A1_O3, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_C_O0, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_C_O1, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_C_O2, //EXTERNAL
        output Tile_X8Y3_FAB2RAM_C_O3, //EXTERNAL
        output Tile_X8Y3_Config_accessC_bit0, //EXTERNAL
        output Tile_X8Y3_Config_accessC_bit1, //EXTERNAL
        output Tile_X8Y3_Config_accessC_bit2, //EXTERNAL
        output Tile_X8Y3_Config_accessC_bit3, //EXTERNAL
        input Tile_X0Y4_A_O_top, //EXTERNAL
        output Tile_X0Y4_A_I_top, //EXTERNAL
        output Tile_X0Y4_A_T_top, //EXTERNAL
        input Tile_X0Y4_B_O_top, //EXTERNAL
        output Tile_X0Y4_B_I_top, //EXTERNAL
        output Tile_X0Y4_B_T_top, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y4_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y4_B_config_C_bit3, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D0_I0, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D0_I1, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D0_I2, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D0_I3, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D1_I0, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D1_I1, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D1_I2, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D1_I3, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D2_I0, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D2_I1, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D2_I2, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D2_I3, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D3_I0, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D3_I1, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D3_I2, //EXTERNAL
        input Tile_X8Y4_RAM2FAB_D3_I3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D0_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D0_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D0_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D0_O3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D1_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D1_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D1_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D1_O3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D2_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D2_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D2_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D2_O3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D3_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D3_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D3_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_D3_O3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A0_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A0_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A0_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A0_O3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A1_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A1_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A1_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_A1_O3, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_C_O0, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_C_O1, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_C_O2, //EXTERNAL
        output Tile_X8Y4_FAB2RAM_C_O3, //EXTERNAL
        output Tile_X8Y4_Config_accessC_bit0, //EXTERNAL
        output Tile_X8Y4_Config_accessC_bit1, //EXTERNAL
        output Tile_X8Y4_Config_accessC_bit2, //EXTERNAL
        output Tile_X8Y4_Config_accessC_bit3, //EXTERNAL
        input Tile_X0Y5_A_O_top, //EXTERNAL
        output Tile_X0Y5_A_I_top, //EXTERNAL
        output Tile_X0Y5_A_T_top, //EXTERNAL
        input Tile_X0Y5_B_O_top, //EXTERNAL
        output Tile_X0Y5_B_I_top, //EXTERNAL
        output Tile_X0Y5_B_T_top, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y5_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y5_B_config_C_bit3, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D0_I0, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D0_I1, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D0_I2, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D0_I3, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D1_I0, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D1_I1, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D1_I2, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D1_I3, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D2_I0, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D2_I1, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D2_I2, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D2_I3, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D3_I0, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D3_I1, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D3_I2, //EXTERNAL
        input Tile_X8Y5_RAM2FAB_D3_I3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D0_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D0_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D0_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D0_O3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D1_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D1_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D1_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D1_O3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D2_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D2_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D2_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D2_O3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D3_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D3_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D3_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_D3_O3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A0_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A0_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A0_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A0_O3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A1_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A1_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A1_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_A1_O3, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_C_O0, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_C_O1, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_C_O2, //EXTERNAL
        output Tile_X8Y5_FAB2RAM_C_O3, //EXTERNAL
        output Tile_X8Y5_Config_accessC_bit0, //EXTERNAL
        output Tile_X8Y5_Config_accessC_bit1, //EXTERNAL
        output Tile_X8Y5_Config_accessC_bit2, //EXTERNAL
        output Tile_X8Y5_Config_accessC_bit3, //EXTERNAL
        input Tile_X0Y6_A_O_top, //EXTERNAL
        output Tile_X0Y6_A_I_top, //EXTERNAL
        output Tile_X0Y6_A_T_top, //EXTERNAL
        input Tile_X0Y6_B_O_top, //EXTERNAL
        output Tile_X0Y6_B_I_top, //EXTERNAL
        output Tile_X0Y6_B_T_top, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit0, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit1, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit2, //EXTERNAL
        output Tile_X0Y6_A_config_C_bit3, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit0, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit1, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit2, //EXTERNAL
        output Tile_X0Y6_B_config_C_bit3, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D0_I0, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D0_I1, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D0_I2, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D0_I3, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D1_I0, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D1_I1, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D1_I2, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D1_I3, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D2_I0, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D2_I1, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D2_I2, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D2_I3, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D3_I0, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D3_I1, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D3_I2, //EXTERNAL
        input Tile_X8Y6_RAM2FAB_D3_I3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D0_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D0_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D0_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D0_O3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D1_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D1_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D1_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D1_O3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D2_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D2_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D2_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D2_O3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D3_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D3_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D3_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_D3_O3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A0_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A0_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A0_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A0_O3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A1_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A1_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A1_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_A1_O3, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_C_O0, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_C_O1, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_C_O2, //EXTERNAL
        output Tile_X8Y6_FAB2RAM_C_O3, //EXTERNAL
        output Tile_X8Y6_Config_accessC_bit0, //EXTERNAL
        output Tile_X8Y6_Config_accessC_bit1, //EXTERNAL
        output Tile_X8Y6_Config_accessC_bit2, //EXTERNAL
        output Tile_X8Y6_Config_accessC_bit3, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X1Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X1Y7_UIO_BOT_UOUT9, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X2Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X2Y7_UIO_BOT_UOUT9, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X3Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X3Y7_UIO_BOT_UOUT9, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X4Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X4Y7_UIO_BOT_UOUT9, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X5Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X5Y7_UIO_BOT_UOUT9, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X6Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X6Y7_UIO_BOT_UOUT9, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN0, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN1, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN10, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN11, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN12, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN13, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN14, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN15, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN16, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN17, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN18, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN19, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN2, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN3, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN4, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN5, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN6, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN7, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN8, //EXTERNAL
        input Tile_X7Y7_UIO_BOT_UIN9, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT0, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT1, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT10, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT11, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT12, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT13, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT14, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT15, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT16, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT17, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT18, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT19, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT2, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT3, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT4, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT5, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT6, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT7, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT8, //EXTERNAL
        output Tile_X7Y7_UIO_BOT_UOUT9, //EXTERNAL
        input [(FrameBitsPerRow*8)-1:0] FrameData, //CONFIG_PORT
        input [(MaxFramesPerCol*9)-1:0] FrameStrobe, //CONFIG_PORT
        input UserCLK
);

 //signal declarations

wire Tile_X0Y0_UserCLKo;
wire Tile_X1Y0_UserCLKo;
wire Tile_X2Y0_UserCLKo;
wire Tile_X3Y0_UserCLKo;
wire Tile_X4Y0_UserCLKo;
wire Tile_X5Y0_UserCLKo;
wire Tile_X6Y0_UserCLKo;
wire Tile_X7Y0_UserCLKo;
wire Tile_X8Y0_UserCLKo;
wire Tile_X0Y1_UserCLKo;
wire Tile_X1Y1_UserCLKo;
wire Tile_X2Y1_UserCLKo;
wire Tile_X3Y1_UserCLKo;
wire Tile_X4Y1_UserCLKo;
wire Tile_X5Y1_UserCLKo;
wire Tile_X6Y1_UserCLKo;
wire Tile_X7Y1_UserCLKo;
wire Tile_X8Y1_UserCLKo;
wire Tile_X0Y2_UserCLKo;
wire Tile_X1Y2_UserCLKo;
wire Tile_X2Y2_UserCLKo;
wire Tile_X3Y2_UserCLKo;
wire Tile_X4Y2_UserCLKo;
wire Tile_X5Y2_UserCLKo;
wire Tile_X6Y2_UserCLKo;
wire Tile_X7Y2_UserCLKo;
wire Tile_X8Y2_UserCLKo;
wire Tile_X0Y3_UserCLKo;
wire Tile_X1Y3_UserCLKo;
wire Tile_X2Y3_UserCLKo;
wire Tile_X3Y3_UserCLKo;
wire Tile_X4Y3_UserCLKo;
wire Tile_X5Y3_UserCLKo;
wire Tile_X6Y3_UserCLKo;
wire Tile_X7Y3_UserCLKo;
wire Tile_X8Y3_UserCLKo;
wire Tile_X0Y4_UserCLKo;
wire Tile_X1Y4_UserCLKo;
wire Tile_X2Y4_UserCLKo;
wire Tile_X3Y4_UserCLKo;
wire Tile_X4Y4_UserCLKo;
wire Tile_X5Y4_UserCLKo;
wire Tile_X6Y4_UserCLKo;
wire Tile_X7Y4_UserCLKo;
wire Tile_X8Y4_UserCLKo;
wire Tile_X0Y5_UserCLKo;
wire Tile_X1Y5_UserCLKo;
wire Tile_X2Y5_UserCLKo;
wire Tile_X3Y5_UserCLKo;
wire Tile_X4Y5_UserCLKo;
wire Tile_X5Y5_UserCLKo;
wire Tile_X6Y5_UserCLKo;
wire Tile_X7Y5_UserCLKo;
wire Tile_X8Y5_UserCLKo;
wire Tile_X0Y6_UserCLKo;
wire Tile_X1Y6_UserCLKo;
wire Tile_X2Y6_UserCLKo;
wire Tile_X3Y6_UserCLKo;
wire Tile_X4Y6_UserCLKo;
wire Tile_X5Y6_UserCLKo;
wire Tile_X6Y6_UserCLKo;
wire Tile_X7Y6_UserCLKo;
wire Tile_X8Y6_UserCLKo;
wire Tile_X0Y7_UserCLKo;
wire Tile_X1Y7_UserCLKo;
wire Tile_X2Y7_UserCLKo;
wire Tile_X3Y7_UserCLKo;
wire Tile_X4Y7_UserCLKo;
wire Tile_X5Y7_UserCLKo;
wire Tile_X6Y7_UserCLKo;
wire Tile_X7Y7_UserCLKo;
wire Tile_X8Y7_UserCLKo;
 //configuration signal declarations

wire[FrameBitsPerRow -1:0] Tile_Y0_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y1_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y2_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y3_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y4_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y5_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y6_FrameData;
wire[FrameBitsPerRow -1:0] Tile_Y7_FrameData;
wire[MaxFramesPerCol - 1:0] Tile_X0_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X1_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X2_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X3_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X4_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X5_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X6_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X7_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Tile_X8_FrameStrobe;
wire[FrameBitsPerRow - 1:0] Tile_X0Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X6Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X7Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X8Y7_FrameData_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X6Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X7Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X8Y8_FrameStrobe_O;
 //tile-to-tile signal declarations
wire[3:0] Tile_X1Y0_S1BEG;
wire[7:0] Tile_X1Y0_S2BEG;
wire[7:0] Tile_X1Y0_S2BEGb;
wire[15:0] Tile_X1Y0_S4BEG;
wire[15:0] Tile_X1Y0_SS4BEG;
wire[3:0] Tile_X2Y0_S1BEG;
wire[7:0] Tile_X2Y0_S2BEG;
wire[7:0] Tile_X2Y0_S2BEGb;
wire[15:0] Tile_X2Y0_S4BEG;
wire[15:0] Tile_X2Y0_SS4BEG;
wire[3:0] Tile_X3Y0_S1BEG;
wire[7:0] Tile_X3Y0_S2BEG;
wire[7:0] Tile_X3Y0_S2BEGb;
wire[15:0] Tile_X3Y0_S4BEG;
wire[15:0] Tile_X3Y0_SS4BEG;
wire[3:0] Tile_X4Y0_S1BEG;
wire[7:0] Tile_X4Y0_S2BEG;
wire[7:0] Tile_X4Y0_S2BEGb;
wire[15:0] Tile_X4Y0_S4BEG;
wire[15:0] Tile_X4Y0_SS4BEG;
wire[3:0] Tile_X5Y0_S1BEG;
wire[7:0] Tile_X5Y0_S2BEG;
wire[7:0] Tile_X5Y0_S2BEGb;
wire[15:0] Tile_X5Y0_S4BEG;
wire[15:0] Tile_X5Y0_SS4BEG;
wire[3:0] Tile_X6Y0_S1BEG;
wire[7:0] Tile_X6Y0_S2BEG;
wire[7:0] Tile_X6Y0_S2BEGb;
wire[15:0] Tile_X6Y0_S4BEG;
wire[15:0] Tile_X6Y0_SS4BEG;
wire[3:0] Tile_X7Y0_S1BEG;
wire[7:0] Tile_X7Y0_S2BEG;
wire[7:0] Tile_X7Y0_S2BEGb;
wire[15:0] Tile_X7Y0_S4BEG;
wire[15:0] Tile_X7Y0_SS4BEG;
wire[3:0] Tile_X8Y0_S1BEG;
wire[7:0] Tile_X8Y0_S2BEG;
wire[7:0] Tile_X8Y0_S2BEGb;
wire[15:0] Tile_X8Y0_S4BEG;
wire[3:0] Tile_X0Y1_E1BEG;
wire[7:0] Tile_X0Y1_E2BEG;
wire[7:0] Tile_X0Y1_E2BEGb;
wire[15:0] Tile_X0Y1_EE4BEG;
wire[11:0] Tile_X0Y1_E6BEG;
wire[3:0] Tile_X1Y1_N1BEG;
wire[7:0] Tile_X1Y1_N2BEG;
wire[7:0] Tile_X1Y1_N2BEGb;
wire[15:0] Tile_X1Y1_N4BEG;
wire[15:0] Tile_X1Y1_NN4BEG;
wire[0:0] Tile_X1Y1_Co;
wire[3:0] Tile_X1Y1_E1BEG;
wire[7:0] Tile_X1Y1_E2BEG;
wire[7:0] Tile_X1Y1_E2BEGb;
wire[15:0] Tile_X1Y1_EE4BEG;
wire[11:0] Tile_X1Y1_E6BEG;
wire[3:0] Tile_X1Y1_S1BEG;
wire[7:0] Tile_X1Y1_S2BEG;
wire[7:0] Tile_X1Y1_S2BEGb;
wire[15:0] Tile_X1Y1_S4BEG;
wire[15:0] Tile_X1Y1_SS4BEG;
wire[3:0] Tile_X1Y1_W1BEG;
wire[7:0] Tile_X1Y1_W2BEG;
wire[7:0] Tile_X1Y1_W2BEGb;
wire[15:0] Tile_X1Y1_WW4BEG;
wire[11:0] Tile_X1Y1_W6BEG;
wire[3:0] Tile_X2Y1_N1BEG;
wire[7:0] Tile_X2Y1_N2BEG;
wire[7:0] Tile_X2Y1_N2BEGb;
wire[15:0] Tile_X2Y1_N4BEG;
wire[15:0] Tile_X2Y1_NN4BEG;
wire[0:0] Tile_X2Y1_Co;
wire[3:0] Tile_X2Y1_E1BEG;
wire[7:0] Tile_X2Y1_E2BEG;
wire[7:0] Tile_X2Y1_E2BEGb;
wire[15:0] Tile_X2Y1_EE4BEG;
wire[11:0] Tile_X2Y1_E6BEG;
wire[3:0] Tile_X2Y1_S1BEG;
wire[7:0] Tile_X2Y1_S2BEG;
wire[7:0] Tile_X2Y1_S2BEGb;
wire[15:0] Tile_X2Y1_S4BEG;
wire[15:0] Tile_X2Y1_SS4BEG;
wire[3:0] Tile_X2Y1_W1BEG;
wire[7:0] Tile_X2Y1_W2BEG;
wire[7:0] Tile_X2Y1_W2BEGb;
wire[15:0] Tile_X2Y1_WW4BEG;
wire[11:0] Tile_X2Y1_W6BEG;
wire[3:0] Tile_X3Y1_N1BEG;
wire[7:0] Tile_X3Y1_N2BEG;
wire[7:0] Tile_X3Y1_N2BEGb;
wire[15:0] Tile_X3Y1_N4BEG;
wire[15:0] Tile_X3Y1_NN4BEG;
wire[0:0] Tile_X3Y1_Co;
wire[3:0] Tile_X3Y1_E1BEG;
wire[7:0] Tile_X3Y1_E2BEG;
wire[7:0] Tile_X3Y1_E2BEGb;
wire[15:0] Tile_X3Y1_EE4BEG;
wire[11:0] Tile_X3Y1_E6BEG;
wire[3:0] Tile_X3Y1_S1BEG;
wire[7:0] Tile_X3Y1_S2BEG;
wire[7:0] Tile_X3Y1_S2BEGb;
wire[15:0] Tile_X3Y1_S4BEG;
wire[15:0] Tile_X3Y1_SS4BEG;
wire[3:0] Tile_X3Y1_W1BEG;
wire[7:0] Tile_X3Y1_W2BEG;
wire[7:0] Tile_X3Y1_W2BEGb;
wire[15:0] Tile_X3Y1_WW4BEG;
wire[11:0] Tile_X3Y1_W6BEG;
wire[3:0] Tile_X4Y1_N1BEG;
wire[7:0] Tile_X4Y1_N2BEG;
wire[7:0] Tile_X4Y1_N2BEGb;
wire[15:0] Tile_X4Y1_N4BEG;
wire[15:0] Tile_X4Y1_NN4BEG;
wire[0:0] Tile_X4Y1_Co;
wire[3:0] Tile_X4Y1_E1BEG;
wire[7:0] Tile_X4Y1_E2BEG;
wire[7:0] Tile_X4Y1_E2BEGb;
wire[15:0] Tile_X4Y1_EE4BEG;
wire[11:0] Tile_X4Y1_E6BEG;
wire[3:0] Tile_X4Y1_S1BEG;
wire[7:0] Tile_X4Y1_S2BEG;
wire[7:0] Tile_X4Y1_S2BEGb;
wire[15:0] Tile_X4Y1_S4BEG;
wire[15:0] Tile_X4Y1_SS4BEG;
wire[3:0] Tile_X4Y1_W1BEG;
wire[7:0] Tile_X4Y1_W2BEG;
wire[7:0] Tile_X4Y1_W2BEGb;
wire[15:0] Tile_X4Y1_WW4BEG;
wire[11:0] Tile_X4Y1_W6BEG;
wire[3:0] Tile_X5Y1_N1BEG;
wire[7:0] Tile_X5Y1_N2BEG;
wire[7:0] Tile_X5Y1_N2BEGb;
wire[15:0] Tile_X5Y1_N4BEG;
wire[15:0] Tile_X5Y1_NN4BEG;
wire[0:0] Tile_X5Y1_Co;
wire[3:0] Tile_X5Y1_E1BEG;
wire[7:0] Tile_X5Y1_E2BEG;
wire[7:0] Tile_X5Y1_E2BEGb;
wire[15:0] Tile_X5Y1_EE4BEG;
wire[11:0] Tile_X5Y1_E6BEG;
wire[3:0] Tile_X5Y1_S1BEG;
wire[7:0] Tile_X5Y1_S2BEG;
wire[7:0] Tile_X5Y1_S2BEGb;
wire[15:0] Tile_X5Y1_S4BEG;
wire[15:0] Tile_X5Y1_SS4BEG;
wire[3:0] Tile_X5Y1_W1BEG;
wire[7:0] Tile_X5Y1_W2BEG;
wire[7:0] Tile_X5Y1_W2BEGb;
wire[15:0] Tile_X5Y1_WW4BEG;
wire[11:0] Tile_X5Y1_W6BEG;
wire[3:0] Tile_X6Y1_N1BEG;
wire[7:0] Tile_X6Y1_N2BEG;
wire[7:0] Tile_X6Y1_N2BEGb;
wire[15:0] Tile_X6Y1_N4BEG;
wire[15:0] Tile_X6Y1_NN4BEG;
wire[0:0] Tile_X6Y1_Co;
wire[3:0] Tile_X6Y1_E1BEG;
wire[7:0] Tile_X6Y1_E2BEG;
wire[7:0] Tile_X6Y1_E2BEGb;
wire[15:0] Tile_X6Y1_EE4BEG;
wire[11:0] Tile_X6Y1_E6BEG;
wire[3:0] Tile_X6Y1_S1BEG;
wire[7:0] Tile_X6Y1_S2BEG;
wire[7:0] Tile_X6Y1_S2BEGb;
wire[15:0] Tile_X6Y1_S4BEG;
wire[15:0] Tile_X6Y1_SS4BEG;
wire[3:0] Tile_X6Y1_W1BEG;
wire[7:0] Tile_X6Y1_W2BEG;
wire[7:0] Tile_X6Y1_W2BEGb;
wire[15:0] Tile_X6Y1_WW4BEG;
wire[11:0] Tile_X6Y1_W6BEG;
wire[3:0] Tile_X7Y1_N1BEG;
wire[7:0] Tile_X7Y1_N2BEG;
wire[7:0] Tile_X7Y1_N2BEGb;
wire[15:0] Tile_X7Y1_N4BEG;
wire[15:0] Tile_X7Y1_NN4BEG;
wire[0:0] Tile_X7Y1_Co;
wire[3:0] Tile_X7Y1_E1BEG;
wire[7:0] Tile_X7Y1_E2BEG;
wire[7:0] Tile_X7Y1_E2BEGb;
wire[15:0] Tile_X7Y1_EE4BEG;
wire[11:0] Tile_X7Y1_E6BEG;
wire[3:0] Tile_X7Y1_S1BEG;
wire[7:0] Tile_X7Y1_S2BEG;
wire[7:0] Tile_X7Y1_S2BEGb;
wire[15:0] Tile_X7Y1_S4BEG;
wire[15:0] Tile_X7Y1_SS4BEG;
wire[3:0] Tile_X7Y1_W1BEG;
wire[7:0] Tile_X7Y1_W2BEG;
wire[7:0] Tile_X7Y1_W2BEGb;
wire[15:0] Tile_X7Y1_WW4BEG;
wire[11:0] Tile_X7Y1_W6BEG;
wire[3:0] Tile_X8Y1_N1BEG;
wire[7:0] Tile_X8Y1_N2BEG;
wire[7:0] Tile_X8Y1_N2BEGb;
wire[15:0] Tile_X8Y1_N4BEG;
wire[3:0] Tile_X8Y1_S1BEG;
wire[7:0] Tile_X8Y1_S2BEG;
wire[7:0] Tile_X8Y1_S2BEGb;
wire[15:0] Tile_X8Y1_S4BEG;
wire[3:0] Tile_X8Y1_W1BEG;
wire[7:0] Tile_X8Y1_W2BEG;
wire[7:0] Tile_X8Y1_W2BEGb;
wire[15:0] Tile_X8Y1_WW4BEG;
wire[11:0] Tile_X8Y1_W6BEG;
wire[3:0] Tile_X0Y2_E1BEG;
wire[7:0] Tile_X0Y2_E2BEG;
wire[7:0] Tile_X0Y2_E2BEGb;
wire[15:0] Tile_X0Y2_EE4BEG;
wire[11:0] Tile_X0Y2_E6BEG;
wire[3:0] Tile_X1Y2_N1BEG;
wire[7:0] Tile_X1Y2_N2BEG;
wire[7:0] Tile_X1Y2_N2BEGb;
wire[15:0] Tile_X1Y2_N4BEG;
wire[15:0] Tile_X1Y2_NN4BEG;
wire[0:0] Tile_X1Y2_Co;
wire[3:0] Tile_X1Y2_E1BEG;
wire[7:0] Tile_X1Y2_E2BEG;
wire[7:0] Tile_X1Y2_E2BEGb;
wire[15:0] Tile_X1Y2_EE4BEG;
wire[11:0] Tile_X1Y2_E6BEG;
wire[3:0] Tile_X1Y2_S1BEG;
wire[7:0] Tile_X1Y2_S2BEG;
wire[7:0] Tile_X1Y2_S2BEGb;
wire[15:0] Tile_X1Y2_S4BEG;
wire[15:0] Tile_X1Y2_SS4BEG;
wire[3:0] Tile_X1Y2_W1BEG;
wire[7:0] Tile_X1Y2_W2BEG;
wire[7:0] Tile_X1Y2_W2BEGb;
wire[15:0] Tile_X1Y2_WW4BEG;
wire[11:0] Tile_X1Y2_W6BEG;
wire[3:0] Tile_X2Y2_N1BEG;
wire[7:0] Tile_X2Y2_N2BEG;
wire[7:0] Tile_X2Y2_N2BEGb;
wire[15:0] Tile_X2Y2_N4BEG;
wire[15:0] Tile_X2Y2_NN4BEG;
wire[0:0] Tile_X2Y2_Co;
wire[3:0] Tile_X2Y2_E1BEG;
wire[7:0] Tile_X2Y2_E2BEG;
wire[7:0] Tile_X2Y2_E2BEGb;
wire[15:0] Tile_X2Y2_EE4BEG;
wire[11:0] Tile_X2Y2_E6BEG;
wire[3:0] Tile_X2Y2_S1BEG;
wire[7:0] Tile_X2Y2_S2BEG;
wire[7:0] Tile_X2Y2_S2BEGb;
wire[15:0] Tile_X2Y2_S4BEG;
wire[15:0] Tile_X2Y2_SS4BEG;
wire[3:0] Tile_X2Y2_W1BEG;
wire[7:0] Tile_X2Y2_W2BEG;
wire[7:0] Tile_X2Y2_W2BEGb;
wire[15:0] Tile_X2Y2_WW4BEG;
wire[11:0] Tile_X2Y2_W6BEG;
wire[3:0] Tile_X3Y2_N1BEG;
wire[7:0] Tile_X3Y2_N2BEG;
wire[7:0] Tile_X3Y2_N2BEGb;
wire[15:0] Tile_X3Y2_N4BEG;
wire[15:0] Tile_X3Y2_NN4BEG;
wire[0:0] Tile_X3Y2_Co;
wire[3:0] Tile_X3Y2_E1BEG;
wire[7:0] Tile_X3Y2_E2BEG;
wire[7:0] Tile_X3Y2_E2BEGb;
wire[15:0] Tile_X3Y2_EE4BEG;
wire[11:0] Tile_X3Y2_E6BEG;
wire[3:0] Tile_X3Y2_S1BEG;
wire[7:0] Tile_X3Y2_S2BEG;
wire[7:0] Tile_X3Y2_S2BEGb;
wire[15:0] Tile_X3Y2_S4BEG;
wire[15:0] Tile_X3Y2_SS4BEG;
wire[3:0] Tile_X3Y2_W1BEG;
wire[7:0] Tile_X3Y2_W2BEG;
wire[7:0] Tile_X3Y2_W2BEGb;
wire[15:0] Tile_X3Y2_WW4BEG;
wire[11:0] Tile_X3Y2_W6BEG;
wire[3:0] Tile_X4Y2_N1BEG;
wire[7:0] Tile_X4Y2_N2BEG;
wire[7:0] Tile_X4Y2_N2BEGb;
wire[15:0] Tile_X4Y2_N4BEG;
wire[15:0] Tile_X4Y2_NN4BEG;
wire[0:0] Tile_X4Y2_Co;
wire[3:0] Tile_X4Y2_E1BEG;
wire[7:0] Tile_X4Y2_E2BEG;
wire[7:0] Tile_X4Y2_E2BEGb;
wire[15:0] Tile_X4Y2_EE4BEG;
wire[11:0] Tile_X4Y2_E6BEG;
wire[3:0] Tile_X4Y2_S1BEG;
wire[7:0] Tile_X4Y2_S2BEG;
wire[7:0] Tile_X4Y2_S2BEGb;
wire[15:0] Tile_X4Y2_S4BEG;
wire[15:0] Tile_X4Y2_SS4BEG;
wire[3:0] Tile_X4Y2_W1BEG;
wire[7:0] Tile_X4Y2_W2BEG;
wire[7:0] Tile_X4Y2_W2BEGb;
wire[15:0] Tile_X4Y2_WW4BEG;
wire[11:0] Tile_X4Y2_W6BEG;
wire[3:0] Tile_X5Y2_N1BEG;
wire[7:0] Tile_X5Y2_N2BEG;
wire[7:0] Tile_X5Y2_N2BEGb;
wire[15:0] Tile_X5Y2_N4BEG;
wire[15:0] Tile_X5Y2_NN4BEG;
wire[0:0] Tile_X5Y2_Co;
wire[3:0] Tile_X5Y2_E1BEG;
wire[7:0] Tile_X5Y2_E2BEG;
wire[7:0] Tile_X5Y2_E2BEGb;
wire[15:0] Tile_X5Y2_EE4BEG;
wire[11:0] Tile_X5Y2_E6BEG;
wire[3:0] Tile_X5Y2_S1BEG;
wire[7:0] Tile_X5Y2_S2BEG;
wire[7:0] Tile_X5Y2_S2BEGb;
wire[15:0] Tile_X5Y2_S4BEG;
wire[15:0] Tile_X5Y2_SS4BEG;
wire[3:0] Tile_X5Y2_W1BEG;
wire[7:0] Tile_X5Y2_W2BEG;
wire[7:0] Tile_X5Y2_W2BEGb;
wire[15:0] Tile_X5Y2_WW4BEG;
wire[11:0] Tile_X5Y2_W6BEG;
wire[3:0] Tile_X6Y2_N1BEG;
wire[7:0] Tile_X6Y2_N2BEG;
wire[7:0] Tile_X6Y2_N2BEGb;
wire[15:0] Tile_X6Y2_N4BEG;
wire[15:0] Tile_X6Y2_NN4BEG;
wire[0:0] Tile_X6Y2_Co;
wire[3:0] Tile_X6Y2_E1BEG;
wire[7:0] Tile_X6Y2_E2BEG;
wire[7:0] Tile_X6Y2_E2BEGb;
wire[15:0] Tile_X6Y2_EE4BEG;
wire[11:0] Tile_X6Y2_E6BEG;
wire[3:0] Tile_X6Y2_S1BEG;
wire[7:0] Tile_X6Y2_S2BEG;
wire[7:0] Tile_X6Y2_S2BEGb;
wire[15:0] Tile_X6Y2_S4BEG;
wire[15:0] Tile_X6Y2_SS4BEG;
wire[3:0] Tile_X6Y2_W1BEG;
wire[7:0] Tile_X6Y2_W2BEG;
wire[7:0] Tile_X6Y2_W2BEGb;
wire[15:0] Tile_X6Y2_WW4BEG;
wire[11:0] Tile_X6Y2_W6BEG;
wire[3:0] Tile_X7Y2_N1BEG;
wire[7:0] Tile_X7Y2_N2BEG;
wire[7:0] Tile_X7Y2_N2BEGb;
wire[15:0] Tile_X7Y2_N4BEG;
wire[15:0] Tile_X7Y2_NN4BEG;
wire[0:0] Tile_X7Y2_Co;
wire[3:0] Tile_X7Y2_E1BEG;
wire[7:0] Tile_X7Y2_E2BEG;
wire[7:0] Tile_X7Y2_E2BEGb;
wire[15:0] Tile_X7Y2_EE4BEG;
wire[11:0] Tile_X7Y2_E6BEG;
wire[3:0] Tile_X7Y2_S1BEG;
wire[7:0] Tile_X7Y2_S2BEG;
wire[7:0] Tile_X7Y2_S2BEGb;
wire[15:0] Tile_X7Y2_S4BEG;
wire[15:0] Tile_X7Y2_SS4BEG;
wire[3:0] Tile_X7Y2_W1BEG;
wire[7:0] Tile_X7Y2_W2BEG;
wire[7:0] Tile_X7Y2_W2BEGb;
wire[15:0] Tile_X7Y2_WW4BEG;
wire[11:0] Tile_X7Y2_W6BEG;
wire[3:0] Tile_X8Y2_N1BEG;
wire[7:0] Tile_X8Y2_N2BEG;
wire[7:0] Tile_X8Y2_N2BEGb;
wire[15:0] Tile_X8Y2_N4BEG;
wire[3:0] Tile_X8Y2_S1BEG;
wire[7:0] Tile_X8Y2_S2BEG;
wire[7:0] Tile_X8Y2_S2BEGb;
wire[15:0] Tile_X8Y2_S4BEG;
wire[3:0] Tile_X8Y2_W1BEG;
wire[7:0] Tile_X8Y2_W2BEG;
wire[7:0] Tile_X8Y2_W2BEGb;
wire[15:0] Tile_X8Y2_WW4BEG;
wire[11:0] Tile_X8Y2_W6BEG;
wire[3:0] Tile_X0Y3_E1BEG;
wire[7:0] Tile_X0Y3_E2BEG;
wire[7:0] Tile_X0Y3_E2BEGb;
wire[15:0] Tile_X0Y3_EE4BEG;
wire[11:0] Tile_X0Y3_E6BEG;
wire[3:0] Tile_X1Y3_N1BEG;
wire[7:0] Tile_X1Y3_N2BEG;
wire[7:0] Tile_X1Y3_N2BEGb;
wire[15:0] Tile_X1Y3_N4BEG;
wire[15:0] Tile_X1Y3_NN4BEG;
wire[0:0] Tile_X1Y3_Co;
wire[3:0] Tile_X1Y3_E1BEG;
wire[7:0] Tile_X1Y3_E2BEG;
wire[7:0] Tile_X1Y3_E2BEGb;
wire[15:0] Tile_X1Y3_EE4BEG;
wire[11:0] Tile_X1Y3_E6BEG;
wire[3:0] Tile_X1Y3_S1BEG;
wire[7:0] Tile_X1Y3_S2BEG;
wire[7:0] Tile_X1Y3_S2BEGb;
wire[15:0] Tile_X1Y3_S4BEG;
wire[15:0] Tile_X1Y3_SS4BEG;
wire[3:0] Tile_X1Y3_W1BEG;
wire[7:0] Tile_X1Y3_W2BEG;
wire[7:0] Tile_X1Y3_W2BEGb;
wire[15:0] Tile_X1Y3_WW4BEG;
wire[11:0] Tile_X1Y3_W6BEG;
wire[3:0] Tile_X2Y3_N1BEG;
wire[7:0] Tile_X2Y3_N2BEG;
wire[7:0] Tile_X2Y3_N2BEGb;
wire[15:0] Tile_X2Y3_N4BEG;
wire[15:0] Tile_X2Y3_NN4BEG;
wire[0:0] Tile_X2Y3_Co;
wire[3:0] Tile_X2Y3_E1BEG;
wire[7:0] Tile_X2Y3_E2BEG;
wire[7:0] Tile_X2Y3_E2BEGb;
wire[15:0] Tile_X2Y3_EE4BEG;
wire[11:0] Tile_X2Y3_E6BEG;
wire[3:0] Tile_X2Y3_S1BEG;
wire[7:0] Tile_X2Y3_S2BEG;
wire[7:0] Tile_X2Y3_S2BEGb;
wire[15:0] Tile_X2Y3_S4BEG;
wire[15:0] Tile_X2Y3_SS4BEG;
wire[3:0] Tile_X2Y3_W1BEG;
wire[7:0] Tile_X2Y3_W2BEG;
wire[7:0] Tile_X2Y3_W2BEGb;
wire[15:0] Tile_X2Y3_WW4BEG;
wire[11:0] Tile_X2Y3_W6BEG;
wire[3:0] Tile_X3Y3_N1BEG;
wire[7:0] Tile_X3Y3_N2BEG;
wire[7:0] Tile_X3Y3_N2BEGb;
wire[15:0] Tile_X3Y3_N4BEG;
wire[15:0] Tile_X3Y3_NN4BEG;
wire[0:0] Tile_X3Y3_Co;
wire[3:0] Tile_X3Y3_E1BEG;
wire[7:0] Tile_X3Y3_E2BEG;
wire[7:0] Tile_X3Y3_E2BEGb;
wire[15:0] Tile_X3Y3_EE4BEG;
wire[11:0] Tile_X3Y3_E6BEG;
wire[3:0] Tile_X3Y3_S1BEG;
wire[7:0] Tile_X3Y3_S2BEG;
wire[7:0] Tile_X3Y3_S2BEGb;
wire[15:0] Tile_X3Y3_S4BEG;
wire[15:0] Tile_X3Y3_SS4BEG;
wire[3:0] Tile_X3Y3_W1BEG;
wire[7:0] Tile_X3Y3_W2BEG;
wire[7:0] Tile_X3Y3_W2BEGb;
wire[15:0] Tile_X3Y3_WW4BEG;
wire[11:0] Tile_X3Y3_W6BEG;
wire[3:0] Tile_X4Y3_N1BEG;
wire[7:0] Tile_X4Y3_N2BEG;
wire[7:0] Tile_X4Y3_N2BEGb;
wire[15:0] Tile_X4Y3_N4BEG;
wire[15:0] Tile_X4Y3_NN4BEG;
wire[0:0] Tile_X4Y3_Co;
wire[3:0] Tile_X4Y3_E1BEG;
wire[7:0] Tile_X4Y3_E2BEG;
wire[7:0] Tile_X4Y3_E2BEGb;
wire[15:0] Tile_X4Y3_EE4BEG;
wire[11:0] Tile_X4Y3_E6BEG;
wire[3:0] Tile_X4Y3_S1BEG;
wire[7:0] Tile_X4Y3_S2BEG;
wire[7:0] Tile_X4Y3_S2BEGb;
wire[15:0] Tile_X4Y3_S4BEG;
wire[15:0] Tile_X4Y3_SS4BEG;
wire[3:0] Tile_X4Y3_W1BEG;
wire[7:0] Tile_X4Y3_W2BEG;
wire[7:0] Tile_X4Y3_W2BEGb;
wire[15:0] Tile_X4Y3_WW4BEG;
wire[11:0] Tile_X4Y3_W6BEG;
wire[3:0] Tile_X5Y3_N1BEG;
wire[7:0] Tile_X5Y3_N2BEG;
wire[7:0] Tile_X5Y3_N2BEGb;
wire[15:0] Tile_X5Y3_N4BEG;
wire[15:0] Tile_X5Y3_NN4BEG;
wire[0:0] Tile_X5Y3_Co;
wire[3:0] Tile_X5Y3_E1BEG;
wire[7:0] Tile_X5Y3_E2BEG;
wire[7:0] Tile_X5Y3_E2BEGb;
wire[15:0] Tile_X5Y3_EE4BEG;
wire[11:0] Tile_X5Y3_E6BEG;
wire[3:0] Tile_X5Y3_S1BEG;
wire[7:0] Tile_X5Y3_S2BEG;
wire[7:0] Tile_X5Y3_S2BEGb;
wire[15:0] Tile_X5Y3_S4BEG;
wire[15:0] Tile_X5Y3_SS4BEG;
wire[3:0] Tile_X5Y3_W1BEG;
wire[7:0] Tile_X5Y3_W2BEG;
wire[7:0] Tile_X5Y3_W2BEGb;
wire[15:0] Tile_X5Y3_WW4BEG;
wire[11:0] Tile_X5Y3_W6BEG;
wire[3:0] Tile_X6Y3_N1BEG;
wire[7:0] Tile_X6Y3_N2BEG;
wire[7:0] Tile_X6Y3_N2BEGb;
wire[15:0] Tile_X6Y3_N4BEG;
wire[15:0] Tile_X6Y3_NN4BEG;
wire[0:0] Tile_X6Y3_Co;
wire[3:0] Tile_X6Y3_E1BEG;
wire[7:0] Tile_X6Y3_E2BEG;
wire[7:0] Tile_X6Y3_E2BEGb;
wire[15:0] Tile_X6Y3_EE4BEG;
wire[11:0] Tile_X6Y3_E6BEG;
wire[3:0] Tile_X6Y3_S1BEG;
wire[7:0] Tile_X6Y3_S2BEG;
wire[7:0] Tile_X6Y3_S2BEGb;
wire[15:0] Tile_X6Y3_S4BEG;
wire[15:0] Tile_X6Y3_SS4BEG;
wire[3:0] Tile_X6Y3_W1BEG;
wire[7:0] Tile_X6Y3_W2BEG;
wire[7:0] Tile_X6Y3_W2BEGb;
wire[15:0] Tile_X6Y3_WW4BEG;
wire[11:0] Tile_X6Y3_W6BEG;
wire[3:0] Tile_X7Y3_N1BEG;
wire[7:0] Tile_X7Y3_N2BEG;
wire[7:0] Tile_X7Y3_N2BEGb;
wire[15:0] Tile_X7Y3_N4BEG;
wire[15:0] Tile_X7Y3_NN4BEG;
wire[0:0] Tile_X7Y3_Co;
wire[3:0] Tile_X7Y3_E1BEG;
wire[7:0] Tile_X7Y3_E2BEG;
wire[7:0] Tile_X7Y3_E2BEGb;
wire[15:0] Tile_X7Y3_EE4BEG;
wire[11:0] Tile_X7Y3_E6BEG;
wire[3:0] Tile_X7Y3_S1BEG;
wire[7:0] Tile_X7Y3_S2BEG;
wire[7:0] Tile_X7Y3_S2BEGb;
wire[15:0] Tile_X7Y3_S4BEG;
wire[15:0] Tile_X7Y3_SS4BEG;
wire[3:0] Tile_X7Y3_W1BEG;
wire[7:0] Tile_X7Y3_W2BEG;
wire[7:0] Tile_X7Y3_W2BEGb;
wire[15:0] Tile_X7Y3_WW4BEG;
wire[11:0] Tile_X7Y3_W6BEG;
wire[3:0] Tile_X8Y3_N1BEG;
wire[7:0] Tile_X8Y3_N2BEG;
wire[7:0] Tile_X8Y3_N2BEGb;
wire[15:0] Tile_X8Y3_N4BEG;
wire[3:0] Tile_X8Y3_S1BEG;
wire[7:0] Tile_X8Y3_S2BEG;
wire[7:0] Tile_X8Y3_S2BEGb;
wire[15:0] Tile_X8Y3_S4BEG;
wire[3:0] Tile_X8Y3_W1BEG;
wire[7:0] Tile_X8Y3_W2BEG;
wire[7:0] Tile_X8Y3_W2BEGb;
wire[15:0] Tile_X8Y3_WW4BEG;
wire[11:0] Tile_X8Y3_W6BEG;
wire[3:0] Tile_X0Y4_E1BEG;
wire[7:0] Tile_X0Y4_E2BEG;
wire[7:0] Tile_X0Y4_E2BEGb;
wire[15:0] Tile_X0Y4_EE4BEG;
wire[11:0] Tile_X0Y4_E6BEG;
wire[3:0] Tile_X1Y4_N1BEG;
wire[7:0] Tile_X1Y4_N2BEG;
wire[7:0] Tile_X1Y4_N2BEGb;
wire[15:0] Tile_X1Y4_N4BEG;
wire[15:0] Tile_X1Y4_NN4BEG;
wire[0:0] Tile_X1Y4_Co;
wire[3:0] Tile_X1Y4_E1BEG;
wire[7:0] Tile_X1Y4_E2BEG;
wire[7:0] Tile_X1Y4_E2BEGb;
wire[15:0] Tile_X1Y4_EE4BEG;
wire[11:0] Tile_X1Y4_E6BEG;
wire[3:0] Tile_X1Y4_S1BEG;
wire[7:0] Tile_X1Y4_S2BEG;
wire[7:0] Tile_X1Y4_S2BEGb;
wire[15:0] Tile_X1Y4_S4BEG;
wire[15:0] Tile_X1Y4_SS4BEG;
wire[3:0] Tile_X1Y4_W1BEG;
wire[7:0] Tile_X1Y4_W2BEG;
wire[7:0] Tile_X1Y4_W2BEGb;
wire[15:0] Tile_X1Y4_WW4BEG;
wire[11:0] Tile_X1Y4_W6BEG;
wire[3:0] Tile_X2Y4_N1BEG;
wire[7:0] Tile_X2Y4_N2BEG;
wire[7:0] Tile_X2Y4_N2BEGb;
wire[15:0] Tile_X2Y4_N4BEG;
wire[15:0] Tile_X2Y4_NN4BEG;
wire[0:0] Tile_X2Y4_Co;
wire[3:0] Tile_X2Y4_E1BEG;
wire[7:0] Tile_X2Y4_E2BEG;
wire[7:0] Tile_X2Y4_E2BEGb;
wire[15:0] Tile_X2Y4_EE4BEG;
wire[11:0] Tile_X2Y4_E6BEG;
wire[3:0] Tile_X2Y4_S1BEG;
wire[7:0] Tile_X2Y4_S2BEG;
wire[7:0] Tile_X2Y4_S2BEGb;
wire[15:0] Tile_X2Y4_S4BEG;
wire[15:0] Tile_X2Y4_SS4BEG;
wire[3:0] Tile_X2Y4_W1BEG;
wire[7:0] Tile_X2Y4_W2BEG;
wire[7:0] Tile_X2Y4_W2BEGb;
wire[15:0] Tile_X2Y4_WW4BEG;
wire[11:0] Tile_X2Y4_W6BEG;
wire[3:0] Tile_X3Y4_N1BEG;
wire[7:0] Tile_X3Y4_N2BEG;
wire[7:0] Tile_X3Y4_N2BEGb;
wire[15:0] Tile_X3Y4_N4BEG;
wire[15:0] Tile_X3Y4_NN4BEG;
wire[0:0] Tile_X3Y4_Co;
wire[3:0] Tile_X3Y4_E1BEG;
wire[7:0] Tile_X3Y4_E2BEG;
wire[7:0] Tile_X3Y4_E2BEGb;
wire[15:0] Tile_X3Y4_EE4BEG;
wire[11:0] Tile_X3Y4_E6BEG;
wire[3:0] Tile_X3Y4_S1BEG;
wire[7:0] Tile_X3Y4_S2BEG;
wire[7:0] Tile_X3Y4_S2BEGb;
wire[15:0] Tile_X3Y4_S4BEG;
wire[15:0] Tile_X3Y4_SS4BEG;
wire[3:0] Tile_X3Y4_W1BEG;
wire[7:0] Tile_X3Y4_W2BEG;
wire[7:0] Tile_X3Y4_W2BEGb;
wire[15:0] Tile_X3Y4_WW4BEG;
wire[11:0] Tile_X3Y4_W6BEG;
wire[3:0] Tile_X4Y4_N1BEG;
wire[7:0] Tile_X4Y4_N2BEG;
wire[7:0] Tile_X4Y4_N2BEGb;
wire[15:0] Tile_X4Y4_N4BEG;
wire[15:0] Tile_X4Y4_NN4BEG;
wire[0:0] Tile_X4Y4_Co;
wire[3:0] Tile_X4Y4_E1BEG;
wire[7:0] Tile_X4Y4_E2BEG;
wire[7:0] Tile_X4Y4_E2BEGb;
wire[15:0] Tile_X4Y4_EE4BEG;
wire[11:0] Tile_X4Y4_E6BEG;
wire[3:0] Tile_X4Y4_S1BEG;
wire[7:0] Tile_X4Y4_S2BEG;
wire[7:0] Tile_X4Y4_S2BEGb;
wire[15:0] Tile_X4Y4_S4BEG;
wire[15:0] Tile_X4Y4_SS4BEG;
wire[3:0] Tile_X4Y4_W1BEG;
wire[7:0] Tile_X4Y4_W2BEG;
wire[7:0] Tile_X4Y4_W2BEGb;
wire[15:0] Tile_X4Y4_WW4BEG;
wire[11:0] Tile_X4Y4_W6BEG;
wire[3:0] Tile_X5Y4_N1BEG;
wire[7:0] Tile_X5Y4_N2BEG;
wire[7:0] Tile_X5Y4_N2BEGb;
wire[15:0] Tile_X5Y4_N4BEG;
wire[15:0] Tile_X5Y4_NN4BEG;
wire[0:0] Tile_X5Y4_Co;
wire[3:0] Tile_X5Y4_E1BEG;
wire[7:0] Tile_X5Y4_E2BEG;
wire[7:0] Tile_X5Y4_E2BEGb;
wire[15:0] Tile_X5Y4_EE4BEG;
wire[11:0] Tile_X5Y4_E6BEG;
wire[3:0] Tile_X5Y4_S1BEG;
wire[7:0] Tile_X5Y4_S2BEG;
wire[7:0] Tile_X5Y4_S2BEGb;
wire[15:0] Tile_X5Y4_S4BEG;
wire[15:0] Tile_X5Y4_SS4BEG;
wire[3:0] Tile_X5Y4_W1BEG;
wire[7:0] Tile_X5Y4_W2BEG;
wire[7:0] Tile_X5Y4_W2BEGb;
wire[15:0] Tile_X5Y4_WW4BEG;
wire[11:0] Tile_X5Y4_W6BEG;
wire[3:0] Tile_X6Y4_N1BEG;
wire[7:0] Tile_X6Y4_N2BEG;
wire[7:0] Tile_X6Y4_N2BEGb;
wire[15:0] Tile_X6Y4_N4BEG;
wire[15:0] Tile_X6Y4_NN4BEG;
wire[0:0] Tile_X6Y4_Co;
wire[3:0] Tile_X6Y4_E1BEG;
wire[7:0] Tile_X6Y4_E2BEG;
wire[7:0] Tile_X6Y4_E2BEGb;
wire[15:0] Tile_X6Y4_EE4BEG;
wire[11:0] Tile_X6Y4_E6BEG;
wire[3:0] Tile_X6Y4_S1BEG;
wire[7:0] Tile_X6Y4_S2BEG;
wire[7:0] Tile_X6Y4_S2BEGb;
wire[15:0] Tile_X6Y4_S4BEG;
wire[15:0] Tile_X6Y4_SS4BEG;
wire[3:0] Tile_X6Y4_W1BEG;
wire[7:0] Tile_X6Y4_W2BEG;
wire[7:0] Tile_X6Y4_W2BEGb;
wire[15:0] Tile_X6Y4_WW4BEG;
wire[11:0] Tile_X6Y4_W6BEG;
wire[3:0] Tile_X7Y4_N1BEG;
wire[7:0] Tile_X7Y4_N2BEG;
wire[7:0] Tile_X7Y4_N2BEGb;
wire[15:0] Tile_X7Y4_N4BEG;
wire[15:0] Tile_X7Y4_NN4BEG;
wire[0:0] Tile_X7Y4_Co;
wire[3:0] Tile_X7Y4_E1BEG;
wire[7:0] Tile_X7Y4_E2BEG;
wire[7:0] Tile_X7Y4_E2BEGb;
wire[15:0] Tile_X7Y4_EE4BEG;
wire[11:0] Tile_X7Y4_E6BEG;
wire[3:0] Tile_X7Y4_S1BEG;
wire[7:0] Tile_X7Y4_S2BEG;
wire[7:0] Tile_X7Y4_S2BEGb;
wire[15:0] Tile_X7Y4_S4BEG;
wire[15:0] Tile_X7Y4_SS4BEG;
wire[3:0] Tile_X7Y4_W1BEG;
wire[7:0] Tile_X7Y4_W2BEG;
wire[7:0] Tile_X7Y4_W2BEGb;
wire[15:0] Tile_X7Y4_WW4BEG;
wire[11:0] Tile_X7Y4_W6BEG;
wire[3:0] Tile_X8Y4_N1BEG;
wire[7:0] Tile_X8Y4_N2BEG;
wire[7:0] Tile_X8Y4_N2BEGb;
wire[15:0] Tile_X8Y4_N4BEG;
wire[3:0] Tile_X8Y4_S1BEG;
wire[7:0] Tile_X8Y4_S2BEG;
wire[7:0] Tile_X8Y4_S2BEGb;
wire[15:0] Tile_X8Y4_S4BEG;
wire[3:0] Tile_X8Y4_W1BEG;
wire[7:0] Tile_X8Y4_W2BEG;
wire[7:0] Tile_X8Y4_W2BEGb;
wire[15:0] Tile_X8Y4_WW4BEG;
wire[11:0] Tile_X8Y4_W6BEG;
wire[3:0] Tile_X0Y5_E1BEG;
wire[7:0] Tile_X0Y5_E2BEG;
wire[7:0] Tile_X0Y5_E2BEGb;
wire[15:0] Tile_X0Y5_EE4BEG;
wire[11:0] Tile_X0Y5_E6BEG;
wire[3:0] Tile_X1Y5_N1BEG;
wire[7:0] Tile_X1Y5_N2BEG;
wire[7:0] Tile_X1Y5_N2BEGb;
wire[15:0] Tile_X1Y5_N4BEG;
wire[15:0] Tile_X1Y5_NN4BEG;
wire[0:0] Tile_X1Y5_Co;
wire[3:0] Tile_X1Y5_E1BEG;
wire[7:0] Tile_X1Y5_E2BEG;
wire[7:0] Tile_X1Y5_E2BEGb;
wire[15:0] Tile_X1Y5_EE4BEG;
wire[11:0] Tile_X1Y5_E6BEG;
wire[3:0] Tile_X1Y5_S1BEG;
wire[7:0] Tile_X1Y5_S2BEG;
wire[7:0] Tile_X1Y5_S2BEGb;
wire[15:0] Tile_X1Y5_S4BEG;
wire[15:0] Tile_X1Y5_SS4BEG;
wire[3:0] Tile_X1Y5_W1BEG;
wire[7:0] Tile_X1Y5_W2BEG;
wire[7:0] Tile_X1Y5_W2BEGb;
wire[15:0] Tile_X1Y5_WW4BEG;
wire[11:0] Tile_X1Y5_W6BEG;
wire[3:0] Tile_X2Y5_N1BEG;
wire[7:0] Tile_X2Y5_N2BEG;
wire[7:0] Tile_X2Y5_N2BEGb;
wire[15:0] Tile_X2Y5_N4BEG;
wire[15:0] Tile_X2Y5_NN4BEG;
wire[0:0] Tile_X2Y5_Co;
wire[3:0] Tile_X2Y5_E1BEG;
wire[7:0] Tile_X2Y5_E2BEG;
wire[7:0] Tile_X2Y5_E2BEGb;
wire[15:0] Tile_X2Y5_EE4BEG;
wire[11:0] Tile_X2Y5_E6BEG;
wire[3:0] Tile_X2Y5_S1BEG;
wire[7:0] Tile_X2Y5_S2BEG;
wire[7:0] Tile_X2Y5_S2BEGb;
wire[15:0] Tile_X2Y5_S4BEG;
wire[15:0] Tile_X2Y5_SS4BEG;
wire[3:0] Tile_X2Y5_W1BEG;
wire[7:0] Tile_X2Y5_W2BEG;
wire[7:0] Tile_X2Y5_W2BEGb;
wire[15:0] Tile_X2Y5_WW4BEG;
wire[11:0] Tile_X2Y5_W6BEG;
wire[3:0] Tile_X3Y5_N1BEG;
wire[7:0] Tile_X3Y5_N2BEG;
wire[7:0] Tile_X3Y5_N2BEGb;
wire[15:0] Tile_X3Y5_N4BEG;
wire[15:0] Tile_X3Y5_NN4BEG;
wire[0:0] Tile_X3Y5_Co;
wire[3:0] Tile_X3Y5_E1BEG;
wire[7:0] Tile_X3Y5_E2BEG;
wire[7:0] Tile_X3Y5_E2BEGb;
wire[15:0] Tile_X3Y5_EE4BEG;
wire[11:0] Tile_X3Y5_E6BEG;
wire[3:0] Tile_X3Y5_S1BEG;
wire[7:0] Tile_X3Y5_S2BEG;
wire[7:0] Tile_X3Y5_S2BEGb;
wire[15:0] Tile_X3Y5_S4BEG;
wire[15:0] Tile_X3Y5_SS4BEG;
wire[3:0] Tile_X3Y5_W1BEG;
wire[7:0] Tile_X3Y5_W2BEG;
wire[7:0] Tile_X3Y5_W2BEGb;
wire[15:0] Tile_X3Y5_WW4BEG;
wire[11:0] Tile_X3Y5_W6BEG;
wire[3:0] Tile_X4Y5_N1BEG;
wire[7:0] Tile_X4Y5_N2BEG;
wire[7:0] Tile_X4Y5_N2BEGb;
wire[15:0] Tile_X4Y5_N4BEG;
wire[15:0] Tile_X4Y5_NN4BEG;
wire[0:0] Tile_X4Y5_Co;
wire[3:0] Tile_X4Y5_E1BEG;
wire[7:0] Tile_X4Y5_E2BEG;
wire[7:0] Tile_X4Y5_E2BEGb;
wire[15:0] Tile_X4Y5_EE4BEG;
wire[11:0] Tile_X4Y5_E6BEG;
wire[3:0] Tile_X4Y5_S1BEG;
wire[7:0] Tile_X4Y5_S2BEG;
wire[7:0] Tile_X4Y5_S2BEGb;
wire[15:0] Tile_X4Y5_S4BEG;
wire[15:0] Tile_X4Y5_SS4BEG;
wire[3:0] Tile_X4Y5_W1BEG;
wire[7:0] Tile_X4Y5_W2BEG;
wire[7:0] Tile_X4Y5_W2BEGb;
wire[15:0] Tile_X4Y5_WW4BEG;
wire[11:0] Tile_X4Y5_W6BEG;
wire[3:0] Tile_X5Y5_N1BEG;
wire[7:0] Tile_X5Y5_N2BEG;
wire[7:0] Tile_X5Y5_N2BEGb;
wire[15:0] Tile_X5Y5_N4BEG;
wire[15:0] Tile_X5Y5_NN4BEG;
wire[0:0] Tile_X5Y5_Co;
wire[3:0] Tile_X5Y5_E1BEG;
wire[7:0] Tile_X5Y5_E2BEG;
wire[7:0] Tile_X5Y5_E2BEGb;
wire[15:0] Tile_X5Y5_EE4BEG;
wire[11:0] Tile_X5Y5_E6BEG;
wire[3:0] Tile_X5Y5_S1BEG;
wire[7:0] Tile_X5Y5_S2BEG;
wire[7:0] Tile_X5Y5_S2BEGb;
wire[15:0] Tile_X5Y5_S4BEG;
wire[15:0] Tile_X5Y5_SS4BEG;
wire[3:0] Tile_X5Y5_W1BEG;
wire[7:0] Tile_X5Y5_W2BEG;
wire[7:0] Tile_X5Y5_W2BEGb;
wire[15:0] Tile_X5Y5_WW4BEG;
wire[11:0] Tile_X5Y5_W6BEG;
wire[3:0] Tile_X6Y5_N1BEG;
wire[7:0] Tile_X6Y5_N2BEG;
wire[7:0] Tile_X6Y5_N2BEGb;
wire[15:0] Tile_X6Y5_N4BEG;
wire[15:0] Tile_X6Y5_NN4BEG;
wire[0:0] Tile_X6Y5_Co;
wire[3:0] Tile_X6Y5_E1BEG;
wire[7:0] Tile_X6Y5_E2BEG;
wire[7:0] Tile_X6Y5_E2BEGb;
wire[15:0] Tile_X6Y5_EE4BEG;
wire[11:0] Tile_X6Y5_E6BEG;
wire[3:0] Tile_X6Y5_S1BEG;
wire[7:0] Tile_X6Y5_S2BEG;
wire[7:0] Tile_X6Y5_S2BEGb;
wire[15:0] Tile_X6Y5_S4BEG;
wire[15:0] Tile_X6Y5_SS4BEG;
wire[3:0] Tile_X6Y5_W1BEG;
wire[7:0] Tile_X6Y5_W2BEG;
wire[7:0] Tile_X6Y5_W2BEGb;
wire[15:0] Tile_X6Y5_WW4BEG;
wire[11:0] Tile_X6Y5_W6BEG;
wire[3:0] Tile_X7Y5_N1BEG;
wire[7:0] Tile_X7Y5_N2BEG;
wire[7:0] Tile_X7Y5_N2BEGb;
wire[15:0] Tile_X7Y5_N4BEG;
wire[15:0] Tile_X7Y5_NN4BEG;
wire[0:0] Tile_X7Y5_Co;
wire[3:0] Tile_X7Y5_E1BEG;
wire[7:0] Tile_X7Y5_E2BEG;
wire[7:0] Tile_X7Y5_E2BEGb;
wire[15:0] Tile_X7Y5_EE4BEG;
wire[11:0] Tile_X7Y5_E6BEG;
wire[3:0] Tile_X7Y5_S1BEG;
wire[7:0] Tile_X7Y5_S2BEG;
wire[7:0] Tile_X7Y5_S2BEGb;
wire[15:0] Tile_X7Y5_S4BEG;
wire[15:0] Tile_X7Y5_SS4BEG;
wire[3:0] Tile_X7Y5_W1BEG;
wire[7:0] Tile_X7Y5_W2BEG;
wire[7:0] Tile_X7Y5_W2BEGb;
wire[15:0] Tile_X7Y5_WW4BEG;
wire[11:0] Tile_X7Y5_W6BEG;
wire[3:0] Tile_X8Y5_N1BEG;
wire[7:0] Tile_X8Y5_N2BEG;
wire[7:0] Tile_X8Y5_N2BEGb;
wire[15:0] Tile_X8Y5_N4BEG;
wire[3:0] Tile_X8Y5_S1BEG;
wire[7:0] Tile_X8Y5_S2BEG;
wire[7:0] Tile_X8Y5_S2BEGb;
wire[15:0] Tile_X8Y5_S4BEG;
wire[3:0] Tile_X8Y5_W1BEG;
wire[7:0] Tile_X8Y5_W2BEG;
wire[7:0] Tile_X8Y5_W2BEGb;
wire[15:0] Tile_X8Y5_WW4BEG;
wire[11:0] Tile_X8Y5_W6BEG;
wire[3:0] Tile_X0Y6_E1BEG;
wire[7:0] Tile_X0Y6_E2BEG;
wire[7:0] Tile_X0Y6_E2BEGb;
wire[15:0] Tile_X0Y6_EE4BEG;
wire[11:0] Tile_X0Y6_E6BEG;
wire[3:0] Tile_X1Y6_N1BEG;
wire[7:0] Tile_X1Y6_N2BEG;
wire[7:0] Tile_X1Y6_N2BEGb;
wire[15:0] Tile_X1Y6_N4BEG;
wire[15:0] Tile_X1Y6_NN4BEG;
wire[0:0] Tile_X1Y6_Co;
wire[3:0] Tile_X1Y6_E1BEG;
wire[7:0] Tile_X1Y6_E2BEG;
wire[7:0] Tile_X1Y6_E2BEGb;
wire[15:0] Tile_X1Y6_EE4BEG;
wire[11:0] Tile_X1Y6_E6BEG;
wire[3:0] Tile_X1Y6_S1BEG;
wire[7:0] Tile_X1Y6_S2BEG;
wire[7:0] Tile_X1Y6_S2BEGb;
wire[15:0] Tile_X1Y6_S4BEG;
wire[15:0] Tile_X1Y6_SS4BEG;
wire[3:0] Tile_X1Y6_W1BEG;
wire[7:0] Tile_X1Y6_W2BEG;
wire[7:0] Tile_X1Y6_W2BEGb;
wire[15:0] Tile_X1Y6_WW4BEG;
wire[11:0] Tile_X1Y6_W6BEG;
wire[3:0] Tile_X2Y6_N1BEG;
wire[7:0] Tile_X2Y6_N2BEG;
wire[7:0] Tile_X2Y6_N2BEGb;
wire[15:0] Tile_X2Y6_N4BEG;
wire[15:0] Tile_X2Y6_NN4BEG;
wire[0:0] Tile_X2Y6_Co;
wire[3:0] Tile_X2Y6_E1BEG;
wire[7:0] Tile_X2Y6_E2BEG;
wire[7:0] Tile_X2Y6_E2BEGb;
wire[15:0] Tile_X2Y6_EE4BEG;
wire[11:0] Tile_X2Y6_E6BEG;
wire[3:0] Tile_X2Y6_S1BEG;
wire[7:0] Tile_X2Y6_S2BEG;
wire[7:0] Tile_X2Y6_S2BEGb;
wire[15:0] Tile_X2Y6_S4BEG;
wire[15:0] Tile_X2Y6_SS4BEG;
wire[3:0] Tile_X2Y6_W1BEG;
wire[7:0] Tile_X2Y6_W2BEG;
wire[7:0] Tile_X2Y6_W2BEGb;
wire[15:0] Tile_X2Y6_WW4BEG;
wire[11:0] Tile_X2Y6_W6BEG;
wire[3:0] Tile_X3Y6_N1BEG;
wire[7:0] Tile_X3Y6_N2BEG;
wire[7:0] Tile_X3Y6_N2BEGb;
wire[15:0] Tile_X3Y6_N4BEG;
wire[15:0] Tile_X3Y6_NN4BEG;
wire[0:0] Tile_X3Y6_Co;
wire[3:0] Tile_X3Y6_E1BEG;
wire[7:0] Tile_X3Y6_E2BEG;
wire[7:0] Tile_X3Y6_E2BEGb;
wire[15:0] Tile_X3Y6_EE4BEG;
wire[11:0] Tile_X3Y6_E6BEG;
wire[3:0] Tile_X3Y6_S1BEG;
wire[7:0] Tile_X3Y6_S2BEG;
wire[7:0] Tile_X3Y6_S2BEGb;
wire[15:0] Tile_X3Y6_S4BEG;
wire[15:0] Tile_X3Y6_SS4BEG;
wire[3:0] Tile_X3Y6_W1BEG;
wire[7:0] Tile_X3Y6_W2BEG;
wire[7:0] Tile_X3Y6_W2BEGb;
wire[15:0] Tile_X3Y6_WW4BEG;
wire[11:0] Tile_X3Y6_W6BEG;
wire[3:0] Tile_X4Y6_N1BEG;
wire[7:0] Tile_X4Y6_N2BEG;
wire[7:0] Tile_X4Y6_N2BEGb;
wire[15:0] Tile_X4Y6_N4BEG;
wire[15:0] Tile_X4Y6_NN4BEG;
wire[0:0] Tile_X4Y6_Co;
wire[3:0] Tile_X4Y6_E1BEG;
wire[7:0] Tile_X4Y6_E2BEG;
wire[7:0] Tile_X4Y6_E2BEGb;
wire[15:0] Tile_X4Y6_EE4BEG;
wire[11:0] Tile_X4Y6_E6BEG;
wire[3:0] Tile_X4Y6_S1BEG;
wire[7:0] Tile_X4Y6_S2BEG;
wire[7:0] Tile_X4Y6_S2BEGb;
wire[15:0] Tile_X4Y6_S4BEG;
wire[15:0] Tile_X4Y6_SS4BEG;
wire[3:0] Tile_X4Y6_W1BEG;
wire[7:0] Tile_X4Y6_W2BEG;
wire[7:0] Tile_X4Y6_W2BEGb;
wire[15:0] Tile_X4Y6_WW4BEG;
wire[11:0] Tile_X4Y6_W6BEG;
wire[3:0] Tile_X5Y6_N1BEG;
wire[7:0] Tile_X5Y6_N2BEG;
wire[7:0] Tile_X5Y6_N2BEGb;
wire[15:0] Tile_X5Y6_N4BEG;
wire[15:0] Tile_X5Y6_NN4BEG;
wire[0:0] Tile_X5Y6_Co;
wire[3:0] Tile_X5Y6_E1BEG;
wire[7:0] Tile_X5Y6_E2BEG;
wire[7:0] Tile_X5Y6_E2BEGb;
wire[15:0] Tile_X5Y6_EE4BEG;
wire[11:0] Tile_X5Y6_E6BEG;
wire[3:0] Tile_X5Y6_S1BEG;
wire[7:0] Tile_X5Y6_S2BEG;
wire[7:0] Tile_X5Y6_S2BEGb;
wire[15:0] Tile_X5Y6_S4BEG;
wire[15:0] Tile_X5Y6_SS4BEG;
wire[3:0] Tile_X5Y6_W1BEG;
wire[7:0] Tile_X5Y6_W2BEG;
wire[7:0] Tile_X5Y6_W2BEGb;
wire[15:0] Tile_X5Y6_WW4BEG;
wire[11:0] Tile_X5Y6_W6BEG;
wire[3:0] Tile_X6Y6_N1BEG;
wire[7:0] Tile_X6Y6_N2BEG;
wire[7:0] Tile_X6Y6_N2BEGb;
wire[15:0] Tile_X6Y6_N4BEG;
wire[15:0] Tile_X6Y6_NN4BEG;
wire[0:0] Tile_X6Y6_Co;
wire[3:0] Tile_X6Y6_E1BEG;
wire[7:0] Tile_X6Y6_E2BEG;
wire[7:0] Tile_X6Y6_E2BEGb;
wire[15:0] Tile_X6Y6_EE4BEG;
wire[11:0] Tile_X6Y6_E6BEG;
wire[3:0] Tile_X6Y6_S1BEG;
wire[7:0] Tile_X6Y6_S2BEG;
wire[7:0] Tile_X6Y6_S2BEGb;
wire[15:0] Tile_X6Y6_S4BEG;
wire[15:0] Tile_X6Y6_SS4BEG;
wire[3:0] Tile_X6Y6_W1BEG;
wire[7:0] Tile_X6Y6_W2BEG;
wire[7:0] Tile_X6Y6_W2BEGb;
wire[15:0] Tile_X6Y6_WW4BEG;
wire[11:0] Tile_X6Y6_W6BEG;
wire[3:0] Tile_X7Y6_N1BEG;
wire[7:0] Tile_X7Y6_N2BEG;
wire[7:0] Tile_X7Y6_N2BEGb;
wire[15:0] Tile_X7Y6_N4BEG;
wire[15:0] Tile_X7Y6_NN4BEG;
wire[0:0] Tile_X7Y6_Co;
wire[3:0] Tile_X7Y6_E1BEG;
wire[7:0] Tile_X7Y6_E2BEG;
wire[7:0] Tile_X7Y6_E2BEGb;
wire[15:0] Tile_X7Y6_EE4BEG;
wire[11:0] Tile_X7Y6_E6BEG;
wire[3:0] Tile_X7Y6_S1BEG;
wire[7:0] Tile_X7Y6_S2BEG;
wire[7:0] Tile_X7Y6_S2BEGb;
wire[15:0] Tile_X7Y6_S4BEG;
wire[15:0] Tile_X7Y6_SS4BEG;
wire[3:0] Tile_X7Y6_W1BEG;
wire[7:0] Tile_X7Y6_W2BEG;
wire[7:0] Tile_X7Y6_W2BEGb;
wire[15:0] Tile_X7Y6_WW4BEG;
wire[11:0] Tile_X7Y6_W6BEG;
wire[3:0] Tile_X8Y6_N1BEG;
wire[7:0] Tile_X8Y6_N2BEG;
wire[7:0] Tile_X8Y6_N2BEGb;
wire[15:0] Tile_X8Y6_N4BEG;
wire[3:0] Tile_X8Y6_S1BEG;
wire[7:0] Tile_X8Y6_S2BEG;
wire[7:0] Tile_X8Y6_S2BEGb;
wire[15:0] Tile_X8Y6_S4BEG;
wire[3:0] Tile_X8Y6_W1BEG;
wire[7:0] Tile_X8Y6_W2BEG;
wire[7:0] Tile_X8Y6_W2BEGb;
wire[15:0] Tile_X8Y6_WW4BEG;
wire[11:0] Tile_X8Y6_W6BEG;
wire[3:0] Tile_X1Y7_N1BEG;
wire[7:0] Tile_X1Y7_N2BEG;
wire[7:0] Tile_X1Y7_N2BEGb;
wire[15:0] Tile_X1Y7_N4BEG;
wire[15:0] Tile_X1Y7_NN4BEG;
wire[0:0] Tile_X1Y7_Co;
wire[3:0] Tile_X2Y7_N1BEG;
wire[7:0] Tile_X2Y7_N2BEG;
wire[7:0] Tile_X2Y7_N2BEGb;
wire[15:0] Tile_X2Y7_N4BEG;
wire[15:0] Tile_X2Y7_NN4BEG;
wire[0:0] Tile_X2Y7_Co;
wire[3:0] Tile_X3Y7_N1BEG;
wire[7:0] Tile_X3Y7_N2BEG;
wire[7:0] Tile_X3Y7_N2BEGb;
wire[15:0] Tile_X3Y7_N4BEG;
wire[15:0] Tile_X3Y7_NN4BEG;
wire[0:0] Tile_X3Y7_Co;
wire[3:0] Tile_X4Y7_N1BEG;
wire[7:0] Tile_X4Y7_N2BEG;
wire[7:0] Tile_X4Y7_N2BEGb;
wire[15:0] Tile_X4Y7_N4BEG;
wire[15:0] Tile_X4Y7_NN4BEG;
wire[0:0] Tile_X4Y7_Co;
wire[3:0] Tile_X5Y7_N1BEG;
wire[7:0] Tile_X5Y7_N2BEG;
wire[7:0] Tile_X5Y7_N2BEGb;
wire[15:0] Tile_X5Y7_N4BEG;
wire[15:0] Tile_X5Y7_NN4BEG;
wire[0:0] Tile_X5Y7_Co;
wire[3:0] Tile_X6Y7_N1BEG;
wire[7:0] Tile_X6Y7_N2BEG;
wire[7:0] Tile_X6Y7_N2BEGb;
wire[15:0] Tile_X6Y7_N4BEG;
wire[15:0] Tile_X6Y7_NN4BEG;
wire[0:0] Tile_X6Y7_Co;
wire[3:0] Tile_X7Y7_N1BEG;
wire[7:0] Tile_X7Y7_N2BEG;
wire[7:0] Tile_X7Y7_N2BEGb;
wire[15:0] Tile_X7Y7_N4BEG;
wire[15:0] Tile_X7Y7_NN4BEG;
wire[0:0] Tile_X7Y7_Co;
wire[3:0] Tile_X8Y7_N1BEG;
wire[7:0] Tile_X8Y7_N2BEG;
wire[7:0] Tile_X8Y7_N2BEGb;
wire[15:0] Tile_X8Y7_N4BEG;

assign Tile_Y1_FrameData = FrameData[FrameBitsPerRow*(1+1)-1:FrameBitsPerRow*1];
assign Tile_Y2_FrameData = FrameData[FrameBitsPerRow*(2+1)-1:FrameBitsPerRow*2];
assign Tile_Y3_FrameData = FrameData[FrameBitsPerRow*(3+1)-1:FrameBitsPerRow*3];
assign Tile_Y4_FrameData = FrameData[FrameBitsPerRow*(4+1)-1:FrameBitsPerRow*4];
assign Tile_Y5_FrameData = FrameData[FrameBitsPerRow*(5+1)-1:FrameBitsPerRow*5];
assign Tile_Y6_FrameData = FrameData[FrameBitsPerRow*(6+1)-1:FrameBitsPerRow*6];
assign Tile_X0_FrameStrobe = FrameStrobe[MaxFramesPerCol*(0+1)-1:MaxFramesPerCol*0];
assign Tile_X1_FrameStrobe = FrameStrobe[MaxFramesPerCol*(1+1)-1:MaxFramesPerCol*1];
assign Tile_X2_FrameStrobe = FrameStrobe[MaxFramesPerCol*(2+1)-1:MaxFramesPerCol*2];
assign Tile_X3_FrameStrobe = FrameStrobe[MaxFramesPerCol*(3+1)-1:MaxFramesPerCol*3];
assign Tile_X4_FrameStrobe = FrameStrobe[MaxFramesPerCol*(4+1)-1:MaxFramesPerCol*4];
assign Tile_X5_FrameStrobe = FrameStrobe[MaxFramesPerCol*(5+1)-1:MaxFramesPerCol*5];
assign Tile_X6_FrameStrobe = FrameStrobe[MaxFramesPerCol*(6+1)-1:MaxFramesPerCol*6];
assign Tile_X7_FrameStrobe = FrameStrobe[MaxFramesPerCol*(7+1)-1:MaxFramesPerCol*7];
assign Tile_X8_FrameStrobe = FrameStrobe[MaxFramesPerCol*(8+1)-1:MaxFramesPerCol*8];

 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X1Y0_N_term_single (
    .N1END(Tile_X1Y1_N1BEG),
    .N2MID(Tile_X1Y1_N2BEG),
    .N2END(Tile_X1Y1_N2BEGb),
    .N4END(Tile_X1Y1_N4BEG),
    .NN4END(Tile_X1Y1_NN4BEG),
    .Ci(Tile_X1Y1_Co),
    .S1BEG(Tile_X1Y0_S1BEG),
    .S2BEG(Tile_X1Y0_S2BEG),
    .S2BEGb(Tile_X1Y0_S2BEGb),
    .S4BEG(Tile_X1Y0_S4BEG),
    .SS4BEG(Tile_X1Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X1Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X1Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X1Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X1Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X1Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X1Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X1Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X1Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X1Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X1Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X1Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X1Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X1Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X1Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X1Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X1Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X1Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X1Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X1Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X1Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X1Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X1Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X1Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X1Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X1Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X1Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X1Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X1Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X1Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X1Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X1Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X1Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X1Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X1Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X1Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X1Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X1Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X1Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X1Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X1Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X1Y1_UserCLKo),
    .UserCLKo(Tile_X1Y0_UserCLKo),
    .FrameStrobe(Tile_X1Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X2Y0_N_term_single (
    .N1END(Tile_X2Y1_N1BEG),
    .N2MID(Tile_X2Y1_N2BEG),
    .N2END(Tile_X2Y1_N2BEGb),
    .N4END(Tile_X2Y1_N4BEG),
    .NN4END(Tile_X2Y1_NN4BEG),
    .Ci(Tile_X2Y1_Co),
    .S1BEG(Tile_X2Y0_S1BEG),
    .S2BEG(Tile_X2Y0_S2BEG),
    .S2BEGb(Tile_X2Y0_S2BEGb),
    .S4BEG(Tile_X2Y0_S4BEG),
    .SS4BEG(Tile_X2Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X2Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X2Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X2Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X2Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X2Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X2Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X2Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X2Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X2Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X2Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X2Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X2Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X2Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X2Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X2Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X2Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X2Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X2Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X2Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X2Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X2Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X2Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X2Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X2Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X2Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X2Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X2Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X2Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X2Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X2Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X2Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X2Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X2Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X2Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X2Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X2Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X2Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X2Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X2Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X2Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X2Y1_UserCLKo),
    .UserCLKo(Tile_X2Y0_UserCLKo),
    .FrameStrobe(Tile_X2Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X3Y0_N_term_single (
    .N1END(Tile_X3Y1_N1BEG),
    .N2MID(Tile_X3Y1_N2BEG),
    .N2END(Tile_X3Y1_N2BEGb),
    .N4END(Tile_X3Y1_N4BEG),
    .NN4END(Tile_X3Y1_NN4BEG),
    .Ci(Tile_X3Y1_Co),
    .S1BEG(Tile_X3Y0_S1BEG),
    .S2BEG(Tile_X3Y0_S2BEG),
    .S2BEGb(Tile_X3Y0_S2BEGb),
    .S4BEG(Tile_X3Y0_S4BEG),
    .SS4BEG(Tile_X3Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X3Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X3Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X3Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X3Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X3Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X3Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X3Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X3Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X3Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X3Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X3Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X3Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X3Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X3Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X3Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X3Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X3Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X3Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X3Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X3Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X3Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X3Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X3Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X3Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X3Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X3Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X3Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X3Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X3Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X3Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X3Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X3Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X3Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X3Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X3Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X3Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X3Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X3Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X3Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X3Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X3Y1_UserCLKo),
    .UserCLKo(Tile_X3Y0_UserCLKo),
    .FrameStrobe(Tile_X3Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X4Y0_N_term_single (
    .N1END(Tile_X4Y1_N1BEG),
    .N2MID(Tile_X4Y1_N2BEG),
    .N2END(Tile_X4Y1_N2BEGb),
    .N4END(Tile_X4Y1_N4BEG),
    .NN4END(Tile_X4Y1_NN4BEG),
    .Ci(Tile_X4Y1_Co),
    .S1BEG(Tile_X4Y0_S1BEG),
    .S2BEG(Tile_X4Y0_S2BEG),
    .S2BEGb(Tile_X4Y0_S2BEGb),
    .S4BEG(Tile_X4Y0_S4BEG),
    .SS4BEG(Tile_X4Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X4Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X4Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X4Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X4Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X4Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X4Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X4Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X4Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X4Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X4Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X4Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X4Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X4Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X4Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X4Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X4Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X4Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X4Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X4Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X4Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X4Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X4Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X4Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X4Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X4Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X4Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X4Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X4Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X4Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X4Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X4Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X4Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X4Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X4Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X4Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X4Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X4Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X4Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X4Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X4Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X4Y1_UserCLKo),
    .UserCLKo(Tile_X4Y0_UserCLKo),
    .FrameStrobe(Tile_X4Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X5Y0_N_term_single (
    .N1END(Tile_X5Y1_N1BEG),
    .N2MID(Tile_X5Y1_N2BEG),
    .N2END(Tile_X5Y1_N2BEGb),
    .N4END(Tile_X5Y1_N4BEG),
    .NN4END(Tile_X5Y1_NN4BEG),
    .Ci(Tile_X5Y1_Co),
    .S1BEG(Tile_X5Y0_S1BEG),
    .S2BEG(Tile_X5Y0_S2BEG),
    .S2BEGb(Tile_X5Y0_S2BEGb),
    .S4BEG(Tile_X5Y0_S4BEG),
    .SS4BEG(Tile_X5Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X5Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X5Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X5Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X5Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X5Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X5Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X5Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X5Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X5Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X5Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X5Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X5Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X5Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X5Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X5Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X5Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X5Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X5Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X5Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X5Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X5Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X5Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X5Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X5Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X5Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X5Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X5Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X5Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X5Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X5Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X5Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X5Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X5Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X5Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X5Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X5Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X5Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X5Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X5Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X5Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X5Y1_UserCLKo),
    .UserCLKo(Tile_X5Y0_UserCLKo),
    .FrameStrobe(Tile_X5Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X6Y0_N_term_single (
    .N1END(Tile_X6Y1_N1BEG),
    .N2MID(Tile_X6Y1_N2BEG),
    .N2END(Tile_X6Y1_N2BEGb),
    .N4END(Tile_X6Y1_N4BEG),
    .NN4END(Tile_X6Y1_NN4BEG),
    .Ci(Tile_X6Y1_Co),
    .S1BEG(Tile_X6Y0_S1BEG),
    .S2BEG(Tile_X6Y0_S2BEG),
    .S2BEGb(Tile_X6Y0_S2BEGb),
    .S4BEG(Tile_X6Y0_S4BEG),
    .SS4BEG(Tile_X6Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X6Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X6Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X6Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X6Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X6Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X6Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X6Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X6Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X6Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X6Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X6Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X6Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X6Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X6Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X6Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X6Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X6Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X6Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X6Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X6Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X6Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X6Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X6Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X6Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X6Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X6Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X6Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X6Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X6Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X6Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X6Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X6Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X6Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X6Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X6Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X6Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X6Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X6Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X6Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X6Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X6Y1_UserCLKo),
    .UserCLKo(Tile_X6Y0_UserCLKo),
    .FrameStrobe(Tile_X6Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_single Tile_X7Y0_N_term_single (
    .N1END(Tile_X7Y1_N1BEG),
    .N2MID(Tile_X7Y1_N2BEG),
    .N2END(Tile_X7Y1_N2BEGb),
    .N4END(Tile_X7Y1_N4BEG),
    .NN4END(Tile_X7Y1_NN4BEG),
    .Ci(Tile_X7Y1_Co),
    .S1BEG(Tile_X7Y0_S1BEG),
    .S2BEG(Tile_X7Y0_S2BEG),
    .S2BEGb(Tile_X7Y0_S2BEGb),
    .S4BEG(Tile_X7Y0_S4BEG),
    .SS4BEG(Tile_X7Y0_SS4BEG),
    .UIO_TOP_UIN0(Tile_X7Y0_UIO_TOP_UIN0),
    .UIO_TOP_UIN1(Tile_X7Y0_UIO_TOP_UIN1),
    .UIO_TOP_UIN10(Tile_X7Y0_UIO_TOP_UIN10),
    .UIO_TOP_UIN11(Tile_X7Y0_UIO_TOP_UIN11),
    .UIO_TOP_UIN12(Tile_X7Y0_UIO_TOP_UIN12),
    .UIO_TOP_UIN13(Tile_X7Y0_UIO_TOP_UIN13),
    .UIO_TOP_UIN14(Tile_X7Y0_UIO_TOP_UIN14),
    .UIO_TOP_UIN15(Tile_X7Y0_UIO_TOP_UIN15),
    .UIO_TOP_UIN16(Tile_X7Y0_UIO_TOP_UIN16),
    .UIO_TOP_UIN17(Tile_X7Y0_UIO_TOP_UIN17),
    .UIO_TOP_UIN18(Tile_X7Y0_UIO_TOP_UIN18),
    .UIO_TOP_UIN19(Tile_X7Y0_UIO_TOP_UIN19),
    .UIO_TOP_UIN2(Tile_X7Y0_UIO_TOP_UIN2),
    .UIO_TOP_UIN3(Tile_X7Y0_UIO_TOP_UIN3),
    .UIO_TOP_UIN4(Tile_X7Y0_UIO_TOP_UIN4),
    .UIO_TOP_UIN5(Tile_X7Y0_UIO_TOP_UIN5),
    .UIO_TOP_UIN6(Tile_X7Y0_UIO_TOP_UIN6),
    .UIO_TOP_UIN7(Tile_X7Y0_UIO_TOP_UIN7),
    .UIO_TOP_UIN8(Tile_X7Y0_UIO_TOP_UIN8),
    .UIO_TOP_UIN9(Tile_X7Y0_UIO_TOP_UIN9),
    .UIO_TOP_UOUT0(Tile_X7Y0_UIO_TOP_UOUT0),
    .UIO_TOP_UOUT1(Tile_X7Y0_UIO_TOP_UOUT1),
    .UIO_TOP_UOUT10(Tile_X7Y0_UIO_TOP_UOUT10),
    .UIO_TOP_UOUT11(Tile_X7Y0_UIO_TOP_UOUT11),
    .UIO_TOP_UOUT12(Tile_X7Y0_UIO_TOP_UOUT12),
    .UIO_TOP_UOUT13(Tile_X7Y0_UIO_TOP_UOUT13),
    .UIO_TOP_UOUT14(Tile_X7Y0_UIO_TOP_UOUT14),
    .UIO_TOP_UOUT15(Tile_X7Y0_UIO_TOP_UOUT15),
    .UIO_TOP_UOUT16(Tile_X7Y0_UIO_TOP_UOUT16),
    .UIO_TOP_UOUT17(Tile_X7Y0_UIO_TOP_UOUT17),
    .UIO_TOP_UOUT18(Tile_X7Y0_UIO_TOP_UOUT18),
    .UIO_TOP_UOUT19(Tile_X7Y0_UIO_TOP_UOUT19),
    .UIO_TOP_UOUT2(Tile_X7Y0_UIO_TOP_UOUT2),
    .UIO_TOP_UOUT3(Tile_X7Y0_UIO_TOP_UOUT3),
    .UIO_TOP_UOUT4(Tile_X7Y0_UIO_TOP_UOUT4),
    .UIO_TOP_UOUT5(Tile_X7Y0_UIO_TOP_UOUT5),
    .UIO_TOP_UOUT6(Tile_X7Y0_UIO_TOP_UOUT6),
    .UIO_TOP_UOUT7(Tile_X7Y0_UIO_TOP_UOUT7),
    .UIO_TOP_UOUT8(Tile_X7Y0_UIO_TOP_UOUT8),
    .UIO_TOP_UOUT9(Tile_X7Y0_UIO_TOP_UOUT9),
    .UserCLK(Tile_X7Y1_UserCLKo),
    .UserCLKo(Tile_X7Y0_UserCLKo),
    .FrameStrobe(Tile_X7Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_term_RAM_IO Tile_X8Y0_N_term_RAM_IO (
    .N1END(Tile_X8Y1_N1BEG),
    .N2MID(Tile_X8Y1_N2BEG),
    .N2END(Tile_X8Y1_N2BEGb),
    .N4END(Tile_X8Y1_N4BEG),
    .S1BEG(Tile_X8Y0_S1BEG),
    .S2BEG(Tile_X8Y0_S2BEG),
    .S2BEGb(Tile_X8Y0_S2BEGb),
    .S4BEG(Tile_X8Y0_S4BEG),
    .UserCLK(Tile_X8Y1_UserCLKo),
    .UserCLKo(Tile_X8Y0_UserCLKo),
    .FrameStrobe(Tile_X8Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y1_Emulate_Bitstream)
    )
`endif
    Tile_X0Y1_W_IO
    (
    .W1END(Tile_X1Y1_W1BEG),
    .W2MID(Tile_X1Y1_W2BEG),
    .W2END(Tile_X1Y1_W2BEGb),
    .WW4END(Tile_X1Y1_WW4BEG),
    .W6END(Tile_X1Y1_W6BEG),
    .E1BEG(Tile_X0Y1_E1BEG),
    .E2BEG(Tile_X0Y1_E2BEG),
    .E2BEGb(Tile_X0Y1_E2BEGb),
    .EE4BEG(Tile_X0Y1_EE4BEG),
    .E6BEG(Tile_X0Y1_E6BEG),
    .A_O_top(Tile_X0Y1_A_O_top),
    .A_I_top(Tile_X0Y1_A_I_top),
    .A_T_top(Tile_X0Y1_A_T_top),
    .B_O_top(Tile_X0Y1_B_O_top),
    .B_I_top(Tile_X0Y1_B_I_top),
    .B_T_top(Tile_X0Y1_B_T_top),
    .A_config_C_bit0(Tile_X0Y1_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y1_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y1_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y1_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y1_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y1_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y1_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y1_B_config_C_bit3),
    .UserCLK(Tile_X0Y2_UserCLKo),
    .UserCLKo(Tile_X0Y1_UserCLKo),
    .FrameData(Tile_Y1_FrameData),
    .FrameData_O(Tile_X0Y1_FrameData_O),
    .FrameStrobe(Tile_X0Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y1_Emulate_Bitstream)
    )
`endif
    Tile_X1Y1_LUT4AB
    (
    .N1END(Tile_X1Y2_N1BEG),
    .N2MID(Tile_X1Y2_N2BEG),
    .N2END(Tile_X1Y2_N2BEGb),
    .N4END(Tile_X1Y2_N4BEG),
    .NN4END(Tile_X1Y2_NN4BEG),
    .Ci(Tile_X1Y2_Co),
    .E1END(Tile_X0Y1_E1BEG),
    .E2MID(Tile_X0Y1_E2BEG),
    .E2END(Tile_X0Y1_E2BEGb),
    .EE4END(Tile_X0Y1_EE4BEG),
    .E6END(Tile_X0Y1_E6BEG),
    .S1END(Tile_X1Y0_S1BEG),
    .S2MID(Tile_X1Y0_S2BEG),
    .S2END(Tile_X1Y0_S2BEGb),
    .S4END(Tile_X1Y0_S4BEG),
    .SS4END(Tile_X1Y0_SS4BEG),
    .W1END(Tile_X2Y1_W1BEG),
    .W2MID(Tile_X2Y1_W2BEG),
    .W2END(Tile_X2Y1_W2BEGb),
    .WW4END(Tile_X2Y1_WW4BEG),
    .W6END(Tile_X2Y1_W6BEG),
    .N1BEG(Tile_X1Y1_N1BEG),
    .N2BEG(Tile_X1Y1_N2BEG),
    .N2BEGb(Tile_X1Y1_N2BEGb),
    .N4BEG(Tile_X1Y1_N4BEG),
    .NN4BEG(Tile_X1Y1_NN4BEG),
    .Co(Tile_X1Y1_Co),
    .E1BEG(Tile_X1Y1_E1BEG),
    .E2BEG(Tile_X1Y1_E2BEG),
    .E2BEGb(Tile_X1Y1_E2BEGb),
    .EE4BEG(Tile_X1Y1_EE4BEG),
    .E6BEG(Tile_X1Y1_E6BEG),
    .S1BEG(Tile_X1Y1_S1BEG),
    .S2BEG(Tile_X1Y1_S2BEG),
    .S2BEGb(Tile_X1Y1_S2BEGb),
    .S4BEG(Tile_X1Y1_S4BEG),
    .SS4BEG(Tile_X1Y1_SS4BEG),
    .W1BEG(Tile_X1Y1_W1BEG),
    .W2BEG(Tile_X1Y1_W2BEG),
    .W2BEGb(Tile_X1Y1_W2BEGb),
    .WW4BEG(Tile_X1Y1_WW4BEG),
    .W6BEG(Tile_X1Y1_W6BEG),
    .UserCLK(Tile_X1Y2_UserCLKo),
    .UserCLKo(Tile_X1Y1_UserCLKo),
    .FrameData(Tile_X0Y1_FrameData_O),
    .FrameData_O(Tile_X1Y1_FrameData_O),
    .FrameStrobe(Tile_X1Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y1_Emulate_Bitstream)
    )
`endif
    Tile_X2Y1_LUT4AB
    (
    .N1END(Tile_X2Y2_N1BEG),
    .N2MID(Tile_X2Y2_N2BEG),
    .N2END(Tile_X2Y2_N2BEGb),
    .N4END(Tile_X2Y2_N4BEG),
    .NN4END(Tile_X2Y2_NN4BEG),
    .Ci(Tile_X2Y2_Co),
    .E1END(Tile_X1Y1_E1BEG),
    .E2MID(Tile_X1Y1_E2BEG),
    .E2END(Tile_X1Y1_E2BEGb),
    .EE4END(Tile_X1Y1_EE4BEG),
    .E6END(Tile_X1Y1_E6BEG),
    .S1END(Tile_X2Y0_S1BEG),
    .S2MID(Tile_X2Y0_S2BEG),
    .S2END(Tile_X2Y0_S2BEGb),
    .S4END(Tile_X2Y0_S4BEG),
    .SS4END(Tile_X2Y0_SS4BEG),
    .W1END(Tile_X3Y1_W1BEG),
    .W2MID(Tile_X3Y1_W2BEG),
    .W2END(Tile_X3Y1_W2BEGb),
    .WW4END(Tile_X3Y1_WW4BEG),
    .W6END(Tile_X3Y1_W6BEG),
    .N1BEG(Tile_X2Y1_N1BEG),
    .N2BEG(Tile_X2Y1_N2BEG),
    .N2BEGb(Tile_X2Y1_N2BEGb),
    .N4BEG(Tile_X2Y1_N4BEG),
    .NN4BEG(Tile_X2Y1_NN4BEG),
    .Co(Tile_X2Y1_Co),
    .E1BEG(Tile_X2Y1_E1BEG),
    .E2BEG(Tile_X2Y1_E2BEG),
    .E2BEGb(Tile_X2Y1_E2BEGb),
    .EE4BEG(Tile_X2Y1_EE4BEG),
    .E6BEG(Tile_X2Y1_E6BEG),
    .S1BEG(Tile_X2Y1_S1BEG),
    .S2BEG(Tile_X2Y1_S2BEG),
    .S2BEGb(Tile_X2Y1_S2BEGb),
    .S4BEG(Tile_X2Y1_S4BEG),
    .SS4BEG(Tile_X2Y1_SS4BEG),
    .W1BEG(Tile_X2Y1_W1BEG),
    .W2BEG(Tile_X2Y1_W2BEG),
    .W2BEGb(Tile_X2Y1_W2BEGb),
    .WW4BEG(Tile_X2Y1_WW4BEG),
    .W6BEG(Tile_X2Y1_W6BEG),
    .UserCLK(Tile_X2Y2_UserCLKo),
    .UserCLKo(Tile_X2Y1_UserCLKo),
    .FrameData(Tile_X1Y1_FrameData_O),
    .FrameData_O(Tile_X2Y1_FrameData_O),
    .FrameStrobe(Tile_X2Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y1_Emulate_Bitstream)
    )
`endif
    Tile_X3Y1_LUT4AB
    (
    .N1END(Tile_X3Y2_N1BEG),
    .N2MID(Tile_X3Y2_N2BEG),
    .N2END(Tile_X3Y2_N2BEGb),
    .N4END(Tile_X3Y2_N4BEG),
    .NN4END(Tile_X3Y2_NN4BEG),
    .Ci(Tile_X3Y2_Co),
    .E1END(Tile_X2Y1_E1BEG),
    .E2MID(Tile_X2Y1_E2BEG),
    .E2END(Tile_X2Y1_E2BEGb),
    .EE4END(Tile_X2Y1_EE4BEG),
    .E6END(Tile_X2Y1_E6BEG),
    .S1END(Tile_X3Y0_S1BEG),
    .S2MID(Tile_X3Y0_S2BEG),
    .S2END(Tile_X3Y0_S2BEGb),
    .S4END(Tile_X3Y0_S4BEG),
    .SS4END(Tile_X3Y0_SS4BEG),
    .W1END(Tile_X4Y1_W1BEG),
    .W2MID(Tile_X4Y1_W2BEG),
    .W2END(Tile_X4Y1_W2BEGb),
    .WW4END(Tile_X4Y1_WW4BEG),
    .W6END(Tile_X4Y1_W6BEG),
    .N1BEG(Tile_X3Y1_N1BEG),
    .N2BEG(Tile_X3Y1_N2BEG),
    .N2BEGb(Tile_X3Y1_N2BEGb),
    .N4BEG(Tile_X3Y1_N4BEG),
    .NN4BEG(Tile_X3Y1_NN4BEG),
    .Co(Tile_X3Y1_Co),
    .E1BEG(Tile_X3Y1_E1BEG),
    .E2BEG(Tile_X3Y1_E2BEG),
    .E2BEGb(Tile_X3Y1_E2BEGb),
    .EE4BEG(Tile_X3Y1_EE4BEG),
    .E6BEG(Tile_X3Y1_E6BEG),
    .S1BEG(Tile_X3Y1_S1BEG),
    .S2BEG(Tile_X3Y1_S2BEG),
    .S2BEGb(Tile_X3Y1_S2BEGb),
    .S4BEG(Tile_X3Y1_S4BEG),
    .SS4BEG(Tile_X3Y1_SS4BEG),
    .W1BEG(Tile_X3Y1_W1BEG),
    .W2BEG(Tile_X3Y1_W2BEG),
    .W2BEGb(Tile_X3Y1_W2BEGb),
    .WW4BEG(Tile_X3Y1_WW4BEG),
    .W6BEG(Tile_X3Y1_W6BEG),
    .UserCLK(Tile_X3Y2_UserCLKo),
    .UserCLKo(Tile_X3Y1_UserCLKo),
    .FrameData(Tile_X2Y1_FrameData_O),
    .FrameData_O(Tile_X3Y1_FrameData_O),
    .FrameStrobe(Tile_X3Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y1_Emulate_Bitstream)
    )
`endif
    Tile_X4Y1_LUT4AB
    (
    .N1END(Tile_X4Y2_N1BEG),
    .N2MID(Tile_X4Y2_N2BEG),
    .N2END(Tile_X4Y2_N2BEGb),
    .N4END(Tile_X4Y2_N4BEG),
    .NN4END(Tile_X4Y2_NN4BEG),
    .Ci(Tile_X4Y2_Co),
    .E1END(Tile_X3Y1_E1BEG),
    .E2MID(Tile_X3Y1_E2BEG),
    .E2END(Tile_X3Y1_E2BEGb),
    .EE4END(Tile_X3Y1_EE4BEG),
    .E6END(Tile_X3Y1_E6BEG),
    .S1END(Tile_X4Y0_S1BEG),
    .S2MID(Tile_X4Y0_S2BEG),
    .S2END(Tile_X4Y0_S2BEGb),
    .S4END(Tile_X4Y0_S4BEG),
    .SS4END(Tile_X4Y0_SS4BEG),
    .W1END(Tile_X5Y1_W1BEG),
    .W2MID(Tile_X5Y1_W2BEG),
    .W2END(Tile_X5Y1_W2BEGb),
    .WW4END(Tile_X5Y1_WW4BEG),
    .W6END(Tile_X5Y1_W6BEG),
    .N1BEG(Tile_X4Y1_N1BEG),
    .N2BEG(Tile_X4Y1_N2BEG),
    .N2BEGb(Tile_X4Y1_N2BEGb),
    .N4BEG(Tile_X4Y1_N4BEG),
    .NN4BEG(Tile_X4Y1_NN4BEG),
    .Co(Tile_X4Y1_Co),
    .E1BEG(Tile_X4Y1_E1BEG),
    .E2BEG(Tile_X4Y1_E2BEG),
    .E2BEGb(Tile_X4Y1_E2BEGb),
    .EE4BEG(Tile_X4Y1_EE4BEG),
    .E6BEG(Tile_X4Y1_E6BEG),
    .S1BEG(Tile_X4Y1_S1BEG),
    .S2BEG(Tile_X4Y1_S2BEG),
    .S2BEGb(Tile_X4Y1_S2BEGb),
    .S4BEG(Tile_X4Y1_S4BEG),
    .SS4BEG(Tile_X4Y1_SS4BEG),
    .W1BEG(Tile_X4Y1_W1BEG),
    .W2BEG(Tile_X4Y1_W2BEG),
    .W2BEGb(Tile_X4Y1_W2BEGb),
    .WW4BEG(Tile_X4Y1_WW4BEG),
    .W6BEG(Tile_X4Y1_W6BEG),
    .UserCLK(Tile_X4Y2_UserCLKo),
    .UserCLKo(Tile_X4Y1_UserCLKo),
    .FrameData(Tile_X3Y1_FrameData_O),
    .FrameData_O(Tile_X4Y1_FrameData_O),
    .FrameStrobe(Tile_X4Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y1_Emulate_Bitstream)
    )
`endif
    Tile_X5Y1_LUT4AB
    (
    .N1END(Tile_X5Y2_N1BEG),
    .N2MID(Tile_X5Y2_N2BEG),
    .N2END(Tile_X5Y2_N2BEGb),
    .N4END(Tile_X5Y2_N4BEG),
    .NN4END(Tile_X5Y2_NN4BEG),
    .Ci(Tile_X5Y2_Co),
    .E1END(Tile_X4Y1_E1BEG),
    .E2MID(Tile_X4Y1_E2BEG),
    .E2END(Tile_X4Y1_E2BEGb),
    .EE4END(Tile_X4Y1_EE4BEG),
    .E6END(Tile_X4Y1_E6BEG),
    .S1END(Tile_X5Y0_S1BEG),
    .S2MID(Tile_X5Y0_S2BEG),
    .S2END(Tile_X5Y0_S2BEGb),
    .S4END(Tile_X5Y0_S4BEG),
    .SS4END(Tile_X5Y0_SS4BEG),
    .W1END(Tile_X6Y1_W1BEG),
    .W2MID(Tile_X6Y1_W2BEG),
    .W2END(Tile_X6Y1_W2BEGb),
    .WW4END(Tile_X6Y1_WW4BEG),
    .W6END(Tile_X6Y1_W6BEG),
    .N1BEG(Tile_X5Y1_N1BEG),
    .N2BEG(Tile_X5Y1_N2BEG),
    .N2BEGb(Tile_X5Y1_N2BEGb),
    .N4BEG(Tile_X5Y1_N4BEG),
    .NN4BEG(Tile_X5Y1_NN4BEG),
    .Co(Tile_X5Y1_Co),
    .E1BEG(Tile_X5Y1_E1BEG),
    .E2BEG(Tile_X5Y1_E2BEG),
    .E2BEGb(Tile_X5Y1_E2BEGb),
    .EE4BEG(Tile_X5Y1_EE4BEG),
    .E6BEG(Tile_X5Y1_E6BEG),
    .S1BEG(Tile_X5Y1_S1BEG),
    .S2BEG(Tile_X5Y1_S2BEG),
    .S2BEGb(Tile_X5Y1_S2BEGb),
    .S4BEG(Tile_X5Y1_S4BEG),
    .SS4BEG(Tile_X5Y1_SS4BEG),
    .W1BEG(Tile_X5Y1_W1BEG),
    .W2BEG(Tile_X5Y1_W2BEG),
    .W2BEGb(Tile_X5Y1_W2BEGb),
    .WW4BEG(Tile_X5Y1_WW4BEG),
    .W6BEG(Tile_X5Y1_W6BEG),
    .UserCLK(Tile_X5Y2_UserCLKo),
    .UserCLKo(Tile_X5Y1_UserCLKo),
    .FrameData(Tile_X4Y1_FrameData_O),
    .FrameData_O(Tile_X5Y1_FrameData_O),
    .FrameStrobe(Tile_X5Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y1_Emulate_Bitstream)
    )
`endif
    Tile_X6Y1_LUT4AB
    (
    .N1END(Tile_X6Y2_N1BEG),
    .N2MID(Tile_X6Y2_N2BEG),
    .N2END(Tile_X6Y2_N2BEGb),
    .N4END(Tile_X6Y2_N4BEG),
    .NN4END(Tile_X6Y2_NN4BEG),
    .Ci(Tile_X6Y2_Co),
    .E1END(Tile_X5Y1_E1BEG),
    .E2MID(Tile_X5Y1_E2BEG),
    .E2END(Tile_X5Y1_E2BEGb),
    .EE4END(Tile_X5Y1_EE4BEG),
    .E6END(Tile_X5Y1_E6BEG),
    .S1END(Tile_X6Y0_S1BEG),
    .S2MID(Tile_X6Y0_S2BEG),
    .S2END(Tile_X6Y0_S2BEGb),
    .S4END(Tile_X6Y0_S4BEG),
    .SS4END(Tile_X6Y0_SS4BEG),
    .W1END(Tile_X7Y1_W1BEG),
    .W2MID(Tile_X7Y1_W2BEG),
    .W2END(Tile_X7Y1_W2BEGb),
    .WW4END(Tile_X7Y1_WW4BEG),
    .W6END(Tile_X7Y1_W6BEG),
    .N1BEG(Tile_X6Y1_N1BEG),
    .N2BEG(Tile_X6Y1_N2BEG),
    .N2BEGb(Tile_X6Y1_N2BEGb),
    .N4BEG(Tile_X6Y1_N4BEG),
    .NN4BEG(Tile_X6Y1_NN4BEG),
    .Co(Tile_X6Y1_Co),
    .E1BEG(Tile_X6Y1_E1BEG),
    .E2BEG(Tile_X6Y1_E2BEG),
    .E2BEGb(Tile_X6Y1_E2BEGb),
    .EE4BEG(Tile_X6Y1_EE4BEG),
    .E6BEG(Tile_X6Y1_E6BEG),
    .S1BEG(Tile_X6Y1_S1BEG),
    .S2BEG(Tile_X6Y1_S2BEG),
    .S2BEGb(Tile_X6Y1_S2BEGb),
    .S4BEG(Tile_X6Y1_S4BEG),
    .SS4BEG(Tile_X6Y1_SS4BEG),
    .W1BEG(Tile_X6Y1_W1BEG),
    .W2BEG(Tile_X6Y1_W2BEG),
    .W2BEGb(Tile_X6Y1_W2BEGb),
    .WW4BEG(Tile_X6Y1_WW4BEG),
    .W6BEG(Tile_X6Y1_W6BEG),
    .UserCLK(Tile_X6Y2_UserCLKo),
    .UserCLKo(Tile_X6Y1_UserCLKo),
    .FrameData(Tile_X5Y1_FrameData_O),
    .FrameData_O(Tile_X6Y1_FrameData_O),
    .FrameStrobe(Tile_X6Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y1_Emulate_Bitstream)
    )
`endif
    Tile_X7Y1_LUT4AB
    (
    .N1END(Tile_X7Y2_N1BEG),
    .N2MID(Tile_X7Y2_N2BEG),
    .N2END(Tile_X7Y2_N2BEGb),
    .N4END(Tile_X7Y2_N4BEG),
    .NN4END(Tile_X7Y2_NN4BEG),
    .Ci(Tile_X7Y2_Co),
    .E1END(Tile_X6Y1_E1BEG),
    .E2MID(Tile_X6Y1_E2BEG),
    .E2END(Tile_X6Y1_E2BEGb),
    .EE4END(Tile_X6Y1_EE4BEG),
    .E6END(Tile_X6Y1_E6BEG),
    .S1END(Tile_X7Y0_S1BEG),
    .S2MID(Tile_X7Y0_S2BEG),
    .S2END(Tile_X7Y0_S2BEGb),
    .S4END(Tile_X7Y0_S4BEG),
    .SS4END(Tile_X7Y0_SS4BEG),
    .W1END(Tile_X8Y1_W1BEG),
    .W2MID(Tile_X8Y1_W2BEG),
    .W2END(Tile_X8Y1_W2BEGb),
    .WW4END(Tile_X8Y1_WW4BEG),
    .W6END(Tile_X8Y1_W6BEG),
    .N1BEG(Tile_X7Y1_N1BEG),
    .N2BEG(Tile_X7Y1_N2BEG),
    .N2BEGb(Tile_X7Y1_N2BEGb),
    .N4BEG(Tile_X7Y1_N4BEG),
    .NN4BEG(Tile_X7Y1_NN4BEG),
    .Co(Tile_X7Y1_Co),
    .E1BEG(Tile_X7Y1_E1BEG),
    .E2BEG(Tile_X7Y1_E2BEG),
    .E2BEGb(Tile_X7Y1_E2BEGb),
    .EE4BEG(Tile_X7Y1_EE4BEG),
    .E6BEG(Tile_X7Y1_E6BEG),
    .S1BEG(Tile_X7Y1_S1BEG),
    .S2BEG(Tile_X7Y1_S2BEG),
    .S2BEGb(Tile_X7Y1_S2BEGb),
    .S4BEG(Tile_X7Y1_S4BEG),
    .SS4BEG(Tile_X7Y1_SS4BEG),
    .W1BEG(Tile_X7Y1_W1BEG),
    .W2BEG(Tile_X7Y1_W2BEG),
    .W2BEGb(Tile_X7Y1_W2BEGb),
    .WW4BEG(Tile_X7Y1_WW4BEG),
    .W6BEG(Tile_X7Y1_W6BEG),
    .UserCLK(Tile_X7Y2_UserCLKo),
    .UserCLKo(Tile_X7Y1_UserCLKo),
    .FrameData(Tile_X6Y1_FrameData_O),
    .FrameData_O(Tile_X7Y1_FrameData_O),
    .FrameStrobe(Tile_X7Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RAM_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y1_Emulate_Bitstream)
    )
`endif
    Tile_X8Y1_RAM_IO
    (
    .N1END(Tile_X8Y2_N1BEG),
    .N2MID(Tile_X8Y2_N2BEG),
    .N2END(Tile_X8Y2_N2BEGb),
    .N4END(Tile_X8Y2_N4BEG),
    .E1END(Tile_X7Y1_E1BEG),
    .E2MID(Tile_X7Y1_E2BEG),
    .E2END(Tile_X7Y1_E2BEGb),
    .EE4END(Tile_X7Y1_EE4BEG),
    .E6END(Tile_X7Y1_E6BEG),
    .S1END(Tile_X8Y0_S1BEG),
    .S2MID(Tile_X8Y0_S2BEG),
    .S2END(Tile_X8Y0_S2BEGb),
    .S4END(Tile_X8Y0_S4BEG),
    .N1BEG(Tile_X8Y1_N1BEG),
    .N2BEG(Tile_X8Y1_N2BEG),
    .N2BEGb(Tile_X8Y1_N2BEGb),
    .N4BEG(Tile_X8Y1_N4BEG),
    .S1BEG(Tile_X8Y1_S1BEG),
    .S2BEG(Tile_X8Y1_S2BEG),
    .S2BEGb(Tile_X8Y1_S2BEGb),
    .S4BEG(Tile_X8Y1_S4BEG),
    .W1BEG(Tile_X8Y1_W1BEG),
    .W2BEG(Tile_X8Y1_W2BEG),
    .W2BEGb(Tile_X8Y1_W2BEGb),
    .WW4BEG(Tile_X8Y1_WW4BEG),
    .W6BEG(Tile_X8Y1_W6BEG),
    .RAM2FAB_D0_I0(Tile_X8Y1_RAM2FAB_D0_I0),
    .RAM2FAB_D0_I1(Tile_X8Y1_RAM2FAB_D0_I1),
    .RAM2FAB_D0_I2(Tile_X8Y1_RAM2FAB_D0_I2),
    .RAM2FAB_D0_I3(Tile_X8Y1_RAM2FAB_D0_I3),
    .RAM2FAB_D1_I0(Tile_X8Y1_RAM2FAB_D1_I0),
    .RAM2FAB_D1_I1(Tile_X8Y1_RAM2FAB_D1_I1),
    .RAM2FAB_D1_I2(Tile_X8Y1_RAM2FAB_D1_I2),
    .RAM2FAB_D1_I3(Tile_X8Y1_RAM2FAB_D1_I3),
    .RAM2FAB_D2_I0(Tile_X8Y1_RAM2FAB_D2_I0),
    .RAM2FAB_D2_I1(Tile_X8Y1_RAM2FAB_D2_I1),
    .RAM2FAB_D2_I2(Tile_X8Y1_RAM2FAB_D2_I2),
    .RAM2FAB_D2_I3(Tile_X8Y1_RAM2FAB_D2_I3),
    .RAM2FAB_D3_I0(Tile_X8Y1_RAM2FAB_D3_I0),
    .RAM2FAB_D3_I1(Tile_X8Y1_RAM2FAB_D3_I1),
    .RAM2FAB_D3_I2(Tile_X8Y1_RAM2FAB_D3_I2),
    .RAM2FAB_D3_I3(Tile_X8Y1_RAM2FAB_D3_I3),
    .FAB2RAM_D0_O0(Tile_X8Y1_FAB2RAM_D0_O0),
    .FAB2RAM_D0_O1(Tile_X8Y1_FAB2RAM_D0_O1),
    .FAB2RAM_D0_O2(Tile_X8Y1_FAB2RAM_D0_O2),
    .FAB2RAM_D0_O3(Tile_X8Y1_FAB2RAM_D0_O3),
    .FAB2RAM_D1_O0(Tile_X8Y1_FAB2RAM_D1_O0),
    .FAB2RAM_D1_O1(Tile_X8Y1_FAB2RAM_D1_O1),
    .FAB2RAM_D1_O2(Tile_X8Y1_FAB2RAM_D1_O2),
    .FAB2RAM_D1_O3(Tile_X8Y1_FAB2RAM_D1_O3),
    .FAB2RAM_D2_O0(Tile_X8Y1_FAB2RAM_D2_O0),
    .FAB2RAM_D2_O1(Tile_X8Y1_FAB2RAM_D2_O1),
    .FAB2RAM_D2_O2(Tile_X8Y1_FAB2RAM_D2_O2),
    .FAB2RAM_D2_O3(Tile_X8Y1_FAB2RAM_D2_O3),
    .FAB2RAM_D3_O0(Tile_X8Y1_FAB2RAM_D3_O0),
    .FAB2RAM_D3_O1(Tile_X8Y1_FAB2RAM_D3_O1),
    .FAB2RAM_D3_O2(Tile_X8Y1_FAB2RAM_D3_O2),
    .FAB2RAM_D3_O3(Tile_X8Y1_FAB2RAM_D3_O3),
    .FAB2RAM_A0_O0(Tile_X8Y1_FAB2RAM_A0_O0),
    .FAB2RAM_A0_O1(Tile_X8Y1_FAB2RAM_A0_O1),
    .FAB2RAM_A0_O2(Tile_X8Y1_FAB2RAM_A0_O2),
    .FAB2RAM_A0_O3(Tile_X8Y1_FAB2RAM_A0_O3),
    .FAB2RAM_A1_O0(Tile_X8Y1_FAB2RAM_A1_O0),
    .FAB2RAM_A1_O1(Tile_X8Y1_FAB2RAM_A1_O1),
    .FAB2RAM_A1_O2(Tile_X8Y1_FAB2RAM_A1_O2),
    .FAB2RAM_A1_O3(Tile_X8Y1_FAB2RAM_A1_O3),
    .FAB2RAM_C_O0(Tile_X8Y1_FAB2RAM_C_O0),
    .FAB2RAM_C_O1(Tile_X8Y1_FAB2RAM_C_O1),
    .FAB2RAM_C_O2(Tile_X8Y1_FAB2RAM_C_O2),
    .FAB2RAM_C_O3(Tile_X8Y1_FAB2RAM_C_O3),
    .Config_accessC_bit0(Tile_X8Y1_Config_accessC_bit0),
    .Config_accessC_bit1(Tile_X8Y1_Config_accessC_bit1),
    .Config_accessC_bit2(Tile_X8Y1_Config_accessC_bit2),
    .Config_accessC_bit3(Tile_X8Y1_Config_accessC_bit3),
    .UserCLK(Tile_X8Y2_UserCLKo),
    .UserCLKo(Tile_X8Y1_UserCLKo),
    .FrameData(Tile_X7Y1_FrameData_O),
    .FrameData_O(Tile_X8Y1_FrameData_O),
    .FrameStrobe(Tile_X8Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y2_Emulate_Bitstream)
    )
`endif
    Tile_X0Y2_W_IO
    (
    .W1END(Tile_X1Y2_W1BEG),
    .W2MID(Tile_X1Y2_W2BEG),
    .W2END(Tile_X1Y2_W2BEGb),
    .WW4END(Tile_X1Y2_WW4BEG),
    .W6END(Tile_X1Y2_W6BEG),
    .E1BEG(Tile_X0Y2_E1BEG),
    .E2BEG(Tile_X0Y2_E2BEG),
    .E2BEGb(Tile_X0Y2_E2BEGb),
    .EE4BEG(Tile_X0Y2_EE4BEG),
    .E6BEG(Tile_X0Y2_E6BEG),
    .A_O_top(Tile_X0Y2_A_O_top),
    .A_I_top(Tile_X0Y2_A_I_top),
    .A_T_top(Tile_X0Y2_A_T_top),
    .B_O_top(Tile_X0Y2_B_O_top),
    .B_I_top(Tile_X0Y2_B_I_top),
    .B_T_top(Tile_X0Y2_B_T_top),
    .A_config_C_bit0(Tile_X0Y2_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y2_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y2_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y2_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y2_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y2_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y2_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y2_B_config_C_bit3),
    .UserCLK(Tile_X0Y3_UserCLKo),
    .UserCLKo(Tile_X0Y2_UserCLKo),
    .FrameData(Tile_Y2_FrameData),
    .FrameData_O(Tile_X0Y2_FrameData_O),
    .FrameStrobe(Tile_X0Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y2_Emulate_Bitstream)
    )
`endif
    Tile_X1Y2_LUT4AB
    (
    .N1END(Tile_X1Y3_N1BEG),
    .N2MID(Tile_X1Y3_N2BEG),
    .N2END(Tile_X1Y3_N2BEGb),
    .N4END(Tile_X1Y3_N4BEG),
    .NN4END(Tile_X1Y3_NN4BEG),
    .Ci(Tile_X1Y3_Co),
    .E1END(Tile_X0Y2_E1BEG),
    .E2MID(Tile_X0Y2_E2BEG),
    .E2END(Tile_X0Y2_E2BEGb),
    .EE4END(Tile_X0Y2_EE4BEG),
    .E6END(Tile_X0Y2_E6BEG),
    .S1END(Tile_X1Y1_S1BEG),
    .S2MID(Tile_X1Y1_S2BEG),
    .S2END(Tile_X1Y1_S2BEGb),
    .S4END(Tile_X1Y1_S4BEG),
    .SS4END(Tile_X1Y1_SS4BEG),
    .W1END(Tile_X2Y2_W1BEG),
    .W2MID(Tile_X2Y2_W2BEG),
    .W2END(Tile_X2Y2_W2BEGb),
    .WW4END(Tile_X2Y2_WW4BEG),
    .W6END(Tile_X2Y2_W6BEG),
    .N1BEG(Tile_X1Y2_N1BEG),
    .N2BEG(Tile_X1Y2_N2BEG),
    .N2BEGb(Tile_X1Y2_N2BEGb),
    .N4BEG(Tile_X1Y2_N4BEG),
    .NN4BEG(Tile_X1Y2_NN4BEG),
    .Co(Tile_X1Y2_Co),
    .E1BEG(Tile_X1Y2_E1BEG),
    .E2BEG(Tile_X1Y2_E2BEG),
    .E2BEGb(Tile_X1Y2_E2BEGb),
    .EE4BEG(Tile_X1Y2_EE4BEG),
    .E6BEG(Tile_X1Y2_E6BEG),
    .S1BEG(Tile_X1Y2_S1BEG),
    .S2BEG(Tile_X1Y2_S2BEG),
    .S2BEGb(Tile_X1Y2_S2BEGb),
    .S4BEG(Tile_X1Y2_S4BEG),
    .SS4BEG(Tile_X1Y2_SS4BEG),
    .W1BEG(Tile_X1Y2_W1BEG),
    .W2BEG(Tile_X1Y2_W2BEG),
    .W2BEGb(Tile_X1Y2_W2BEGb),
    .WW4BEG(Tile_X1Y2_WW4BEG),
    .W6BEG(Tile_X1Y2_W6BEG),
    .UserCLK(Tile_X1Y3_UserCLKo),
    .UserCLKo(Tile_X1Y2_UserCLKo),
    .FrameData(Tile_X0Y2_FrameData_O),
    .FrameData_O(Tile_X1Y2_FrameData_O),
    .FrameStrobe(Tile_X1Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y2_Emulate_Bitstream)
    )
`endif
    Tile_X2Y2_LUT4AB
    (
    .N1END(Tile_X2Y3_N1BEG),
    .N2MID(Tile_X2Y3_N2BEG),
    .N2END(Tile_X2Y3_N2BEGb),
    .N4END(Tile_X2Y3_N4BEG),
    .NN4END(Tile_X2Y3_NN4BEG),
    .Ci(Tile_X2Y3_Co),
    .E1END(Tile_X1Y2_E1BEG),
    .E2MID(Tile_X1Y2_E2BEG),
    .E2END(Tile_X1Y2_E2BEGb),
    .EE4END(Tile_X1Y2_EE4BEG),
    .E6END(Tile_X1Y2_E6BEG),
    .S1END(Tile_X2Y1_S1BEG),
    .S2MID(Tile_X2Y1_S2BEG),
    .S2END(Tile_X2Y1_S2BEGb),
    .S4END(Tile_X2Y1_S4BEG),
    .SS4END(Tile_X2Y1_SS4BEG),
    .W1END(Tile_X3Y2_W1BEG),
    .W2MID(Tile_X3Y2_W2BEG),
    .W2END(Tile_X3Y2_W2BEGb),
    .WW4END(Tile_X3Y2_WW4BEG),
    .W6END(Tile_X3Y2_W6BEG),
    .N1BEG(Tile_X2Y2_N1BEG),
    .N2BEG(Tile_X2Y2_N2BEG),
    .N2BEGb(Tile_X2Y2_N2BEGb),
    .N4BEG(Tile_X2Y2_N4BEG),
    .NN4BEG(Tile_X2Y2_NN4BEG),
    .Co(Tile_X2Y2_Co),
    .E1BEG(Tile_X2Y2_E1BEG),
    .E2BEG(Tile_X2Y2_E2BEG),
    .E2BEGb(Tile_X2Y2_E2BEGb),
    .EE4BEG(Tile_X2Y2_EE4BEG),
    .E6BEG(Tile_X2Y2_E6BEG),
    .S1BEG(Tile_X2Y2_S1BEG),
    .S2BEG(Tile_X2Y2_S2BEG),
    .S2BEGb(Tile_X2Y2_S2BEGb),
    .S4BEG(Tile_X2Y2_S4BEG),
    .SS4BEG(Tile_X2Y2_SS4BEG),
    .W1BEG(Tile_X2Y2_W1BEG),
    .W2BEG(Tile_X2Y2_W2BEG),
    .W2BEGb(Tile_X2Y2_W2BEGb),
    .WW4BEG(Tile_X2Y2_WW4BEG),
    .W6BEG(Tile_X2Y2_W6BEG),
    .UserCLK(Tile_X2Y3_UserCLKo),
    .UserCLKo(Tile_X2Y2_UserCLKo),
    .FrameData(Tile_X1Y2_FrameData_O),
    .FrameData_O(Tile_X2Y2_FrameData_O),
    .FrameStrobe(Tile_X2Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y2_Emulate_Bitstream)
    )
`endif
    Tile_X3Y2_LUT4AB
    (
    .N1END(Tile_X3Y3_N1BEG),
    .N2MID(Tile_X3Y3_N2BEG),
    .N2END(Tile_X3Y3_N2BEGb),
    .N4END(Tile_X3Y3_N4BEG),
    .NN4END(Tile_X3Y3_NN4BEG),
    .Ci(Tile_X3Y3_Co),
    .E1END(Tile_X2Y2_E1BEG),
    .E2MID(Tile_X2Y2_E2BEG),
    .E2END(Tile_X2Y2_E2BEGb),
    .EE4END(Tile_X2Y2_EE4BEG),
    .E6END(Tile_X2Y2_E6BEG),
    .S1END(Tile_X3Y1_S1BEG),
    .S2MID(Tile_X3Y1_S2BEG),
    .S2END(Tile_X3Y1_S2BEGb),
    .S4END(Tile_X3Y1_S4BEG),
    .SS4END(Tile_X3Y1_SS4BEG),
    .W1END(Tile_X4Y2_W1BEG),
    .W2MID(Tile_X4Y2_W2BEG),
    .W2END(Tile_X4Y2_W2BEGb),
    .WW4END(Tile_X4Y2_WW4BEG),
    .W6END(Tile_X4Y2_W6BEG),
    .N1BEG(Tile_X3Y2_N1BEG),
    .N2BEG(Tile_X3Y2_N2BEG),
    .N2BEGb(Tile_X3Y2_N2BEGb),
    .N4BEG(Tile_X3Y2_N4BEG),
    .NN4BEG(Tile_X3Y2_NN4BEG),
    .Co(Tile_X3Y2_Co),
    .E1BEG(Tile_X3Y2_E1BEG),
    .E2BEG(Tile_X3Y2_E2BEG),
    .E2BEGb(Tile_X3Y2_E2BEGb),
    .EE4BEG(Tile_X3Y2_EE4BEG),
    .E6BEG(Tile_X3Y2_E6BEG),
    .S1BEG(Tile_X3Y2_S1BEG),
    .S2BEG(Tile_X3Y2_S2BEG),
    .S2BEGb(Tile_X3Y2_S2BEGb),
    .S4BEG(Tile_X3Y2_S4BEG),
    .SS4BEG(Tile_X3Y2_SS4BEG),
    .W1BEG(Tile_X3Y2_W1BEG),
    .W2BEG(Tile_X3Y2_W2BEG),
    .W2BEGb(Tile_X3Y2_W2BEGb),
    .WW4BEG(Tile_X3Y2_WW4BEG),
    .W6BEG(Tile_X3Y2_W6BEG),
    .UserCLK(Tile_X3Y3_UserCLKo),
    .UserCLKo(Tile_X3Y2_UserCLKo),
    .FrameData(Tile_X2Y2_FrameData_O),
    .FrameData_O(Tile_X3Y2_FrameData_O),
    .FrameStrobe(Tile_X3Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y2_Emulate_Bitstream)
    )
`endif
    Tile_X4Y2_LUT4AB
    (
    .N1END(Tile_X4Y3_N1BEG),
    .N2MID(Tile_X4Y3_N2BEG),
    .N2END(Tile_X4Y3_N2BEGb),
    .N4END(Tile_X4Y3_N4BEG),
    .NN4END(Tile_X4Y3_NN4BEG),
    .Ci(Tile_X4Y3_Co),
    .E1END(Tile_X3Y2_E1BEG),
    .E2MID(Tile_X3Y2_E2BEG),
    .E2END(Tile_X3Y2_E2BEGb),
    .EE4END(Tile_X3Y2_EE4BEG),
    .E6END(Tile_X3Y2_E6BEG),
    .S1END(Tile_X4Y1_S1BEG),
    .S2MID(Tile_X4Y1_S2BEG),
    .S2END(Tile_X4Y1_S2BEGb),
    .S4END(Tile_X4Y1_S4BEG),
    .SS4END(Tile_X4Y1_SS4BEG),
    .W1END(Tile_X5Y2_W1BEG),
    .W2MID(Tile_X5Y2_W2BEG),
    .W2END(Tile_X5Y2_W2BEGb),
    .WW4END(Tile_X5Y2_WW4BEG),
    .W6END(Tile_X5Y2_W6BEG),
    .N1BEG(Tile_X4Y2_N1BEG),
    .N2BEG(Tile_X4Y2_N2BEG),
    .N2BEGb(Tile_X4Y2_N2BEGb),
    .N4BEG(Tile_X4Y2_N4BEG),
    .NN4BEG(Tile_X4Y2_NN4BEG),
    .Co(Tile_X4Y2_Co),
    .E1BEG(Tile_X4Y2_E1BEG),
    .E2BEG(Tile_X4Y2_E2BEG),
    .E2BEGb(Tile_X4Y2_E2BEGb),
    .EE4BEG(Tile_X4Y2_EE4BEG),
    .E6BEG(Tile_X4Y2_E6BEG),
    .S1BEG(Tile_X4Y2_S1BEG),
    .S2BEG(Tile_X4Y2_S2BEG),
    .S2BEGb(Tile_X4Y2_S2BEGb),
    .S4BEG(Tile_X4Y2_S4BEG),
    .SS4BEG(Tile_X4Y2_SS4BEG),
    .W1BEG(Tile_X4Y2_W1BEG),
    .W2BEG(Tile_X4Y2_W2BEG),
    .W2BEGb(Tile_X4Y2_W2BEGb),
    .WW4BEG(Tile_X4Y2_WW4BEG),
    .W6BEG(Tile_X4Y2_W6BEG),
    .UserCLK(Tile_X4Y3_UserCLKo),
    .UserCLKo(Tile_X4Y2_UserCLKo),
    .FrameData(Tile_X3Y2_FrameData_O),
    .FrameData_O(Tile_X4Y2_FrameData_O),
    .FrameStrobe(Tile_X4Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y2_Emulate_Bitstream)
    )
`endif
    Tile_X5Y2_LUT4AB
    (
    .N1END(Tile_X5Y3_N1BEG),
    .N2MID(Tile_X5Y3_N2BEG),
    .N2END(Tile_X5Y3_N2BEGb),
    .N4END(Tile_X5Y3_N4BEG),
    .NN4END(Tile_X5Y3_NN4BEG),
    .Ci(Tile_X5Y3_Co),
    .E1END(Tile_X4Y2_E1BEG),
    .E2MID(Tile_X4Y2_E2BEG),
    .E2END(Tile_X4Y2_E2BEGb),
    .EE4END(Tile_X4Y2_EE4BEG),
    .E6END(Tile_X4Y2_E6BEG),
    .S1END(Tile_X5Y1_S1BEG),
    .S2MID(Tile_X5Y1_S2BEG),
    .S2END(Tile_X5Y1_S2BEGb),
    .S4END(Tile_X5Y1_S4BEG),
    .SS4END(Tile_X5Y1_SS4BEG),
    .W1END(Tile_X6Y2_W1BEG),
    .W2MID(Tile_X6Y2_W2BEG),
    .W2END(Tile_X6Y2_W2BEGb),
    .WW4END(Tile_X6Y2_WW4BEG),
    .W6END(Tile_X6Y2_W6BEG),
    .N1BEG(Tile_X5Y2_N1BEG),
    .N2BEG(Tile_X5Y2_N2BEG),
    .N2BEGb(Tile_X5Y2_N2BEGb),
    .N4BEG(Tile_X5Y2_N4BEG),
    .NN4BEG(Tile_X5Y2_NN4BEG),
    .Co(Tile_X5Y2_Co),
    .E1BEG(Tile_X5Y2_E1BEG),
    .E2BEG(Tile_X5Y2_E2BEG),
    .E2BEGb(Tile_X5Y2_E2BEGb),
    .EE4BEG(Tile_X5Y2_EE4BEG),
    .E6BEG(Tile_X5Y2_E6BEG),
    .S1BEG(Tile_X5Y2_S1BEG),
    .S2BEG(Tile_X5Y2_S2BEG),
    .S2BEGb(Tile_X5Y2_S2BEGb),
    .S4BEG(Tile_X5Y2_S4BEG),
    .SS4BEG(Tile_X5Y2_SS4BEG),
    .W1BEG(Tile_X5Y2_W1BEG),
    .W2BEG(Tile_X5Y2_W2BEG),
    .W2BEGb(Tile_X5Y2_W2BEGb),
    .WW4BEG(Tile_X5Y2_WW4BEG),
    .W6BEG(Tile_X5Y2_W6BEG),
    .UserCLK(Tile_X5Y3_UserCLKo),
    .UserCLKo(Tile_X5Y2_UserCLKo),
    .FrameData(Tile_X4Y2_FrameData_O),
    .FrameData_O(Tile_X5Y2_FrameData_O),
    .FrameStrobe(Tile_X5Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y2_Emulate_Bitstream)
    )
`endif
    Tile_X6Y2_LUT4AB
    (
    .N1END(Tile_X6Y3_N1BEG),
    .N2MID(Tile_X6Y3_N2BEG),
    .N2END(Tile_X6Y3_N2BEGb),
    .N4END(Tile_X6Y3_N4BEG),
    .NN4END(Tile_X6Y3_NN4BEG),
    .Ci(Tile_X6Y3_Co),
    .E1END(Tile_X5Y2_E1BEG),
    .E2MID(Tile_X5Y2_E2BEG),
    .E2END(Tile_X5Y2_E2BEGb),
    .EE4END(Tile_X5Y2_EE4BEG),
    .E6END(Tile_X5Y2_E6BEG),
    .S1END(Tile_X6Y1_S1BEG),
    .S2MID(Tile_X6Y1_S2BEG),
    .S2END(Tile_X6Y1_S2BEGb),
    .S4END(Tile_X6Y1_S4BEG),
    .SS4END(Tile_X6Y1_SS4BEG),
    .W1END(Tile_X7Y2_W1BEG),
    .W2MID(Tile_X7Y2_W2BEG),
    .W2END(Tile_X7Y2_W2BEGb),
    .WW4END(Tile_X7Y2_WW4BEG),
    .W6END(Tile_X7Y2_W6BEG),
    .N1BEG(Tile_X6Y2_N1BEG),
    .N2BEG(Tile_X6Y2_N2BEG),
    .N2BEGb(Tile_X6Y2_N2BEGb),
    .N4BEG(Tile_X6Y2_N4BEG),
    .NN4BEG(Tile_X6Y2_NN4BEG),
    .Co(Tile_X6Y2_Co),
    .E1BEG(Tile_X6Y2_E1BEG),
    .E2BEG(Tile_X6Y2_E2BEG),
    .E2BEGb(Tile_X6Y2_E2BEGb),
    .EE4BEG(Tile_X6Y2_EE4BEG),
    .E6BEG(Tile_X6Y2_E6BEG),
    .S1BEG(Tile_X6Y2_S1BEG),
    .S2BEG(Tile_X6Y2_S2BEG),
    .S2BEGb(Tile_X6Y2_S2BEGb),
    .S4BEG(Tile_X6Y2_S4BEG),
    .SS4BEG(Tile_X6Y2_SS4BEG),
    .W1BEG(Tile_X6Y2_W1BEG),
    .W2BEG(Tile_X6Y2_W2BEG),
    .W2BEGb(Tile_X6Y2_W2BEGb),
    .WW4BEG(Tile_X6Y2_WW4BEG),
    .W6BEG(Tile_X6Y2_W6BEG),
    .UserCLK(Tile_X6Y3_UserCLKo),
    .UserCLKo(Tile_X6Y2_UserCLKo),
    .FrameData(Tile_X5Y2_FrameData_O),
    .FrameData_O(Tile_X6Y2_FrameData_O),
    .FrameStrobe(Tile_X6Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y2_Emulate_Bitstream)
    )
`endif
    Tile_X7Y2_LUT4AB
    (
    .N1END(Tile_X7Y3_N1BEG),
    .N2MID(Tile_X7Y3_N2BEG),
    .N2END(Tile_X7Y3_N2BEGb),
    .N4END(Tile_X7Y3_N4BEG),
    .NN4END(Tile_X7Y3_NN4BEG),
    .Ci(Tile_X7Y3_Co),
    .E1END(Tile_X6Y2_E1BEG),
    .E2MID(Tile_X6Y2_E2BEG),
    .E2END(Tile_X6Y2_E2BEGb),
    .EE4END(Tile_X6Y2_EE4BEG),
    .E6END(Tile_X6Y2_E6BEG),
    .S1END(Tile_X7Y1_S1BEG),
    .S2MID(Tile_X7Y1_S2BEG),
    .S2END(Tile_X7Y1_S2BEGb),
    .S4END(Tile_X7Y1_S4BEG),
    .SS4END(Tile_X7Y1_SS4BEG),
    .W1END(Tile_X8Y2_W1BEG),
    .W2MID(Tile_X8Y2_W2BEG),
    .W2END(Tile_X8Y2_W2BEGb),
    .WW4END(Tile_X8Y2_WW4BEG),
    .W6END(Tile_X8Y2_W6BEG),
    .N1BEG(Tile_X7Y2_N1BEG),
    .N2BEG(Tile_X7Y2_N2BEG),
    .N2BEGb(Tile_X7Y2_N2BEGb),
    .N4BEG(Tile_X7Y2_N4BEG),
    .NN4BEG(Tile_X7Y2_NN4BEG),
    .Co(Tile_X7Y2_Co),
    .E1BEG(Tile_X7Y2_E1BEG),
    .E2BEG(Tile_X7Y2_E2BEG),
    .E2BEGb(Tile_X7Y2_E2BEGb),
    .EE4BEG(Tile_X7Y2_EE4BEG),
    .E6BEG(Tile_X7Y2_E6BEG),
    .S1BEG(Tile_X7Y2_S1BEG),
    .S2BEG(Tile_X7Y2_S2BEG),
    .S2BEGb(Tile_X7Y2_S2BEGb),
    .S4BEG(Tile_X7Y2_S4BEG),
    .SS4BEG(Tile_X7Y2_SS4BEG),
    .W1BEG(Tile_X7Y2_W1BEG),
    .W2BEG(Tile_X7Y2_W2BEG),
    .W2BEGb(Tile_X7Y2_W2BEGb),
    .WW4BEG(Tile_X7Y2_WW4BEG),
    .W6BEG(Tile_X7Y2_W6BEG),
    .UserCLK(Tile_X7Y3_UserCLKo),
    .UserCLKo(Tile_X7Y2_UserCLKo),
    .FrameData(Tile_X6Y2_FrameData_O),
    .FrameData_O(Tile_X7Y2_FrameData_O),
    .FrameStrobe(Tile_X7Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RAM_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y2_Emulate_Bitstream)
    )
`endif
    Tile_X8Y2_RAM_IO
    (
    .N1END(Tile_X8Y3_N1BEG),
    .N2MID(Tile_X8Y3_N2BEG),
    .N2END(Tile_X8Y3_N2BEGb),
    .N4END(Tile_X8Y3_N4BEG),
    .E1END(Tile_X7Y2_E1BEG),
    .E2MID(Tile_X7Y2_E2BEG),
    .E2END(Tile_X7Y2_E2BEGb),
    .EE4END(Tile_X7Y2_EE4BEG),
    .E6END(Tile_X7Y2_E6BEG),
    .S1END(Tile_X8Y1_S1BEG),
    .S2MID(Tile_X8Y1_S2BEG),
    .S2END(Tile_X8Y1_S2BEGb),
    .S4END(Tile_X8Y1_S4BEG),
    .N1BEG(Tile_X8Y2_N1BEG),
    .N2BEG(Tile_X8Y2_N2BEG),
    .N2BEGb(Tile_X8Y2_N2BEGb),
    .N4BEG(Tile_X8Y2_N4BEG),
    .S1BEG(Tile_X8Y2_S1BEG),
    .S2BEG(Tile_X8Y2_S2BEG),
    .S2BEGb(Tile_X8Y2_S2BEGb),
    .S4BEG(Tile_X8Y2_S4BEG),
    .W1BEG(Tile_X8Y2_W1BEG),
    .W2BEG(Tile_X8Y2_W2BEG),
    .W2BEGb(Tile_X8Y2_W2BEGb),
    .WW4BEG(Tile_X8Y2_WW4BEG),
    .W6BEG(Tile_X8Y2_W6BEG),
    .RAM2FAB_D0_I0(Tile_X8Y2_RAM2FAB_D0_I0),
    .RAM2FAB_D0_I1(Tile_X8Y2_RAM2FAB_D0_I1),
    .RAM2FAB_D0_I2(Tile_X8Y2_RAM2FAB_D0_I2),
    .RAM2FAB_D0_I3(Tile_X8Y2_RAM2FAB_D0_I3),
    .RAM2FAB_D1_I0(Tile_X8Y2_RAM2FAB_D1_I0),
    .RAM2FAB_D1_I1(Tile_X8Y2_RAM2FAB_D1_I1),
    .RAM2FAB_D1_I2(Tile_X8Y2_RAM2FAB_D1_I2),
    .RAM2FAB_D1_I3(Tile_X8Y2_RAM2FAB_D1_I3),
    .RAM2FAB_D2_I0(Tile_X8Y2_RAM2FAB_D2_I0),
    .RAM2FAB_D2_I1(Tile_X8Y2_RAM2FAB_D2_I1),
    .RAM2FAB_D2_I2(Tile_X8Y2_RAM2FAB_D2_I2),
    .RAM2FAB_D2_I3(Tile_X8Y2_RAM2FAB_D2_I3),
    .RAM2FAB_D3_I0(Tile_X8Y2_RAM2FAB_D3_I0),
    .RAM2FAB_D3_I1(Tile_X8Y2_RAM2FAB_D3_I1),
    .RAM2FAB_D3_I2(Tile_X8Y2_RAM2FAB_D3_I2),
    .RAM2FAB_D3_I3(Tile_X8Y2_RAM2FAB_D3_I3),
    .FAB2RAM_D0_O0(Tile_X8Y2_FAB2RAM_D0_O0),
    .FAB2RAM_D0_O1(Tile_X8Y2_FAB2RAM_D0_O1),
    .FAB2RAM_D0_O2(Tile_X8Y2_FAB2RAM_D0_O2),
    .FAB2RAM_D0_O3(Tile_X8Y2_FAB2RAM_D0_O3),
    .FAB2RAM_D1_O0(Tile_X8Y2_FAB2RAM_D1_O0),
    .FAB2RAM_D1_O1(Tile_X8Y2_FAB2RAM_D1_O1),
    .FAB2RAM_D1_O2(Tile_X8Y2_FAB2RAM_D1_O2),
    .FAB2RAM_D1_O3(Tile_X8Y2_FAB2RAM_D1_O3),
    .FAB2RAM_D2_O0(Tile_X8Y2_FAB2RAM_D2_O0),
    .FAB2RAM_D2_O1(Tile_X8Y2_FAB2RAM_D2_O1),
    .FAB2RAM_D2_O2(Tile_X8Y2_FAB2RAM_D2_O2),
    .FAB2RAM_D2_O3(Tile_X8Y2_FAB2RAM_D2_O3),
    .FAB2RAM_D3_O0(Tile_X8Y2_FAB2RAM_D3_O0),
    .FAB2RAM_D3_O1(Tile_X8Y2_FAB2RAM_D3_O1),
    .FAB2RAM_D3_O2(Tile_X8Y2_FAB2RAM_D3_O2),
    .FAB2RAM_D3_O3(Tile_X8Y2_FAB2RAM_D3_O3),
    .FAB2RAM_A0_O0(Tile_X8Y2_FAB2RAM_A0_O0),
    .FAB2RAM_A0_O1(Tile_X8Y2_FAB2RAM_A0_O1),
    .FAB2RAM_A0_O2(Tile_X8Y2_FAB2RAM_A0_O2),
    .FAB2RAM_A0_O3(Tile_X8Y2_FAB2RAM_A0_O3),
    .FAB2RAM_A1_O0(Tile_X8Y2_FAB2RAM_A1_O0),
    .FAB2RAM_A1_O1(Tile_X8Y2_FAB2RAM_A1_O1),
    .FAB2RAM_A1_O2(Tile_X8Y2_FAB2RAM_A1_O2),
    .FAB2RAM_A1_O3(Tile_X8Y2_FAB2RAM_A1_O3),
    .FAB2RAM_C_O0(Tile_X8Y2_FAB2RAM_C_O0),
    .FAB2RAM_C_O1(Tile_X8Y2_FAB2RAM_C_O1),
    .FAB2RAM_C_O2(Tile_X8Y2_FAB2RAM_C_O2),
    .FAB2RAM_C_O3(Tile_X8Y2_FAB2RAM_C_O3),
    .Config_accessC_bit0(Tile_X8Y2_Config_accessC_bit0),
    .Config_accessC_bit1(Tile_X8Y2_Config_accessC_bit1),
    .Config_accessC_bit2(Tile_X8Y2_Config_accessC_bit2),
    .Config_accessC_bit3(Tile_X8Y2_Config_accessC_bit3),
    .UserCLK(Tile_X8Y3_UserCLKo),
    .UserCLKo(Tile_X8Y2_UserCLKo),
    .FrameData(Tile_X7Y2_FrameData_O),
    .FrameData_O(Tile_X8Y2_FrameData_O),
    .FrameStrobe(Tile_X8Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y3_Emulate_Bitstream)
    )
`endif
    Tile_X0Y3_W_IO
    (
    .W1END(Tile_X1Y3_W1BEG),
    .W2MID(Tile_X1Y3_W2BEG),
    .W2END(Tile_X1Y3_W2BEGb),
    .WW4END(Tile_X1Y3_WW4BEG),
    .W6END(Tile_X1Y3_W6BEG),
    .E1BEG(Tile_X0Y3_E1BEG),
    .E2BEG(Tile_X0Y3_E2BEG),
    .E2BEGb(Tile_X0Y3_E2BEGb),
    .EE4BEG(Tile_X0Y3_EE4BEG),
    .E6BEG(Tile_X0Y3_E6BEG),
    .A_O_top(Tile_X0Y3_A_O_top),
    .A_I_top(Tile_X0Y3_A_I_top),
    .A_T_top(Tile_X0Y3_A_T_top),
    .B_O_top(Tile_X0Y3_B_O_top),
    .B_I_top(Tile_X0Y3_B_I_top),
    .B_T_top(Tile_X0Y3_B_T_top),
    .A_config_C_bit0(Tile_X0Y3_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y3_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y3_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y3_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y3_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y3_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y3_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y3_B_config_C_bit3),
    .UserCLK(Tile_X0Y4_UserCLKo),
    .UserCLKo(Tile_X0Y3_UserCLKo),
    .FrameData(Tile_Y3_FrameData),
    .FrameData_O(Tile_X0Y3_FrameData_O),
    .FrameStrobe(Tile_X0Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y3_Emulate_Bitstream)
    )
`endif
    Tile_X1Y3_LUT4AB
    (
    .N1END(Tile_X1Y4_N1BEG),
    .N2MID(Tile_X1Y4_N2BEG),
    .N2END(Tile_X1Y4_N2BEGb),
    .N4END(Tile_X1Y4_N4BEG),
    .NN4END(Tile_X1Y4_NN4BEG),
    .Ci(Tile_X1Y4_Co),
    .E1END(Tile_X0Y3_E1BEG),
    .E2MID(Tile_X0Y3_E2BEG),
    .E2END(Tile_X0Y3_E2BEGb),
    .EE4END(Tile_X0Y3_EE4BEG),
    .E6END(Tile_X0Y3_E6BEG),
    .S1END(Tile_X1Y2_S1BEG),
    .S2MID(Tile_X1Y2_S2BEG),
    .S2END(Tile_X1Y2_S2BEGb),
    .S4END(Tile_X1Y2_S4BEG),
    .SS4END(Tile_X1Y2_SS4BEG),
    .W1END(Tile_X2Y3_W1BEG),
    .W2MID(Tile_X2Y3_W2BEG),
    .W2END(Tile_X2Y3_W2BEGb),
    .WW4END(Tile_X2Y3_WW4BEG),
    .W6END(Tile_X2Y3_W6BEG),
    .N1BEG(Tile_X1Y3_N1BEG),
    .N2BEG(Tile_X1Y3_N2BEG),
    .N2BEGb(Tile_X1Y3_N2BEGb),
    .N4BEG(Tile_X1Y3_N4BEG),
    .NN4BEG(Tile_X1Y3_NN4BEG),
    .Co(Tile_X1Y3_Co),
    .E1BEG(Tile_X1Y3_E1BEG),
    .E2BEG(Tile_X1Y3_E2BEG),
    .E2BEGb(Tile_X1Y3_E2BEGb),
    .EE4BEG(Tile_X1Y3_EE4BEG),
    .E6BEG(Tile_X1Y3_E6BEG),
    .S1BEG(Tile_X1Y3_S1BEG),
    .S2BEG(Tile_X1Y3_S2BEG),
    .S2BEGb(Tile_X1Y3_S2BEGb),
    .S4BEG(Tile_X1Y3_S4BEG),
    .SS4BEG(Tile_X1Y3_SS4BEG),
    .W1BEG(Tile_X1Y3_W1BEG),
    .W2BEG(Tile_X1Y3_W2BEG),
    .W2BEGb(Tile_X1Y3_W2BEGb),
    .WW4BEG(Tile_X1Y3_WW4BEG),
    .W6BEG(Tile_X1Y3_W6BEG),
    .UserCLK(Tile_X1Y4_UserCLKo),
    .UserCLKo(Tile_X1Y3_UserCLKo),
    .FrameData(Tile_X0Y3_FrameData_O),
    .FrameData_O(Tile_X1Y3_FrameData_O),
    .FrameStrobe(Tile_X1Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y3_Emulate_Bitstream)
    )
`endif
    Tile_X2Y3_LUT4AB
    (
    .N1END(Tile_X2Y4_N1BEG),
    .N2MID(Tile_X2Y4_N2BEG),
    .N2END(Tile_X2Y4_N2BEGb),
    .N4END(Tile_X2Y4_N4BEG),
    .NN4END(Tile_X2Y4_NN4BEG),
    .Ci(Tile_X2Y4_Co),
    .E1END(Tile_X1Y3_E1BEG),
    .E2MID(Tile_X1Y3_E2BEG),
    .E2END(Tile_X1Y3_E2BEGb),
    .EE4END(Tile_X1Y3_EE4BEG),
    .E6END(Tile_X1Y3_E6BEG),
    .S1END(Tile_X2Y2_S1BEG),
    .S2MID(Tile_X2Y2_S2BEG),
    .S2END(Tile_X2Y2_S2BEGb),
    .S4END(Tile_X2Y2_S4BEG),
    .SS4END(Tile_X2Y2_SS4BEG),
    .W1END(Tile_X3Y3_W1BEG),
    .W2MID(Tile_X3Y3_W2BEG),
    .W2END(Tile_X3Y3_W2BEGb),
    .WW4END(Tile_X3Y3_WW4BEG),
    .W6END(Tile_X3Y3_W6BEG),
    .N1BEG(Tile_X2Y3_N1BEG),
    .N2BEG(Tile_X2Y3_N2BEG),
    .N2BEGb(Tile_X2Y3_N2BEGb),
    .N4BEG(Tile_X2Y3_N4BEG),
    .NN4BEG(Tile_X2Y3_NN4BEG),
    .Co(Tile_X2Y3_Co),
    .E1BEG(Tile_X2Y3_E1BEG),
    .E2BEG(Tile_X2Y3_E2BEG),
    .E2BEGb(Tile_X2Y3_E2BEGb),
    .EE4BEG(Tile_X2Y3_EE4BEG),
    .E6BEG(Tile_X2Y3_E6BEG),
    .S1BEG(Tile_X2Y3_S1BEG),
    .S2BEG(Tile_X2Y3_S2BEG),
    .S2BEGb(Tile_X2Y3_S2BEGb),
    .S4BEG(Tile_X2Y3_S4BEG),
    .SS4BEG(Tile_X2Y3_SS4BEG),
    .W1BEG(Tile_X2Y3_W1BEG),
    .W2BEG(Tile_X2Y3_W2BEG),
    .W2BEGb(Tile_X2Y3_W2BEGb),
    .WW4BEG(Tile_X2Y3_WW4BEG),
    .W6BEG(Tile_X2Y3_W6BEG),
    .UserCLK(Tile_X2Y4_UserCLKo),
    .UserCLKo(Tile_X2Y3_UserCLKo),
    .FrameData(Tile_X1Y3_FrameData_O),
    .FrameData_O(Tile_X2Y3_FrameData_O),
    .FrameStrobe(Tile_X2Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y3_Emulate_Bitstream)
    )
`endif
    Tile_X3Y3_LUT4AB
    (
    .N1END(Tile_X3Y4_N1BEG),
    .N2MID(Tile_X3Y4_N2BEG),
    .N2END(Tile_X3Y4_N2BEGb),
    .N4END(Tile_X3Y4_N4BEG),
    .NN4END(Tile_X3Y4_NN4BEG),
    .Ci(Tile_X3Y4_Co),
    .E1END(Tile_X2Y3_E1BEG),
    .E2MID(Tile_X2Y3_E2BEG),
    .E2END(Tile_X2Y3_E2BEGb),
    .EE4END(Tile_X2Y3_EE4BEG),
    .E6END(Tile_X2Y3_E6BEG),
    .S1END(Tile_X3Y2_S1BEG),
    .S2MID(Tile_X3Y2_S2BEG),
    .S2END(Tile_X3Y2_S2BEGb),
    .S4END(Tile_X3Y2_S4BEG),
    .SS4END(Tile_X3Y2_SS4BEG),
    .W1END(Tile_X4Y3_W1BEG),
    .W2MID(Tile_X4Y3_W2BEG),
    .W2END(Tile_X4Y3_W2BEGb),
    .WW4END(Tile_X4Y3_WW4BEG),
    .W6END(Tile_X4Y3_W6BEG),
    .N1BEG(Tile_X3Y3_N1BEG),
    .N2BEG(Tile_X3Y3_N2BEG),
    .N2BEGb(Tile_X3Y3_N2BEGb),
    .N4BEG(Tile_X3Y3_N4BEG),
    .NN4BEG(Tile_X3Y3_NN4BEG),
    .Co(Tile_X3Y3_Co),
    .E1BEG(Tile_X3Y3_E1BEG),
    .E2BEG(Tile_X3Y3_E2BEG),
    .E2BEGb(Tile_X3Y3_E2BEGb),
    .EE4BEG(Tile_X3Y3_EE4BEG),
    .E6BEG(Tile_X3Y3_E6BEG),
    .S1BEG(Tile_X3Y3_S1BEG),
    .S2BEG(Tile_X3Y3_S2BEG),
    .S2BEGb(Tile_X3Y3_S2BEGb),
    .S4BEG(Tile_X3Y3_S4BEG),
    .SS4BEG(Tile_X3Y3_SS4BEG),
    .W1BEG(Tile_X3Y3_W1BEG),
    .W2BEG(Tile_X3Y3_W2BEG),
    .W2BEGb(Tile_X3Y3_W2BEGb),
    .WW4BEG(Tile_X3Y3_WW4BEG),
    .W6BEG(Tile_X3Y3_W6BEG),
    .UserCLK(Tile_X3Y4_UserCLKo),
    .UserCLKo(Tile_X3Y3_UserCLKo),
    .FrameData(Tile_X2Y3_FrameData_O),
    .FrameData_O(Tile_X3Y3_FrameData_O),
    .FrameStrobe(Tile_X3Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y3_Emulate_Bitstream)
    )
`endif
    Tile_X4Y3_LUT4AB
    (
    .N1END(Tile_X4Y4_N1BEG),
    .N2MID(Tile_X4Y4_N2BEG),
    .N2END(Tile_X4Y4_N2BEGb),
    .N4END(Tile_X4Y4_N4BEG),
    .NN4END(Tile_X4Y4_NN4BEG),
    .Ci(Tile_X4Y4_Co),
    .E1END(Tile_X3Y3_E1BEG),
    .E2MID(Tile_X3Y3_E2BEG),
    .E2END(Tile_X3Y3_E2BEGb),
    .EE4END(Tile_X3Y3_EE4BEG),
    .E6END(Tile_X3Y3_E6BEG),
    .S1END(Tile_X4Y2_S1BEG),
    .S2MID(Tile_X4Y2_S2BEG),
    .S2END(Tile_X4Y2_S2BEGb),
    .S4END(Tile_X4Y2_S4BEG),
    .SS4END(Tile_X4Y2_SS4BEG),
    .W1END(Tile_X5Y3_W1BEG),
    .W2MID(Tile_X5Y3_W2BEG),
    .W2END(Tile_X5Y3_W2BEGb),
    .WW4END(Tile_X5Y3_WW4BEG),
    .W6END(Tile_X5Y3_W6BEG),
    .N1BEG(Tile_X4Y3_N1BEG),
    .N2BEG(Tile_X4Y3_N2BEG),
    .N2BEGb(Tile_X4Y3_N2BEGb),
    .N4BEG(Tile_X4Y3_N4BEG),
    .NN4BEG(Tile_X4Y3_NN4BEG),
    .Co(Tile_X4Y3_Co),
    .E1BEG(Tile_X4Y3_E1BEG),
    .E2BEG(Tile_X4Y3_E2BEG),
    .E2BEGb(Tile_X4Y3_E2BEGb),
    .EE4BEG(Tile_X4Y3_EE4BEG),
    .E6BEG(Tile_X4Y3_E6BEG),
    .S1BEG(Tile_X4Y3_S1BEG),
    .S2BEG(Tile_X4Y3_S2BEG),
    .S2BEGb(Tile_X4Y3_S2BEGb),
    .S4BEG(Tile_X4Y3_S4BEG),
    .SS4BEG(Tile_X4Y3_SS4BEG),
    .W1BEG(Tile_X4Y3_W1BEG),
    .W2BEG(Tile_X4Y3_W2BEG),
    .W2BEGb(Tile_X4Y3_W2BEGb),
    .WW4BEG(Tile_X4Y3_WW4BEG),
    .W6BEG(Tile_X4Y3_W6BEG),
    .UserCLK(Tile_X4Y4_UserCLKo),
    .UserCLKo(Tile_X4Y3_UserCLKo),
    .FrameData(Tile_X3Y3_FrameData_O),
    .FrameData_O(Tile_X4Y3_FrameData_O),
    .FrameStrobe(Tile_X4Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y3_Emulate_Bitstream)
    )
`endif
    Tile_X5Y3_LUT4AB
    (
    .N1END(Tile_X5Y4_N1BEG),
    .N2MID(Tile_X5Y4_N2BEG),
    .N2END(Tile_X5Y4_N2BEGb),
    .N4END(Tile_X5Y4_N4BEG),
    .NN4END(Tile_X5Y4_NN4BEG),
    .Ci(Tile_X5Y4_Co),
    .E1END(Tile_X4Y3_E1BEG),
    .E2MID(Tile_X4Y3_E2BEG),
    .E2END(Tile_X4Y3_E2BEGb),
    .EE4END(Tile_X4Y3_EE4BEG),
    .E6END(Tile_X4Y3_E6BEG),
    .S1END(Tile_X5Y2_S1BEG),
    .S2MID(Tile_X5Y2_S2BEG),
    .S2END(Tile_X5Y2_S2BEGb),
    .S4END(Tile_X5Y2_S4BEG),
    .SS4END(Tile_X5Y2_SS4BEG),
    .W1END(Tile_X6Y3_W1BEG),
    .W2MID(Tile_X6Y3_W2BEG),
    .W2END(Tile_X6Y3_W2BEGb),
    .WW4END(Tile_X6Y3_WW4BEG),
    .W6END(Tile_X6Y3_W6BEG),
    .N1BEG(Tile_X5Y3_N1BEG),
    .N2BEG(Tile_X5Y3_N2BEG),
    .N2BEGb(Tile_X5Y3_N2BEGb),
    .N4BEG(Tile_X5Y3_N4BEG),
    .NN4BEG(Tile_X5Y3_NN4BEG),
    .Co(Tile_X5Y3_Co),
    .E1BEG(Tile_X5Y3_E1BEG),
    .E2BEG(Tile_X5Y3_E2BEG),
    .E2BEGb(Tile_X5Y3_E2BEGb),
    .EE4BEG(Tile_X5Y3_EE4BEG),
    .E6BEG(Tile_X5Y3_E6BEG),
    .S1BEG(Tile_X5Y3_S1BEG),
    .S2BEG(Tile_X5Y3_S2BEG),
    .S2BEGb(Tile_X5Y3_S2BEGb),
    .S4BEG(Tile_X5Y3_S4BEG),
    .SS4BEG(Tile_X5Y3_SS4BEG),
    .W1BEG(Tile_X5Y3_W1BEG),
    .W2BEG(Tile_X5Y3_W2BEG),
    .W2BEGb(Tile_X5Y3_W2BEGb),
    .WW4BEG(Tile_X5Y3_WW4BEG),
    .W6BEG(Tile_X5Y3_W6BEG),
    .UserCLK(Tile_X5Y4_UserCLKo),
    .UserCLKo(Tile_X5Y3_UserCLKo),
    .FrameData(Tile_X4Y3_FrameData_O),
    .FrameData_O(Tile_X5Y3_FrameData_O),
    .FrameStrobe(Tile_X5Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y3_Emulate_Bitstream)
    )
`endif
    Tile_X6Y3_LUT4AB
    (
    .N1END(Tile_X6Y4_N1BEG),
    .N2MID(Tile_X6Y4_N2BEG),
    .N2END(Tile_X6Y4_N2BEGb),
    .N4END(Tile_X6Y4_N4BEG),
    .NN4END(Tile_X6Y4_NN4BEG),
    .Ci(Tile_X6Y4_Co),
    .E1END(Tile_X5Y3_E1BEG),
    .E2MID(Tile_X5Y3_E2BEG),
    .E2END(Tile_X5Y3_E2BEGb),
    .EE4END(Tile_X5Y3_EE4BEG),
    .E6END(Tile_X5Y3_E6BEG),
    .S1END(Tile_X6Y2_S1BEG),
    .S2MID(Tile_X6Y2_S2BEG),
    .S2END(Tile_X6Y2_S2BEGb),
    .S4END(Tile_X6Y2_S4BEG),
    .SS4END(Tile_X6Y2_SS4BEG),
    .W1END(Tile_X7Y3_W1BEG),
    .W2MID(Tile_X7Y3_W2BEG),
    .W2END(Tile_X7Y3_W2BEGb),
    .WW4END(Tile_X7Y3_WW4BEG),
    .W6END(Tile_X7Y3_W6BEG),
    .N1BEG(Tile_X6Y3_N1BEG),
    .N2BEG(Tile_X6Y3_N2BEG),
    .N2BEGb(Tile_X6Y3_N2BEGb),
    .N4BEG(Tile_X6Y3_N4BEG),
    .NN4BEG(Tile_X6Y3_NN4BEG),
    .Co(Tile_X6Y3_Co),
    .E1BEG(Tile_X6Y3_E1BEG),
    .E2BEG(Tile_X6Y3_E2BEG),
    .E2BEGb(Tile_X6Y3_E2BEGb),
    .EE4BEG(Tile_X6Y3_EE4BEG),
    .E6BEG(Tile_X6Y3_E6BEG),
    .S1BEG(Tile_X6Y3_S1BEG),
    .S2BEG(Tile_X6Y3_S2BEG),
    .S2BEGb(Tile_X6Y3_S2BEGb),
    .S4BEG(Tile_X6Y3_S4BEG),
    .SS4BEG(Tile_X6Y3_SS4BEG),
    .W1BEG(Tile_X6Y3_W1BEG),
    .W2BEG(Tile_X6Y3_W2BEG),
    .W2BEGb(Tile_X6Y3_W2BEGb),
    .WW4BEG(Tile_X6Y3_WW4BEG),
    .W6BEG(Tile_X6Y3_W6BEG),
    .UserCLK(Tile_X6Y4_UserCLKo),
    .UserCLKo(Tile_X6Y3_UserCLKo),
    .FrameData(Tile_X5Y3_FrameData_O),
    .FrameData_O(Tile_X6Y3_FrameData_O),
    .FrameStrobe(Tile_X6Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y3_Emulate_Bitstream)
    )
`endif
    Tile_X7Y3_LUT4AB
    (
    .N1END(Tile_X7Y4_N1BEG),
    .N2MID(Tile_X7Y4_N2BEG),
    .N2END(Tile_X7Y4_N2BEGb),
    .N4END(Tile_X7Y4_N4BEG),
    .NN4END(Tile_X7Y4_NN4BEG),
    .Ci(Tile_X7Y4_Co),
    .E1END(Tile_X6Y3_E1BEG),
    .E2MID(Tile_X6Y3_E2BEG),
    .E2END(Tile_X6Y3_E2BEGb),
    .EE4END(Tile_X6Y3_EE4BEG),
    .E6END(Tile_X6Y3_E6BEG),
    .S1END(Tile_X7Y2_S1BEG),
    .S2MID(Tile_X7Y2_S2BEG),
    .S2END(Tile_X7Y2_S2BEGb),
    .S4END(Tile_X7Y2_S4BEG),
    .SS4END(Tile_X7Y2_SS4BEG),
    .W1END(Tile_X8Y3_W1BEG),
    .W2MID(Tile_X8Y3_W2BEG),
    .W2END(Tile_X8Y3_W2BEGb),
    .WW4END(Tile_X8Y3_WW4BEG),
    .W6END(Tile_X8Y3_W6BEG),
    .N1BEG(Tile_X7Y3_N1BEG),
    .N2BEG(Tile_X7Y3_N2BEG),
    .N2BEGb(Tile_X7Y3_N2BEGb),
    .N4BEG(Tile_X7Y3_N4BEG),
    .NN4BEG(Tile_X7Y3_NN4BEG),
    .Co(Tile_X7Y3_Co),
    .E1BEG(Tile_X7Y3_E1BEG),
    .E2BEG(Tile_X7Y3_E2BEG),
    .E2BEGb(Tile_X7Y3_E2BEGb),
    .EE4BEG(Tile_X7Y3_EE4BEG),
    .E6BEG(Tile_X7Y3_E6BEG),
    .S1BEG(Tile_X7Y3_S1BEG),
    .S2BEG(Tile_X7Y3_S2BEG),
    .S2BEGb(Tile_X7Y3_S2BEGb),
    .S4BEG(Tile_X7Y3_S4BEG),
    .SS4BEG(Tile_X7Y3_SS4BEG),
    .W1BEG(Tile_X7Y3_W1BEG),
    .W2BEG(Tile_X7Y3_W2BEG),
    .W2BEGb(Tile_X7Y3_W2BEGb),
    .WW4BEG(Tile_X7Y3_WW4BEG),
    .W6BEG(Tile_X7Y3_W6BEG),
    .UserCLK(Tile_X7Y4_UserCLKo),
    .UserCLKo(Tile_X7Y3_UserCLKo),
    .FrameData(Tile_X6Y3_FrameData_O),
    .FrameData_O(Tile_X7Y3_FrameData_O),
    .FrameStrobe(Tile_X7Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RAM_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y3_Emulate_Bitstream)
    )
`endif
    Tile_X8Y3_RAM_IO
    (
    .N1END(Tile_X8Y4_N1BEG),
    .N2MID(Tile_X8Y4_N2BEG),
    .N2END(Tile_X8Y4_N2BEGb),
    .N4END(Tile_X8Y4_N4BEG),
    .E1END(Tile_X7Y3_E1BEG),
    .E2MID(Tile_X7Y3_E2BEG),
    .E2END(Tile_X7Y3_E2BEGb),
    .EE4END(Tile_X7Y3_EE4BEG),
    .E6END(Tile_X7Y3_E6BEG),
    .S1END(Tile_X8Y2_S1BEG),
    .S2MID(Tile_X8Y2_S2BEG),
    .S2END(Tile_X8Y2_S2BEGb),
    .S4END(Tile_X8Y2_S4BEG),
    .N1BEG(Tile_X8Y3_N1BEG),
    .N2BEG(Tile_X8Y3_N2BEG),
    .N2BEGb(Tile_X8Y3_N2BEGb),
    .N4BEG(Tile_X8Y3_N4BEG),
    .S1BEG(Tile_X8Y3_S1BEG),
    .S2BEG(Tile_X8Y3_S2BEG),
    .S2BEGb(Tile_X8Y3_S2BEGb),
    .S4BEG(Tile_X8Y3_S4BEG),
    .W1BEG(Tile_X8Y3_W1BEG),
    .W2BEG(Tile_X8Y3_W2BEG),
    .W2BEGb(Tile_X8Y3_W2BEGb),
    .WW4BEG(Tile_X8Y3_WW4BEG),
    .W6BEG(Tile_X8Y3_W6BEG),
    .RAM2FAB_D0_I0(Tile_X8Y3_RAM2FAB_D0_I0),
    .RAM2FAB_D0_I1(Tile_X8Y3_RAM2FAB_D0_I1),
    .RAM2FAB_D0_I2(Tile_X8Y3_RAM2FAB_D0_I2),
    .RAM2FAB_D0_I3(Tile_X8Y3_RAM2FAB_D0_I3),
    .RAM2FAB_D1_I0(Tile_X8Y3_RAM2FAB_D1_I0),
    .RAM2FAB_D1_I1(Tile_X8Y3_RAM2FAB_D1_I1),
    .RAM2FAB_D1_I2(Tile_X8Y3_RAM2FAB_D1_I2),
    .RAM2FAB_D1_I3(Tile_X8Y3_RAM2FAB_D1_I3),
    .RAM2FAB_D2_I0(Tile_X8Y3_RAM2FAB_D2_I0),
    .RAM2FAB_D2_I1(Tile_X8Y3_RAM2FAB_D2_I1),
    .RAM2FAB_D2_I2(Tile_X8Y3_RAM2FAB_D2_I2),
    .RAM2FAB_D2_I3(Tile_X8Y3_RAM2FAB_D2_I3),
    .RAM2FAB_D3_I0(Tile_X8Y3_RAM2FAB_D3_I0),
    .RAM2FAB_D3_I1(Tile_X8Y3_RAM2FAB_D3_I1),
    .RAM2FAB_D3_I2(Tile_X8Y3_RAM2FAB_D3_I2),
    .RAM2FAB_D3_I3(Tile_X8Y3_RAM2FAB_D3_I3),
    .FAB2RAM_D0_O0(Tile_X8Y3_FAB2RAM_D0_O0),
    .FAB2RAM_D0_O1(Tile_X8Y3_FAB2RAM_D0_O1),
    .FAB2RAM_D0_O2(Tile_X8Y3_FAB2RAM_D0_O2),
    .FAB2RAM_D0_O3(Tile_X8Y3_FAB2RAM_D0_O3),
    .FAB2RAM_D1_O0(Tile_X8Y3_FAB2RAM_D1_O0),
    .FAB2RAM_D1_O1(Tile_X8Y3_FAB2RAM_D1_O1),
    .FAB2RAM_D1_O2(Tile_X8Y3_FAB2RAM_D1_O2),
    .FAB2RAM_D1_O3(Tile_X8Y3_FAB2RAM_D1_O3),
    .FAB2RAM_D2_O0(Tile_X8Y3_FAB2RAM_D2_O0),
    .FAB2RAM_D2_O1(Tile_X8Y3_FAB2RAM_D2_O1),
    .FAB2RAM_D2_O2(Tile_X8Y3_FAB2RAM_D2_O2),
    .FAB2RAM_D2_O3(Tile_X8Y3_FAB2RAM_D2_O3),
    .FAB2RAM_D3_O0(Tile_X8Y3_FAB2RAM_D3_O0),
    .FAB2RAM_D3_O1(Tile_X8Y3_FAB2RAM_D3_O1),
    .FAB2RAM_D3_O2(Tile_X8Y3_FAB2RAM_D3_O2),
    .FAB2RAM_D3_O3(Tile_X8Y3_FAB2RAM_D3_O3),
    .FAB2RAM_A0_O0(Tile_X8Y3_FAB2RAM_A0_O0),
    .FAB2RAM_A0_O1(Tile_X8Y3_FAB2RAM_A0_O1),
    .FAB2RAM_A0_O2(Tile_X8Y3_FAB2RAM_A0_O2),
    .FAB2RAM_A0_O3(Tile_X8Y3_FAB2RAM_A0_O3),
    .FAB2RAM_A1_O0(Tile_X8Y3_FAB2RAM_A1_O0),
    .FAB2RAM_A1_O1(Tile_X8Y3_FAB2RAM_A1_O1),
    .FAB2RAM_A1_O2(Tile_X8Y3_FAB2RAM_A1_O2),
    .FAB2RAM_A1_O3(Tile_X8Y3_FAB2RAM_A1_O3),
    .FAB2RAM_C_O0(Tile_X8Y3_FAB2RAM_C_O0),
    .FAB2RAM_C_O1(Tile_X8Y3_FAB2RAM_C_O1),
    .FAB2RAM_C_O2(Tile_X8Y3_FAB2RAM_C_O2),
    .FAB2RAM_C_O3(Tile_X8Y3_FAB2RAM_C_O3),
    .Config_accessC_bit0(Tile_X8Y3_Config_accessC_bit0),
    .Config_accessC_bit1(Tile_X8Y3_Config_accessC_bit1),
    .Config_accessC_bit2(Tile_X8Y3_Config_accessC_bit2),
    .Config_accessC_bit3(Tile_X8Y3_Config_accessC_bit3),
    .UserCLK(Tile_X8Y4_UserCLKo),
    .UserCLKo(Tile_X8Y3_UserCLKo),
    .FrameData(Tile_X7Y3_FrameData_O),
    .FrameData_O(Tile_X8Y3_FrameData_O),
    .FrameStrobe(Tile_X8Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y4_Emulate_Bitstream)
    )
`endif
    Tile_X0Y4_W_IO
    (
    .W1END(Tile_X1Y4_W1BEG),
    .W2MID(Tile_X1Y4_W2BEG),
    .W2END(Tile_X1Y4_W2BEGb),
    .WW4END(Tile_X1Y4_WW4BEG),
    .W6END(Tile_X1Y4_W6BEG),
    .E1BEG(Tile_X0Y4_E1BEG),
    .E2BEG(Tile_X0Y4_E2BEG),
    .E2BEGb(Tile_X0Y4_E2BEGb),
    .EE4BEG(Tile_X0Y4_EE4BEG),
    .E6BEG(Tile_X0Y4_E6BEG),
    .A_O_top(Tile_X0Y4_A_O_top),
    .A_I_top(Tile_X0Y4_A_I_top),
    .A_T_top(Tile_X0Y4_A_T_top),
    .B_O_top(Tile_X0Y4_B_O_top),
    .B_I_top(Tile_X0Y4_B_I_top),
    .B_T_top(Tile_X0Y4_B_T_top),
    .A_config_C_bit0(Tile_X0Y4_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y4_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y4_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y4_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y4_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y4_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y4_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y4_B_config_C_bit3),
    .UserCLK(Tile_X0Y5_UserCLKo),
    .UserCLKo(Tile_X0Y4_UserCLKo),
    .FrameData(Tile_Y4_FrameData),
    .FrameData_O(Tile_X0Y4_FrameData_O),
    .FrameStrobe(Tile_X0Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y4_Emulate_Bitstream)
    )
`endif
    Tile_X1Y4_LUT4AB
    (
    .N1END(Tile_X1Y5_N1BEG),
    .N2MID(Tile_X1Y5_N2BEG),
    .N2END(Tile_X1Y5_N2BEGb),
    .N4END(Tile_X1Y5_N4BEG),
    .NN4END(Tile_X1Y5_NN4BEG),
    .Ci(Tile_X1Y5_Co),
    .E1END(Tile_X0Y4_E1BEG),
    .E2MID(Tile_X0Y4_E2BEG),
    .E2END(Tile_X0Y4_E2BEGb),
    .EE4END(Tile_X0Y4_EE4BEG),
    .E6END(Tile_X0Y4_E6BEG),
    .S1END(Tile_X1Y3_S1BEG),
    .S2MID(Tile_X1Y3_S2BEG),
    .S2END(Tile_X1Y3_S2BEGb),
    .S4END(Tile_X1Y3_S4BEG),
    .SS4END(Tile_X1Y3_SS4BEG),
    .W1END(Tile_X2Y4_W1BEG),
    .W2MID(Tile_X2Y4_W2BEG),
    .W2END(Tile_X2Y4_W2BEGb),
    .WW4END(Tile_X2Y4_WW4BEG),
    .W6END(Tile_X2Y4_W6BEG),
    .N1BEG(Tile_X1Y4_N1BEG),
    .N2BEG(Tile_X1Y4_N2BEG),
    .N2BEGb(Tile_X1Y4_N2BEGb),
    .N4BEG(Tile_X1Y4_N4BEG),
    .NN4BEG(Tile_X1Y4_NN4BEG),
    .Co(Tile_X1Y4_Co),
    .E1BEG(Tile_X1Y4_E1BEG),
    .E2BEG(Tile_X1Y4_E2BEG),
    .E2BEGb(Tile_X1Y4_E2BEGb),
    .EE4BEG(Tile_X1Y4_EE4BEG),
    .E6BEG(Tile_X1Y4_E6BEG),
    .S1BEG(Tile_X1Y4_S1BEG),
    .S2BEG(Tile_X1Y4_S2BEG),
    .S2BEGb(Tile_X1Y4_S2BEGb),
    .S4BEG(Tile_X1Y4_S4BEG),
    .SS4BEG(Tile_X1Y4_SS4BEG),
    .W1BEG(Tile_X1Y4_W1BEG),
    .W2BEG(Tile_X1Y4_W2BEG),
    .W2BEGb(Tile_X1Y4_W2BEGb),
    .WW4BEG(Tile_X1Y4_WW4BEG),
    .W6BEG(Tile_X1Y4_W6BEG),
    .UserCLK(Tile_X1Y5_UserCLKo),
    .UserCLKo(Tile_X1Y4_UserCLKo),
    .FrameData(Tile_X0Y4_FrameData_O),
    .FrameData_O(Tile_X1Y4_FrameData_O),
    .FrameStrobe(Tile_X1Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y4_Emulate_Bitstream)
    )
`endif
    Tile_X2Y4_LUT4AB
    (
    .N1END(Tile_X2Y5_N1BEG),
    .N2MID(Tile_X2Y5_N2BEG),
    .N2END(Tile_X2Y5_N2BEGb),
    .N4END(Tile_X2Y5_N4BEG),
    .NN4END(Tile_X2Y5_NN4BEG),
    .Ci(Tile_X2Y5_Co),
    .E1END(Tile_X1Y4_E1BEG),
    .E2MID(Tile_X1Y4_E2BEG),
    .E2END(Tile_X1Y4_E2BEGb),
    .EE4END(Tile_X1Y4_EE4BEG),
    .E6END(Tile_X1Y4_E6BEG),
    .S1END(Tile_X2Y3_S1BEG),
    .S2MID(Tile_X2Y3_S2BEG),
    .S2END(Tile_X2Y3_S2BEGb),
    .S4END(Tile_X2Y3_S4BEG),
    .SS4END(Tile_X2Y3_SS4BEG),
    .W1END(Tile_X3Y4_W1BEG),
    .W2MID(Tile_X3Y4_W2BEG),
    .W2END(Tile_X3Y4_W2BEGb),
    .WW4END(Tile_X3Y4_WW4BEG),
    .W6END(Tile_X3Y4_W6BEG),
    .N1BEG(Tile_X2Y4_N1BEG),
    .N2BEG(Tile_X2Y4_N2BEG),
    .N2BEGb(Tile_X2Y4_N2BEGb),
    .N4BEG(Tile_X2Y4_N4BEG),
    .NN4BEG(Tile_X2Y4_NN4BEG),
    .Co(Tile_X2Y4_Co),
    .E1BEG(Tile_X2Y4_E1BEG),
    .E2BEG(Tile_X2Y4_E2BEG),
    .E2BEGb(Tile_X2Y4_E2BEGb),
    .EE4BEG(Tile_X2Y4_EE4BEG),
    .E6BEG(Tile_X2Y4_E6BEG),
    .S1BEG(Tile_X2Y4_S1BEG),
    .S2BEG(Tile_X2Y4_S2BEG),
    .S2BEGb(Tile_X2Y4_S2BEGb),
    .S4BEG(Tile_X2Y4_S4BEG),
    .SS4BEG(Tile_X2Y4_SS4BEG),
    .W1BEG(Tile_X2Y4_W1BEG),
    .W2BEG(Tile_X2Y4_W2BEG),
    .W2BEGb(Tile_X2Y4_W2BEGb),
    .WW4BEG(Tile_X2Y4_WW4BEG),
    .W6BEG(Tile_X2Y4_W6BEG),
    .UserCLK(Tile_X2Y5_UserCLKo),
    .UserCLKo(Tile_X2Y4_UserCLKo),
    .FrameData(Tile_X1Y4_FrameData_O),
    .FrameData_O(Tile_X2Y4_FrameData_O),
    .FrameStrobe(Tile_X2Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y4_Emulate_Bitstream)
    )
`endif
    Tile_X3Y4_LUT4AB
    (
    .N1END(Tile_X3Y5_N1BEG),
    .N2MID(Tile_X3Y5_N2BEG),
    .N2END(Tile_X3Y5_N2BEGb),
    .N4END(Tile_X3Y5_N4BEG),
    .NN4END(Tile_X3Y5_NN4BEG),
    .Ci(Tile_X3Y5_Co),
    .E1END(Tile_X2Y4_E1BEG),
    .E2MID(Tile_X2Y4_E2BEG),
    .E2END(Tile_X2Y4_E2BEGb),
    .EE4END(Tile_X2Y4_EE4BEG),
    .E6END(Tile_X2Y4_E6BEG),
    .S1END(Tile_X3Y3_S1BEG),
    .S2MID(Tile_X3Y3_S2BEG),
    .S2END(Tile_X3Y3_S2BEGb),
    .S4END(Tile_X3Y3_S4BEG),
    .SS4END(Tile_X3Y3_SS4BEG),
    .W1END(Tile_X4Y4_W1BEG),
    .W2MID(Tile_X4Y4_W2BEG),
    .W2END(Tile_X4Y4_W2BEGb),
    .WW4END(Tile_X4Y4_WW4BEG),
    .W6END(Tile_X4Y4_W6BEG),
    .N1BEG(Tile_X3Y4_N1BEG),
    .N2BEG(Tile_X3Y4_N2BEG),
    .N2BEGb(Tile_X3Y4_N2BEGb),
    .N4BEG(Tile_X3Y4_N4BEG),
    .NN4BEG(Tile_X3Y4_NN4BEG),
    .Co(Tile_X3Y4_Co),
    .E1BEG(Tile_X3Y4_E1BEG),
    .E2BEG(Tile_X3Y4_E2BEG),
    .E2BEGb(Tile_X3Y4_E2BEGb),
    .EE4BEG(Tile_X3Y4_EE4BEG),
    .E6BEG(Tile_X3Y4_E6BEG),
    .S1BEG(Tile_X3Y4_S1BEG),
    .S2BEG(Tile_X3Y4_S2BEG),
    .S2BEGb(Tile_X3Y4_S2BEGb),
    .S4BEG(Tile_X3Y4_S4BEG),
    .SS4BEG(Tile_X3Y4_SS4BEG),
    .W1BEG(Tile_X3Y4_W1BEG),
    .W2BEG(Tile_X3Y4_W2BEG),
    .W2BEGb(Tile_X3Y4_W2BEGb),
    .WW4BEG(Tile_X3Y4_WW4BEG),
    .W6BEG(Tile_X3Y4_W6BEG),
    .UserCLK(Tile_X3Y5_UserCLKo),
    .UserCLKo(Tile_X3Y4_UserCLKo),
    .FrameData(Tile_X2Y4_FrameData_O),
    .FrameData_O(Tile_X3Y4_FrameData_O),
    .FrameStrobe(Tile_X3Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y4_Emulate_Bitstream)
    )
`endif
    Tile_X4Y4_LUT4AB
    (
    .N1END(Tile_X4Y5_N1BEG),
    .N2MID(Tile_X4Y5_N2BEG),
    .N2END(Tile_X4Y5_N2BEGb),
    .N4END(Tile_X4Y5_N4BEG),
    .NN4END(Tile_X4Y5_NN4BEG),
    .Ci(Tile_X4Y5_Co),
    .E1END(Tile_X3Y4_E1BEG),
    .E2MID(Tile_X3Y4_E2BEG),
    .E2END(Tile_X3Y4_E2BEGb),
    .EE4END(Tile_X3Y4_EE4BEG),
    .E6END(Tile_X3Y4_E6BEG),
    .S1END(Tile_X4Y3_S1BEG),
    .S2MID(Tile_X4Y3_S2BEG),
    .S2END(Tile_X4Y3_S2BEGb),
    .S4END(Tile_X4Y3_S4BEG),
    .SS4END(Tile_X4Y3_SS4BEG),
    .W1END(Tile_X5Y4_W1BEG),
    .W2MID(Tile_X5Y4_W2BEG),
    .W2END(Tile_X5Y4_W2BEGb),
    .WW4END(Tile_X5Y4_WW4BEG),
    .W6END(Tile_X5Y4_W6BEG),
    .N1BEG(Tile_X4Y4_N1BEG),
    .N2BEG(Tile_X4Y4_N2BEG),
    .N2BEGb(Tile_X4Y4_N2BEGb),
    .N4BEG(Tile_X4Y4_N4BEG),
    .NN4BEG(Tile_X4Y4_NN4BEG),
    .Co(Tile_X4Y4_Co),
    .E1BEG(Tile_X4Y4_E1BEG),
    .E2BEG(Tile_X4Y4_E2BEG),
    .E2BEGb(Tile_X4Y4_E2BEGb),
    .EE4BEG(Tile_X4Y4_EE4BEG),
    .E6BEG(Tile_X4Y4_E6BEG),
    .S1BEG(Tile_X4Y4_S1BEG),
    .S2BEG(Tile_X4Y4_S2BEG),
    .S2BEGb(Tile_X4Y4_S2BEGb),
    .S4BEG(Tile_X4Y4_S4BEG),
    .SS4BEG(Tile_X4Y4_SS4BEG),
    .W1BEG(Tile_X4Y4_W1BEG),
    .W2BEG(Tile_X4Y4_W2BEG),
    .W2BEGb(Tile_X4Y4_W2BEGb),
    .WW4BEG(Tile_X4Y4_WW4BEG),
    .W6BEG(Tile_X4Y4_W6BEG),
    .UserCLK(Tile_X4Y5_UserCLKo),
    .UserCLKo(Tile_X4Y4_UserCLKo),
    .FrameData(Tile_X3Y4_FrameData_O),
    .FrameData_O(Tile_X4Y4_FrameData_O),
    .FrameStrobe(Tile_X4Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y4_Emulate_Bitstream)
    )
`endif
    Tile_X5Y4_LUT4AB
    (
    .N1END(Tile_X5Y5_N1BEG),
    .N2MID(Tile_X5Y5_N2BEG),
    .N2END(Tile_X5Y5_N2BEGb),
    .N4END(Tile_X5Y5_N4BEG),
    .NN4END(Tile_X5Y5_NN4BEG),
    .Ci(Tile_X5Y5_Co),
    .E1END(Tile_X4Y4_E1BEG),
    .E2MID(Tile_X4Y4_E2BEG),
    .E2END(Tile_X4Y4_E2BEGb),
    .EE4END(Tile_X4Y4_EE4BEG),
    .E6END(Tile_X4Y4_E6BEG),
    .S1END(Tile_X5Y3_S1BEG),
    .S2MID(Tile_X5Y3_S2BEG),
    .S2END(Tile_X5Y3_S2BEGb),
    .S4END(Tile_X5Y3_S4BEG),
    .SS4END(Tile_X5Y3_SS4BEG),
    .W1END(Tile_X6Y4_W1BEG),
    .W2MID(Tile_X6Y4_W2BEG),
    .W2END(Tile_X6Y4_W2BEGb),
    .WW4END(Tile_X6Y4_WW4BEG),
    .W6END(Tile_X6Y4_W6BEG),
    .N1BEG(Tile_X5Y4_N1BEG),
    .N2BEG(Tile_X5Y4_N2BEG),
    .N2BEGb(Tile_X5Y4_N2BEGb),
    .N4BEG(Tile_X5Y4_N4BEG),
    .NN4BEG(Tile_X5Y4_NN4BEG),
    .Co(Tile_X5Y4_Co),
    .E1BEG(Tile_X5Y4_E1BEG),
    .E2BEG(Tile_X5Y4_E2BEG),
    .E2BEGb(Tile_X5Y4_E2BEGb),
    .EE4BEG(Tile_X5Y4_EE4BEG),
    .E6BEG(Tile_X5Y4_E6BEG),
    .S1BEG(Tile_X5Y4_S1BEG),
    .S2BEG(Tile_X5Y4_S2BEG),
    .S2BEGb(Tile_X5Y4_S2BEGb),
    .S4BEG(Tile_X5Y4_S4BEG),
    .SS4BEG(Tile_X5Y4_SS4BEG),
    .W1BEG(Tile_X5Y4_W1BEG),
    .W2BEG(Tile_X5Y4_W2BEG),
    .W2BEGb(Tile_X5Y4_W2BEGb),
    .WW4BEG(Tile_X5Y4_WW4BEG),
    .W6BEG(Tile_X5Y4_W6BEG),
    .UserCLK(Tile_X5Y5_UserCLKo),
    .UserCLKo(Tile_X5Y4_UserCLKo),
    .FrameData(Tile_X4Y4_FrameData_O),
    .FrameData_O(Tile_X5Y4_FrameData_O),
    .FrameStrobe(Tile_X5Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y4_Emulate_Bitstream)
    )
`endif
    Tile_X6Y4_LUT4AB
    (
    .N1END(Tile_X6Y5_N1BEG),
    .N2MID(Tile_X6Y5_N2BEG),
    .N2END(Tile_X6Y5_N2BEGb),
    .N4END(Tile_X6Y5_N4BEG),
    .NN4END(Tile_X6Y5_NN4BEG),
    .Ci(Tile_X6Y5_Co),
    .E1END(Tile_X5Y4_E1BEG),
    .E2MID(Tile_X5Y4_E2BEG),
    .E2END(Tile_X5Y4_E2BEGb),
    .EE4END(Tile_X5Y4_EE4BEG),
    .E6END(Tile_X5Y4_E6BEG),
    .S1END(Tile_X6Y3_S1BEG),
    .S2MID(Tile_X6Y3_S2BEG),
    .S2END(Tile_X6Y3_S2BEGb),
    .S4END(Tile_X6Y3_S4BEG),
    .SS4END(Tile_X6Y3_SS4BEG),
    .W1END(Tile_X7Y4_W1BEG),
    .W2MID(Tile_X7Y4_W2BEG),
    .W2END(Tile_X7Y4_W2BEGb),
    .WW4END(Tile_X7Y4_WW4BEG),
    .W6END(Tile_X7Y4_W6BEG),
    .N1BEG(Tile_X6Y4_N1BEG),
    .N2BEG(Tile_X6Y4_N2BEG),
    .N2BEGb(Tile_X6Y4_N2BEGb),
    .N4BEG(Tile_X6Y4_N4BEG),
    .NN4BEG(Tile_X6Y4_NN4BEG),
    .Co(Tile_X6Y4_Co),
    .E1BEG(Tile_X6Y4_E1BEG),
    .E2BEG(Tile_X6Y4_E2BEG),
    .E2BEGb(Tile_X6Y4_E2BEGb),
    .EE4BEG(Tile_X6Y4_EE4BEG),
    .E6BEG(Tile_X6Y4_E6BEG),
    .S1BEG(Tile_X6Y4_S1BEG),
    .S2BEG(Tile_X6Y4_S2BEG),
    .S2BEGb(Tile_X6Y4_S2BEGb),
    .S4BEG(Tile_X6Y4_S4BEG),
    .SS4BEG(Tile_X6Y4_SS4BEG),
    .W1BEG(Tile_X6Y4_W1BEG),
    .W2BEG(Tile_X6Y4_W2BEG),
    .W2BEGb(Tile_X6Y4_W2BEGb),
    .WW4BEG(Tile_X6Y4_WW4BEG),
    .W6BEG(Tile_X6Y4_W6BEG),
    .UserCLK(Tile_X6Y5_UserCLKo),
    .UserCLKo(Tile_X6Y4_UserCLKo),
    .FrameData(Tile_X5Y4_FrameData_O),
    .FrameData_O(Tile_X6Y4_FrameData_O),
    .FrameStrobe(Tile_X6Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y4_Emulate_Bitstream)
    )
`endif
    Tile_X7Y4_LUT4AB
    (
    .N1END(Tile_X7Y5_N1BEG),
    .N2MID(Tile_X7Y5_N2BEG),
    .N2END(Tile_X7Y5_N2BEGb),
    .N4END(Tile_X7Y5_N4BEG),
    .NN4END(Tile_X7Y5_NN4BEG),
    .Ci(Tile_X7Y5_Co),
    .E1END(Tile_X6Y4_E1BEG),
    .E2MID(Tile_X6Y4_E2BEG),
    .E2END(Tile_X6Y4_E2BEGb),
    .EE4END(Tile_X6Y4_EE4BEG),
    .E6END(Tile_X6Y4_E6BEG),
    .S1END(Tile_X7Y3_S1BEG),
    .S2MID(Tile_X7Y3_S2BEG),
    .S2END(Tile_X7Y3_S2BEGb),
    .S4END(Tile_X7Y3_S4BEG),
    .SS4END(Tile_X7Y3_SS4BEG),
    .W1END(Tile_X8Y4_W1BEG),
    .W2MID(Tile_X8Y4_W2BEG),
    .W2END(Tile_X8Y4_W2BEGb),
    .WW4END(Tile_X8Y4_WW4BEG),
    .W6END(Tile_X8Y4_W6BEG),
    .N1BEG(Tile_X7Y4_N1BEG),
    .N2BEG(Tile_X7Y4_N2BEG),
    .N2BEGb(Tile_X7Y4_N2BEGb),
    .N4BEG(Tile_X7Y4_N4BEG),
    .NN4BEG(Tile_X7Y4_NN4BEG),
    .Co(Tile_X7Y4_Co),
    .E1BEG(Tile_X7Y4_E1BEG),
    .E2BEG(Tile_X7Y4_E2BEG),
    .E2BEGb(Tile_X7Y4_E2BEGb),
    .EE4BEG(Tile_X7Y4_EE4BEG),
    .E6BEG(Tile_X7Y4_E6BEG),
    .S1BEG(Tile_X7Y4_S1BEG),
    .S2BEG(Tile_X7Y4_S2BEG),
    .S2BEGb(Tile_X7Y4_S2BEGb),
    .S4BEG(Tile_X7Y4_S4BEG),
    .SS4BEG(Tile_X7Y4_SS4BEG),
    .W1BEG(Tile_X7Y4_W1BEG),
    .W2BEG(Tile_X7Y4_W2BEG),
    .W2BEGb(Tile_X7Y4_W2BEGb),
    .WW4BEG(Tile_X7Y4_WW4BEG),
    .W6BEG(Tile_X7Y4_W6BEG),
    .UserCLK(Tile_X7Y5_UserCLKo),
    .UserCLKo(Tile_X7Y4_UserCLKo),
    .FrameData(Tile_X6Y4_FrameData_O),
    .FrameData_O(Tile_X7Y4_FrameData_O),
    .FrameStrobe(Tile_X7Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RAM_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y4_Emulate_Bitstream)
    )
`endif
    Tile_X8Y4_RAM_IO
    (
    .N1END(Tile_X8Y5_N1BEG),
    .N2MID(Tile_X8Y5_N2BEG),
    .N2END(Tile_X8Y5_N2BEGb),
    .N4END(Tile_X8Y5_N4BEG),
    .E1END(Tile_X7Y4_E1BEG),
    .E2MID(Tile_X7Y4_E2BEG),
    .E2END(Tile_X7Y4_E2BEGb),
    .EE4END(Tile_X7Y4_EE4BEG),
    .E6END(Tile_X7Y4_E6BEG),
    .S1END(Tile_X8Y3_S1BEG),
    .S2MID(Tile_X8Y3_S2BEG),
    .S2END(Tile_X8Y3_S2BEGb),
    .S4END(Tile_X8Y3_S4BEG),
    .N1BEG(Tile_X8Y4_N1BEG),
    .N2BEG(Tile_X8Y4_N2BEG),
    .N2BEGb(Tile_X8Y4_N2BEGb),
    .N4BEG(Tile_X8Y4_N4BEG),
    .S1BEG(Tile_X8Y4_S1BEG),
    .S2BEG(Tile_X8Y4_S2BEG),
    .S2BEGb(Tile_X8Y4_S2BEGb),
    .S4BEG(Tile_X8Y4_S4BEG),
    .W1BEG(Tile_X8Y4_W1BEG),
    .W2BEG(Tile_X8Y4_W2BEG),
    .W2BEGb(Tile_X8Y4_W2BEGb),
    .WW4BEG(Tile_X8Y4_WW4BEG),
    .W6BEG(Tile_X8Y4_W6BEG),
    .RAM2FAB_D0_I0(Tile_X8Y4_RAM2FAB_D0_I0),
    .RAM2FAB_D0_I1(Tile_X8Y4_RAM2FAB_D0_I1),
    .RAM2FAB_D0_I2(Tile_X8Y4_RAM2FAB_D0_I2),
    .RAM2FAB_D0_I3(Tile_X8Y4_RAM2FAB_D0_I3),
    .RAM2FAB_D1_I0(Tile_X8Y4_RAM2FAB_D1_I0),
    .RAM2FAB_D1_I1(Tile_X8Y4_RAM2FAB_D1_I1),
    .RAM2FAB_D1_I2(Tile_X8Y4_RAM2FAB_D1_I2),
    .RAM2FAB_D1_I3(Tile_X8Y4_RAM2FAB_D1_I3),
    .RAM2FAB_D2_I0(Tile_X8Y4_RAM2FAB_D2_I0),
    .RAM2FAB_D2_I1(Tile_X8Y4_RAM2FAB_D2_I1),
    .RAM2FAB_D2_I2(Tile_X8Y4_RAM2FAB_D2_I2),
    .RAM2FAB_D2_I3(Tile_X8Y4_RAM2FAB_D2_I3),
    .RAM2FAB_D3_I0(Tile_X8Y4_RAM2FAB_D3_I0),
    .RAM2FAB_D3_I1(Tile_X8Y4_RAM2FAB_D3_I1),
    .RAM2FAB_D3_I2(Tile_X8Y4_RAM2FAB_D3_I2),
    .RAM2FAB_D3_I3(Tile_X8Y4_RAM2FAB_D3_I3),
    .FAB2RAM_D0_O0(Tile_X8Y4_FAB2RAM_D0_O0),
    .FAB2RAM_D0_O1(Tile_X8Y4_FAB2RAM_D0_O1),
    .FAB2RAM_D0_O2(Tile_X8Y4_FAB2RAM_D0_O2),
    .FAB2RAM_D0_O3(Tile_X8Y4_FAB2RAM_D0_O3),
    .FAB2RAM_D1_O0(Tile_X8Y4_FAB2RAM_D1_O0),
    .FAB2RAM_D1_O1(Tile_X8Y4_FAB2RAM_D1_O1),
    .FAB2RAM_D1_O2(Tile_X8Y4_FAB2RAM_D1_O2),
    .FAB2RAM_D1_O3(Tile_X8Y4_FAB2RAM_D1_O3),
    .FAB2RAM_D2_O0(Tile_X8Y4_FAB2RAM_D2_O0),
    .FAB2RAM_D2_O1(Tile_X8Y4_FAB2RAM_D2_O1),
    .FAB2RAM_D2_O2(Tile_X8Y4_FAB2RAM_D2_O2),
    .FAB2RAM_D2_O3(Tile_X8Y4_FAB2RAM_D2_O3),
    .FAB2RAM_D3_O0(Tile_X8Y4_FAB2RAM_D3_O0),
    .FAB2RAM_D3_O1(Tile_X8Y4_FAB2RAM_D3_O1),
    .FAB2RAM_D3_O2(Tile_X8Y4_FAB2RAM_D3_O2),
    .FAB2RAM_D3_O3(Tile_X8Y4_FAB2RAM_D3_O3),
    .FAB2RAM_A0_O0(Tile_X8Y4_FAB2RAM_A0_O0),
    .FAB2RAM_A0_O1(Tile_X8Y4_FAB2RAM_A0_O1),
    .FAB2RAM_A0_O2(Tile_X8Y4_FAB2RAM_A0_O2),
    .FAB2RAM_A0_O3(Tile_X8Y4_FAB2RAM_A0_O3),
    .FAB2RAM_A1_O0(Tile_X8Y4_FAB2RAM_A1_O0),
    .FAB2RAM_A1_O1(Tile_X8Y4_FAB2RAM_A1_O1),
    .FAB2RAM_A1_O2(Tile_X8Y4_FAB2RAM_A1_O2),
    .FAB2RAM_A1_O3(Tile_X8Y4_FAB2RAM_A1_O3),
    .FAB2RAM_C_O0(Tile_X8Y4_FAB2RAM_C_O0),
    .FAB2RAM_C_O1(Tile_X8Y4_FAB2RAM_C_O1),
    .FAB2RAM_C_O2(Tile_X8Y4_FAB2RAM_C_O2),
    .FAB2RAM_C_O3(Tile_X8Y4_FAB2RAM_C_O3),
    .Config_accessC_bit0(Tile_X8Y4_Config_accessC_bit0),
    .Config_accessC_bit1(Tile_X8Y4_Config_accessC_bit1),
    .Config_accessC_bit2(Tile_X8Y4_Config_accessC_bit2),
    .Config_accessC_bit3(Tile_X8Y4_Config_accessC_bit3),
    .UserCLK(Tile_X8Y5_UserCLKo),
    .UserCLKo(Tile_X8Y4_UserCLKo),
    .FrameData(Tile_X7Y4_FrameData_O),
    .FrameData_O(Tile_X8Y4_FrameData_O),
    .FrameStrobe(Tile_X8Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y5_Emulate_Bitstream)
    )
`endif
    Tile_X0Y5_W_IO
    (
    .W1END(Tile_X1Y5_W1BEG),
    .W2MID(Tile_X1Y5_W2BEG),
    .W2END(Tile_X1Y5_W2BEGb),
    .WW4END(Tile_X1Y5_WW4BEG),
    .W6END(Tile_X1Y5_W6BEG),
    .E1BEG(Tile_X0Y5_E1BEG),
    .E2BEG(Tile_X0Y5_E2BEG),
    .E2BEGb(Tile_X0Y5_E2BEGb),
    .EE4BEG(Tile_X0Y5_EE4BEG),
    .E6BEG(Tile_X0Y5_E6BEG),
    .A_O_top(Tile_X0Y5_A_O_top),
    .A_I_top(Tile_X0Y5_A_I_top),
    .A_T_top(Tile_X0Y5_A_T_top),
    .B_O_top(Tile_X0Y5_B_O_top),
    .B_I_top(Tile_X0Y5_B_I_top),
    .B_T_top(Tile_X0Y5_B_T_top),
    .A_config_C_bit0(Tile_X0Y5_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y5_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y5_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y5_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y5_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y5_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y5_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y5_B_config_C_bit3),
    .UserCLK(Tile_X0Y6_UserCLKo),
    .UserCLKo(Tile_X0Y5_UserCLKo),
    .FrameData(Tile_Y5_FrameData),
    .FrameData_O(Tile_X0Y5_FrameData_O),
    .FrameStrobe(Tile_X0Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y5_Emulate_Bitstream)
    )
`endif
    Tile_X1Y5_LUT4AB
    (
    .N1END(Tile_X1Y6_N1BEG),
    .N2MID(Tile_X1Y6_N2BEG),
    .N2END(Tile_X1Y6_N2BEGb),
    .N4END(Tile_X1Y6_N4BEG),
    .NN4END(Tile_X1Y6_NN4BEG),
    .Ci(Tile_X1Y6_Co),
    .E1END(Tile_X0Y5_E1BEG),
    .E2MID(Tile_X0Y5_E2BEG),
    .E2END(Tile_X0Y5_E2BEGb),
    .EE4END(Tile_X0Y5_EE4BEG),
    .E6END(Tile_X0Y5_E6BEG),
    .S1END(Tile_X1Y4_S1BEG),
    .S2MID(Tile_X1Y4_S2BEG),
    .S2END(Tile_X1Y4_S2BEGb),
    .S4END(Tile_X1Y4_S4BEG),
    .SS4END(Tile_X1Y4_SS4BEG),
    .W1END(Tile_X2Y5_W1BEG),
    .W2MID(Tile_X2Y5_W2BEG),
    .W2END(Tile_X2Y5_W2BEGb),
    .WW4END(Tile_X2Y5_WW4BEG),
    .W6END(Tile_X2Y5_W6BEG),
    .N1BEG(Tile_X1Y5_N1BEG),
    .N2BEG(Tile_X1Y5_N2BEG),
    .N2BEGb(Tile_X1Y5_N2BEGb),
    .N4BEG(Tile_X1Y5_N4BEG),
    .NN4BEG(Tile_X1Y5_NN4BEG),
    .Co(Tile_X1Y5_Co),
    .E1BEG(Tile_X1Y5_E1BEG),
    .E2BEG(Tile_X1Y5_E2BEG),
    .E2BEGb(Tile_X1Y5_E2BEGb),
    .EE4BEG(Tile_X1Y5_EE4BEG),
    .E6BEG(Tile_X1Y5_E6BEG),
    .S1BEG(Tile_X1Y5_S1BEG),
    .S2BEG(Tile_X1Y5_S2BEG),
    .S2BEGb(Tile_X1Y5_S2BEGb),
    .S4BEG(Tile_X1Y5_S4BEG),
    .SS4BEG(Tile_X1Y5_SS4BEG),
    .W1BEG(Tile_X1Y5_W1BEG),
    .W2BEG(Tile_X1Y5_W2BEG),
    .W2BEGb(Tile_X1Y5_W2BEGb),
    .WW4BEG(Tile_X1Y5_WW4BEG),
    .W6BEG(Tile_X1Y5_W6BEG),
    .UserCLK(Tile_X1Y6_UserCLKo),
    .UserCLKo(Tile_X1Y5_UserCLKo),
    .FrameData(Tile_X0Y5_FrameData_O),
    .FrameData_O(Tile_X1Y5_FrameData_O),
    .FrameStrobe(Tile_X1Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y5_Emulate_Bitstream)
    )
`endif
    Tile_X2Y5_LUT4AB
    (
    .N1END(Tile_X2Y6_N1BEG),
    .N2MID(Tile_X2Y6_N2BEG),
    .N2END(Tile_X2Y6_N2BEGb),
    .N4END(Tile_X2Y6_N4BEG),
    .NN4END(Tile_X2Y6_NN4BEG),
    .Ci(Tile_X2Y6_Co),
    .E1END(Tile_X1Y5_E1BEG),
    .E2MID(Tile_X1Y5_E2BEG),
    .E2END(Tile_X1Y5_E2BEGb),
    .EE4END(Tile_X1Y5_EE4BEG),
    .E6END(Tile_X1Y5_E6BEG),
    .S1END(Tile_X2Y4_S1BEG),
    .S2MID(Tile_X2Y4_S2BEG),
    .S2END(Tile_X2Y4_S2BEGb),
    .S4END(Tile_X2Y4_S4BEG),
    .SS4END(Tile_X2Y4_SS4BEG),
    .W1END(Tile_X3Y5_W1BEG),
    .W2MID(Tile_X3Y5_W2BEG),
    .W2END(Tile_X3Y5_W2BEGb),
    .WW4END(Tile_X3Y5_WW4BEG),
    .W6END(Tile_X3Y5_W6BEG),
    .N1BEG(Tile_X2Y5_N1BEG),
    .N2BEG(Tile_X2Y5_N2BEG),
    .N2BEGb(Tile_X2Y5_N2BEGb),
    .N4BEG(Tile_X2Y5_N4BEG),
    .NN4BEG(Tile_X2Y5_NN4BEG),
    .Co(Tile_X2Y5_Co),
    .E1BEG(Tile_X2Y5_E1BEG),
    .E2BEG(Tile_X2Y5_E2BEG),
    .E2BEGb(Tile_X2Y5_E2BEGb),
    .EE4BEG(Tile_X2Y5_EE4BEG),
    .E6BEG(Tile_X2Y5_E6BEG),
    .S1BEG(Tile_X2Y5_S1BEG),
    .S2BEG(Tile_X2Y5_S2BEG),
    .S2BEGb(Tile_X2Y5_S2BEGb),
    .S4BEG(Tile_X2Y5_S4BEG),
    .SS4BEG(Tile_X2Y5_SS4BEG),
    .W1BEG(Tile_X2Y5_W1BEG),
    .W2BEG(Tile_X2Y5_W2BEG),
    .W2BEGb(Tile_X2Y5_W2BEGb),
    .WW4BEG(Tile_X2Y5_WW4BEG),
    .W6BEG(Tile_X2Y5_W6BEG),
    .UserCLK(Tile_X2Y6_UserCLKo),
    .UserCLKo(Tile_X2Y5_UserCLKo),
    .FrameData(Tile_X1Y5_FrameData_O),
    .FrameData_O(Tile_X2Y5_FrameData_O),
    .FrameStrobe(Tile_X2Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y5_Emulate_Bitstream)
    )
`endif
    Tile_X3Y5_LUT4AB
    (
    .N1END(Tile_X3Y6_N1BEG),
    .N2MID(Tile_X3Y6_N2BEG),
    .N2END(Tile_X3Y6_N2BEGb),
    .N4END(Tile_X3Y6_N4BEG),
    .NN4END(Tile_X3Y6_NN4BEG),
    .Ci(Tile_X3Y6_Co),
    .E1END(Tile_X2Y5_E1BEG),
    .E2MID(Tile_X2Y5_E2BEG),
    .E2END(Tile_X2Y5_E2BEGb),
    .EE4END(Tile_X2Y5_EE4BEG),
    .E6END(Tile_X2Y5_E6BEG),
    .S1END(Tile_X3Y4_S1BEG),
    .S2MID(Tile_X3Y4_S2BEG),
    .S2END(Tile_X3Y4_S2BEGb),
    .S4END(Tile_X3Y4_S4BEG),
    .SS4END(Tile_X3Y4_SS4BEG),
    .W1END(Tile_X4Y5_W1BEG),
    .W2MID(Tile_X4Y5_W2BEG),
    .W2END(Tile_X4Y5_W2BEGb),
    .WW4END(Tile_X4Y5_WW4BEG),
    .W6END(Tile_X4Y5_W6BEG),
    .N1BEG(Tile_X3Y5_N1BEG),
    .N2BEG(Tile_X3Y5_N2BEG),
    .N2BEGb(Tile_X3Y5_N2BEGb),
    .N4BEG(Tile_X3Y5_N4BEG),
    .NN4BEG(Tile_X3Y5_NN4BEG),
    .Co(Tile_X3Y5_Co),
    .E1BEG(Tile_X3Y5_E1BEG),
    .E2BEG(Tile_X3Y5_E2BEG),
    .E2BEGb(Tile_X3Y5_E2BEGb),
    .EE4BEG(Tile_X3Y5_EE4BEG),
    .E6BEG(Tile_X3Y5_E6BEG),
    .S1BEG(Tile_X3Y5_S1BEG),
    .S2BEG(Tile_X3Y5_S2BEG),
    .S2BEGb(Tile_X3Y5_S2BEGb),
    .S4BEG(Tile_X3Y5_S4BEG),
    .SS4BEG(Tile_X3Y5_SS4BEG),
    .W1BEG(Tile_X3Y5_W1BEG),
    .W2BEG(Tile_X3Y5_W2BEG),
    .W2BEGb(Tile_X3Y5_W2BEGb),
    .WW4BEG(Tile_X3Y5_WW4BEG),
    .W6BEG(Tile_X3Y5_W6BEG),
    .UserCLK(Tile_X3Y6_UserCLKo),
    .UserCLKo(Tile_X3Y5_UserCLKo),
    .FrameData(Tile_X2Y5_FrameData_O),
    .FrameData_O(Tile_X3Y5_FrameData_O),
    .FrameStrobe(Tile_X3Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y5_Emulate_Bitstream)
    )
`endif
    Tile_X4Y5_LUT4AB
    (
    .N1END(Tile_X4Y6_N1BEG),
    .N2MID(Tile_X4Y6_N2BEG),
    .N2END(Tile_X4Y6_N2BEGb),
    .N4END(Tile_X4Y6_N4BEG),
    .NN4END(Tile_X4Y6_NN4BEG),
    .Ci(Tile_X4Y6_Co),
    .E1END(Tile_X3Y5_E1BEG),
    .E2MID(Tile_X3Y5_E2BEG),
    .E2END(Tile_X3Y5_E2BEGb),
    .EE4END(Tile_X3Y5_EE4BEG),
    .E6END(Tile_X3Y5_E6BEG),
    .S1END(Tile_X4Y4_S1BEG),
    .S2MID(Tile_X4Y4_S2BEG),
    .S2END(Tile_X4Y4_S2BEGb),
    .S4END(Tile_X4Y4_S4BEG),
    .SS4END(Tile_X4Y4_SS4BEG),
    .W1END(Tile_X5Y5_W1BEG),
    .W2MID(Tile_X5Y5_W2BEG),
    .W2END(Tile_X5Y5_W2BEGb),
    .WW4END(Tile_X5Y5_WW4BEG),
    .W6END(Tile_X5Y5_W6BEG),
    .N1BEG(Tile_X4Y5_N1BEG),
    .N2BEG(Tile_X4Y5_N2BEG),
    .N2BEGb(Tile_X4Y5_N2BEGb),
    .N4BEG(Tile_X4Y5_N4BEG),
    .NN4BEG(Tile_X4Y5_NN4BEG),
    .Co(Tile_X4Y5_Co),
    .E1BEG(Tile_X4Y5_E1BEG),
    .E2BEG(Tile_X4Y5_E2BEG),
    .E2BEGb(Tile_X4Y5_E2BEGb),
    .EE4BEG(Tile_X4Y5_EE4BEG),
    .E6BEG(Tile_X4Y5_E6BEG),
    .S1BEG(Tile_X4Y5_S1BEG),
    .S2BEG(Tile_X4Y5_S2BEG),
    .S2BEGb(Tile_X4Y5_S2BEGb),
    .S4BEG(Tile_X4Y5_S4BEG),
    .SS4BEG(Tile_X4Y5_SS4BEG),
    .W1BEG(Tile_X4Y5_W1BEG),
    .W2BEG(Tile_X4Y5_W2BEG),
    .W2BEGb(Tile_X4Y5_W2BEGb),
    .WW4BEG(Tile_X4Y5_WW4BEG),
    .W6BEG(Tile_X4Y5_W6BEG),
    .UserCLK(Tile_X4Y6_UserCLKo),
    .UserCLKo(Tile_X4Y5_UserCLKo),
    .FrameData(Tile_X3Y5_FrameData_O),
    .FrameData_O(Tile_X4Y5_FrameData_O),
    .FrameStrobe(Tile_X4Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y5_Emulate_Bitstream)
    )
`endif
    Tile_X5Y5_LUT4AB
    (
    .N1END(Tile_X5Y6_N1BEG),
    .N2MID(Tile_X5Y6_N2BEG),
    .N2END(Tile_X5Y6_N2BEGb),
    .N4END(Tile_X5Y6_N4BEG),
    .NN4END(Tile_X5Y6_NN4BEG),
    .Ci(Tile_X5Y6_Co),
    .E1END(Tile_X4Y5_E1BEG),
    .E2MID(Tile_X4Y5_E2BEG),
    .E2END(Tile_X4Y5_E2BEGb),
    .EE4END(Tile_X4Y5_EE4BEG),
    .E6END(Tile_X4Y5_E6BEG),
    .S1END(Tile_X5Y4_S1BEG),
    .S2MID(Tile_X5Y4_S2BEG),
    .S2END(Tile_X5Y4_S2BEGb),
    .S4END(Tile_X5Y4_S4BEG),
    .SS4END(Tile_X5Y4_SS4BEG),
    .W1END(Tile_X6Y5_W1BEG),
    .W2MID(Tile_X6Y5_W2BEG),
    .W2END(Tile_X6Y5_W2BEGb),
    .WW4END(Tile_X6Y5_WW4BEG),
    .W6END(Tile_X6Y5_W6BEG),
    .N1BEG(Tile_X5Y5_N1BEG),
    .N2BEG(Tile_X5Y5_N2BEG),
    .N2BEGb(Tile_X5Y5_N2BEGb),
    .N4BEG(Tile_X5Y5_N4BEG),
    .NN4BEG(Tile_X5Y5_NN4BEG),
    .Co(Tile_X5Y5_Co),
    .E1BEG(Tile_X5Y5_E1BEG),
    .E2BEG(Tile_X5Y5_E2BEG),
    .E2BEGb(Tile_X5Y5_E2BEGb),
    .EE4BEG(Tile_X5Y5_EE4BEG),
    .E6BEG(Tile_X5Y5_E6BEG),
    .S1BEG(Tile_X5Y5_S1BEG),
    .S2BEG(Tile_X5Y5_S2BEG),
    .S2BEGb(Tile_X5Y5_S2BEGb),
    .S4BEG(Tile_X5Y5_S4BEG),
    .SS4BEG(Tile_X5Y5_SS4BEG),
    .W1BEG(Tile_X5Y5_W1BEG),
    .W2BEG(Tile_X5Y5_W2BEG),
    .W2BEGb(Tile_X5Y5_W2BEGb),
    .WW4BEG(Tile_X5Y5_WW4BEG),
    .W6BEG(Tile_X5Y5_W6BEG),
    .UserCLK(Tile_X5Y6_UserCLKo),
    .UserCLKo(Tile_X5Y5_UserCLKo),
    .FrameData(Tile_X4Y5_FrameData_O),
    .FrameData_O(Tile_X5Y5_FrameData_O),
    .FrameStrobe(Tile_X5Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y5_Emulate_Bitstream)
    )
`endif
    Tile_X6Y5_LUT4AB
    (
    .N1END(Tile_X6Y6_N1BEG),
    .N2MID(Tile_X6Y6_N2BEG),
    .N2END(Tile_X6Y6_N2BEGb),
    .N4END(Tile_X6Y6_N4BEG),
    .NN4END(Tile_X6Y6_NN4BEG),
    .Ci(Tile_X6Y6_Co),
    .E1END(Tile_X5Y5_E1BEG),
    .E2MID(Tile_X5Y5_E2BEG),
    .E2END(Tile_X5Y5_E2BEGb),
    .EE4END(Tile_X5Y5_EE4BEG),
    .E6END(Tile_X5Y5_E6BEG),
    .S1END(Tile_X6Y4_S1BEG),
    .S2MID(Tile_X6Y4_S2BEG),
    .S2END(Tile_X6Y4_S2BEGb),
    .S4END(Tile_X6Y4_S4BEG),
    .SS4END(Tile_X6Y4_SS4BEG),
    .W1END(Tile_X7Y5_W1BEG),
    .W2MID(Tile_X7Y5_W2BEG),
    .W2END(Tile_X7Y5_W2BEGb),
    .WW4END(Tile_X7Y5_WW4BEG),
    .W6END(Tile_X7Y5_W6BEG),
    .N1BEG(Tile_X6Y5_N1BEG),
    .N2BEG(Tile_X6Y5_N2BEG),
    .N2BEGb(Tile_X6Y5_N2BEGb),
    .N4BEG(Tile_X6Y5_N4BEG),
    .NN4BEG(Tile_X6Y5_NN4BEG),
    .Co(Tile_X6Y5_Co),
    .E1BEG(Tile_X6Y5_E1BEG),
    .E2BEG(Tile_X6Y5_E2BEG),
    .E2BEGb(Tile_X6Y5_E2BEGb),
    .EE4BEG(Tile_X6Y5_EE4BEG),
    .E6BEG(Tile_X6Y5_E6BEG),
    .S1BEG(Tile_X6Y5_S1BEG),
    .S2BEG(Tile_X6Y5_S2BEG),
    .S2BEGb(Tile_X6Y5_S2BEGb),
    .S4BEG(Tile_X6Y5_S4BEG),
    .SS4BEG(Tile_X6Y5_SS4BEG),
    .W1BEG(Tile_X6Y5_W1BEG),
    .W2BEG(Tile_X6Y5_W2BEG),
    .W2BEGb(Tile_X6Y5_W2BEGb),
    .WW4BEG(Tile_X6Y5_WW4BEG),
    .W6BEG(Tile_X6Y5_W6BEG),
    .UserCLK(Tile_X6Y6_UserCLKo),
    .UserCLKo(Tile_X6Y5_UserCLKo),
    .FrameData(Tile_X5Y5_FrameData_O),
    .FrameData_O(Tile_X6Y5_FrameData_O),
    .FrameStrobe(Tile_X6Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y5_Emulate_Bitstream)
    )
`endif
    Tile_X7Y5_LUT4AB
    (
    .N1END(Tile_X7Y6_N1BEG),
    .N2MID(Tile_X7Y6_N2BEG),
    .N2END(Tile_X7Y6_N2BEGb),
    .N4END(Tile_X7Y6_N4BEG),
    .NN4END(Tile_X7Y6_NN4BEG),
    .Ci(Tile_X7Y6_Co),
    .E1END(Tile_X6Y5_E1BEG),
    .E2MID(Tile_X6Y5_E2BEG),
    .E2END(Tile_X6Y5_E2BEGb),
    .EE4END(Tile_X6Y5_EE4BEG),
    .E6END(Tile_X6Y5_E6BEG),
    .S1END(Tile_X7Y4_S1BEG),
    .S2MID(Tile_X7Y4_S2BEG),
    .S2END(Tile_X7Y4_S2BEGb),
    .S4END(Tile_X7Y4_S4BEG),
    .SS4END(Tile_X7Y4_SS4BEG),
    .W1END(Tile_X8Y5_W1BEG),
    .W2MID(Tile_X8Y5_W2BEG),
    .W2END(Tile_X8Y5_W2BEGb),
    .WW4END(Tile_X8Y5_WW4BEG),
    .W6END(Tile_X8Y5_W6BEG),
    .N1BEG(Tile_X7Y5_N1BEG),
    .N2BEG(Tile_X7Y5_N2BEG),
    .N2BEGb(Tile_X7Y5_N2BEGb),
    .N4BEG(Tile_X7Y5_N4BEG),
    .NN4BEG(Tile_X7Y5_NN4BEG),
    .Co(Tile_X7Y5_Co),
    .E1BEG(Tile_X7Y5_E1BEG),
    .E2BEG(Tile_X7Y5_E2BEG),
    .E2BEGb(Tile_X7Y5_E2BEGb),
    .EE4BEG(Tile_X7Y5_EE4BEG),
    .E6BEG(Tile_X7Y5_E6BEG),
    .S1BEG(Tile_X7Y5_S1BEG),
    .S2BEG(Tile_X7Y5_S2BEG),
    .S2BEGb(Tile_X7Y5_S2BEGb),
    .S4BEG(Tile_X7Y5_S4BEG),
    .SS4BEG(Tile_X7Y5_SS4BEG),
    .W1BEG(Tile_X7Y5_W1BEG),
    .W2BEG(Tile_X7Y5_W2BEG),
    .W2BEGb(Tile_X7Y5_W2BEGb),
    .WW4BEG(Tile_X7Y5_WW4BEG),
    .W6BEG(Tile_X7Y5_W6BEG),
    .UserCLK(Tile_X7Y6_UserCLKo),
    .UserCLKo(Tile_X7Y5_UserCLKo),
    .FrameData(Tile_X6Y5_FrameData_O),
    .FrameData_O(Tile_X7Y5_FrameData_O),
    .FrameStrobe(Tile_X7Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RAM_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y5_Emulate_Bitstream)
    )
`endif
    Tile_X8Y5_RAM_IO
    (
    .N1END(Tile_X8Y6_N1BEG),
    .N2MID(Tile_X8Y6_N2BEG),
    .N2END(Tile_X8Y6_N2BEGb),
    .N4END(Tile_X8Y6_N4BEG),
    .E1END(Tile_X7Y5_E1BEG),
    .E2MID(Tile_X7Y5_E2BEG),
    .E2END(Tile_X7Y5_E2BEGb),
    .EE4END(Tile_X7Y5_EE4BEG),
    .E6END(Tile_X7Y5_E6BEG),
    .S1END(Tile_X8Y4_S1BEG),
    .S2MID(Tile_X8Y4_S2BEG),
    .S2END(Tile_X8Y4_S2BEGb),
    .S4END(Tile_X8Y4_S4BEG),
    .N1BEG(Tile_X8Y5_N1BEG),
    .N2BEG(Tile_X8Y5_N2BEG),
    .N2BEGb(Tile_X8Y5_N2BEGb),
    .N4BEG(Tile_X8Y5_N4BEG),
    .S1BEG(Tile_X8Y5_S1BEG),
    .S2BEG(Tile_X8Y5_S2BEG),
    .S2BEGb(Tile_X8Y5_S2BEGb),
    .S4BEG(Tile_X8Y5_S4BEG),
    .W1BEG(Tile_X8Y5_W1BEG),
    .W2BEG(Tile_X8Y5_W2BEG),
    .W2BEGb(Tile_X8Y5_W2BEGb),
    .WW4BEG(Tile_X8Y5_WW4BEG),
    .W6BEG(Tile_X8Y5_W6BEG),
    .RAM2FAB_D0_I0(Tile_X8Y5_RAM2FAB_D0_I0),
    .RAM2FAB_D0_I1(Tile_X8Y5_RAM2FAB_D0_I1),
    .RAM2FAB_D0_I2(Tile_X8Y5_RAM2FAB_D0_I2),
    .RAM2FAB_D0_I3(Tile_X8Y5_RAM2FAB_D0_I3),
    .RAM2FAB_D1_I0(Tile_X8Y5_RAM2FAB_D1_I0),
    .RAM2FAB_D1_I1(Tile_X8Y5_RAM2FAB_D1_I1),
    .RAM2FAB_D1_I2(Tile_X8Y5_RAM2FAB_D1_I2),
    .RAM2FAB_D1_I3(Tile_X8Y5_RAM2FAB_D1_I3),
    .RAM2FAB_D2_I0(Tile_X8Y5_RAM2FAB_D2_I0),
    .RAM2FAB_D2_I1(Tile_X8Y5_RAM2FAB_D2_I1),
    .RAM2FAB_D2_I2(Tile_X8Y5_RAM2FAB_D2_I2),
    .RAM2FAB_D2_I3(Tile_X8Y5_RAM2FAB_D2_I3),
    .RAM2FAB_D3_I0(Tile_X8Y5_RAM2FAB_D3_I0),
    .RAM2FAB_D3_I1(Tile_X8Y5_RAM2FAB_D3_I1),
    .RAM2FAB_D3_I2(Tile_X8Y5_RAM2FAB_D3_I2),
    .RAM2FAB_D3_I3(Tile_X8Y5_RAM2FAB_D3_I3),
    .FAB2RAM_D0_O0(Tile_X8Y5_FAB2RAM_D0_O0),
    .FAB2RAM_D0_O1(Tile_X8Y5_FAB2RAM_D0_O1),
    .FAB2RAM_D0_O2(Tile_X8Y5_FAB2RAM_D0_O2),
    .FAB2RAM_D0_O3(Tile_X8Y5_FAB2RAM_D0_O3),
    .FAB2RAM_D1_O0(Tile_X8Y5_FAB2RAM_D1_O0),
    .FAB2RAM_D1_O1(Tile_X8Y5_FAB2RAM_D1_O1),
    .FAB2RAM_D1_O2(Tile_X8Y5_FAB2RAM_D1_O2),
    .FAB2RAM_D1_O3(Tile_X8Y5_FAB2RAM_D1_O3),
    .FAB2RAM_D2_O0(Tile_X8Y5_FAB2RAM_D2_O0),
    .FAB2RAM_D2_O1(Tile_X8Y5_FAB2RAM_D2_O1),
    .FAB2RAM_D2_O2(Tile_X8Y5_FAB2RAM_D2_O2),
    .FAB2RAM_D2_O3(Tile_X8Y5_FAB2RAM_D2_O3),
    .FAB2RAM_D3_O0(Tile_X8Y5_FAB2RAM_D3_O0),
    .FAB2RAM_D3_O1(Tile_X8Y5_FAB2RAM_D3_O1),
    .FAB2RAM_D3_O2(Tile_X8Y5_FAB2RAM_D3_O2),
    .FAB2RAM_D3_O3(Tile_X8Y5_FAB2RAM_D3_O3),
    .FAB2RAM_A0_O0(Tile_X8Y5_FAB2RAM_A0_O0),
    .FAB2RAM_A0_O1(Tile_X8Y5_FAB2RAM_A0_O1),
    .FAB2RAM_A0_O2(Tile_X8Y5_FAB2RAM_A0_O2),
    .FAB2RAM_A0_O3(Tile_X8Y5_FAB2RAM_A0_O3),
    .FAB2RAM_A1_O0(Tile_X8Y5_FAB2RAM_A1_O0),
    .FAB2RAM_A1_O1(Tile_X8Y5_FAB2RAM_A1_O1),
    .FAB2RAM_A1_O2(Tile_X8Y5_FAB2RAM_A1_O2),
    .FAB2RAM_A1_O3(Tile_X8Y5_FAB2RAM_A1_O3),
    .FAB2RAM_C_O0(Tile_X8Y5_FAB2RAM_C_O0),
    .FAB2RAM_C_O1(Tile_X8Y5_FAB2RAM_C_O1),
    .FAB2RAM_C_O2(Tile_X8Y5_FAB2RAM_C_O2),
    .FAB2RAM_C_O3(Tile_X8Y5_FAB2RAM_C_O3),
    .Config_accessC_bit0(Tile_X8Y5_Config_accessC_bit0),
    .Config_accessC_bit1(Tile_X8Y5_Config_accessC_bit1),
    .Config_accessC_bit2(Tile_X8Y5_Config_accessC_bit2),
    .Config_accessC_bit3(Tile_X8Y5_Config_accessC_bit3),
    .UserCLK(Tile_X8Y6_UserCLKo),
    .UserCLKo(Tile_X8Y5_UserCLKo),
    .FrameData(Tile_X7Y5_FrameData_O),
    .FrameData_O(Tile_X8Y5_FrameData_O),
    .FrameStrobe(Tile_X8Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y6_Emulate_Bitstream)
    )
`endif
    Tile_X0Y6_W_IO
    (
    .W1END(Tile_X1Y6_W1BEG),
    .W2MID(Tile_X1Y6_W2BEG),
    .W2END(Tile_X1Y6_W2BEGb),
    .WW4END(Tile_X1Y6_WW4BEG),
    .W6END(Tile_X1Y6_W6BEG),
    .E1BEG(Tile_X0Y6_E1BEG),
    .E2BEG(Tile_X0Y6_E2BEG),
    .E2BEGb(Tile_X0Y6_E2BEGb),
    .EE4BEG(Tile_X0Y6_EE4BEG),
    .E6BEG(Tile_X0Y6_E6BEG),
    .A_O_top(Tile_X0Y6_A_O_top),
    .A_I_top(Tile_X0Y6_A_I_top),
    .A_T_top(Tile_X0Y6_A_T_top),
    .B_O_top(Tile_X0Y6_B_O_top),
    .B_I_top(Tile_X0Y6_B_I_top),
    .B_T_top(Tile_X0Y6_B_T_top),
    .A_config_C_bit0(Tile_X0Y6_A_config_C_bit0),
    .A_config_C_bit1(Tile_X0Y6_A_config_C_bit1),
    .A_config_C_bit2(Tile_X0Y6_A_config_C_bit2),
    .A_config_C_bit3(Tile_X0Y6_A_config_C_bit3),
    .B_config_C_bit0(Tile_X0Y6_B_config_C_bit0),
    .B_config_C_bit1(Tile_X0Y6_B_config_C_bit1),
    .B_config_C_bit2(Tile_X0Y6_B_config_C_bit2),
    .B_config_C_bit3(Tile_X0Y6_B_config_C_bit3),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X0Y6_UserCLKo),
    .FrameData(Tile_Y6_FrameData),
    .FrameData_O(Tile_X0Y6_FrameData_O),
    .FrameStrobe(Tile_X0_FrameStrobe),
    .FrameStrobe_O(Tile_X0Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y6_Emulate_Bitstream)
    )
`endif
    Tile_X1Y6_LUT4AB
    (
    .N1END(Tile_X1Y7_N1BEG),
    .N2MID(Tile_X1Y7_N2BEG),
    .N2END(Tile_X1Y7_N2BEGb),
    .N4END(Tile_X1Y7_N4BEG),
    .NN4END(Tile_X1Y7_NN4BEG),
    .Ci(Tile_X1Y7_Co),
    .E1END(Tile_X0Y6_E1BEG),
    .E2MID(Tile_X0Y6_E2BEG),
    .E2END(Tile_X0Y6_E2BEGb),
    .EE4END(Tile_X0Y6_EE4BEG),
    .E6END(Tile_X0Y6_E6BEG),
    .S1END(Tile_X1Y5_S1BEG),
    .S2MID(Tile_X1Y5_S2BEG),
    .S2END(Tile_X1Y5_S2BEGb),
    .S4END(Tile_X1Y5_S4BEG),
    .SS4END(Tile_X1Y5_SS4BEG),
    .W1END(Tile_X2Y6_W1BEG),
    .W2MID(Tile_X2Y6_W2BEG),
    .W2END(Tile_X2Y6_W2BEGb),
    .WW4END(Tile_X2Y6_WW4BEG),
    .W6END(Tile_X2Y6_W6BEG),
    .N1BEG(Tile_X1Y6_N1BEG),
    .N2BEG(Tile_X1Y6_N2BEG),
    .N2BEGb(Tile_X1Y6_N2BEGb),
    .N4BEG(Tile_X1Y6_N4BEG),
    .NN4BEG(Tile_X1Y6_NN4BEG),
    .Co(Tile_X1Y6_Co),
    .E1BEG(Tile_X1Y6_E1BEG),
    .E2BEG(Tile_X1Y6_E2BEG),
    .E2BEGb(Tile_X1Y6_E2BEGb),
    .EE4BEG(Tile_X1Y6_EE4BEG),
    .E6BEG(Tile_X1Y6_E6BEG),
    .S1BEG(Tile_X1Y6_S1BEG),
    .S2BEG(Tile_X1Y6_S2BEG),
    .S2BEGb(Tile_X1Y6_S2BEGb),
    .S4BEG(Tile_X1Y6_S4BEG),
    .SS4BEG(Tile_X1Y6_SS4BEG),
    .W1BEG(Tile_X1Y6_W1BEG),
    .W2BEG(Tile_X1Y6_W2BEG),
    .W2BEGb(Tile_X1Y6_W2BEGb),
    .WW4BEG(Tile_X1Y6_WW4BEG),
    .W6BEG(Tile_X1Y6_W6BEG),
    .UserCLK(Tile_X1Y7_UserCLKo),
    .UserCLKo(Tile_X1Y6_UserCLKo),
    .FrameData(Tile_X0Y6_FrameData_O),
    .FrameData_O(Tile_X1Y6_FrameData_O),
    .FrameStrobe(Tile_X1Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y6_Emulate_Bitstream)
    )
`endif
    Tile_X2Y6_LUT4AB
    (
    .N1END(Tile_X2Y7_N1BEG),
    .N2MID(Tile_X2Y7_N2BEG),
    .N2END(Tile_X2Y7_N2BEGb),
    .N4END(Tile_X2Y7_N4BEG),
    .NN4END(Tile_X2Y7_NN4BEG),
    .Ci(Tile_X2Y7_Co),
    .E1END(Tile_X1Y6_E1BEG),
    .E2MID(Tile_X1Y6_E2BEG),
    .E2END(Tile_X1Y6_E2BEGb),
    .EE4END(Tile_X1Y6_EE4BEG),
    .E6END(Tile_X1Y6_E6BEG),
    .S1END(Tile_X2Y5_S1BEG),
    .S2MID(Tile_X2Y5_S2BEG),
    .S2END(Tile_X2Y5_S2BEGb),
    .S4END(Tile_X2Y5_S4BEG),
    .SS4END(Tile_X2Y5_SS4BEG),
    .W1END(Tile_X3Y6_W1BEG),
    .W2MID(Tile_X3Y6_W2BEG),
    .W2END(Tile_X3Y6_W2BEGb),
    .WW4END(Tile_X3Y6_WW4BEG),
    .W6END(Tile_X3Y6_W6BEG),
    .N1BEG(Tile_X2Y6_N1BEG),
    .N2BEG(Tile_X2Y6_N2BEG),
    .N2BEGb(Tile_X2Y6_N2BEGb),
    .N4BEG(Tile_X2Y6_N4BEG),
    .NN4BEG(Tile_X2Y6_NN4BEG),
    .Co(Tile_X2Y6_Co),
    .E1BEG(Tile_X2Y6_E1BEG),
    .E2BEG(Tile_X2Y6_E2BEG),
    .E2BEGb(Tile_X2Y6_E2BEGb),
    .EE4BEG(Tile_X2Y6_EE4BEG),
    .E6BEG(Tile_X2Y6_E6BEG),
    .S1BEG(Tile_X2Y6_S1BEG),
    .S2BEG(Tile_X2Y6_S2BEG),
    .S2BEGb(Tile_X2Y6_S2BEGb),
    .S4BEG(Tile_X2Y6_S4BEG),
    .SS4BEG(Tile_X2Y6_SS4BEG),
    .W1BEG(Tile_X2Y6_W1BEG),
    .W2BEG(Tile_X2Y6_W2BEG),
    .W2BEGb(Tile_X2Y6_W2BEGb),
    .WW4BEG(Tile_X2Y6_WW4BEG),
    .W6BEG(Tile_X2Y6_W6BEG),
    .UserCLK(Tile_X2Y7_UserCLKo),
    .UserCLKo(Tile_X2Y6_UserCLKo),
    .FrameData(Tile_X1Y6_FrameData_O),
    .FrameData_O(Tile_X2Y6_FrameData_O),
    .FrameStrobe(Tile_X2Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y6_Emulate_Bitstream)
    )
`endif
    Tile_X3Y6_LUT4AB
    (
    .N1END(Tile_X3Y7_N1BEG),
    .N2MID(Tile_X3Y7_N2BEG),
    .N2END(Tile_X3Y7_N2BEGb),
    .N4END(Tile_X3Y7_N4BEG),
    .NN4END(Tile_X3Y7_NN4BEG),
    .Ci(Tile_X3Y7_Co),
    .E1END(Tile_X2Y6_E1BEG),
    .E2MID(Tile_X2Y6_E2BEG),
    .E2END(Tile_X2Y6_E2BEGb),
    .EE4END(Tile_X2Y6_EE4BEG),
    .E6END(Tile_X2Y6_E6BEG),
    .S1END(Tile_X3Y5_S1BEG),
    .S2MID(Tile_X3Y5_S2BEG),
    .S2END(Tile_X3Y5_S2BEGb),
    .S4END(Tile_X3Y5_S4BEG),
    .SS4END(Tile_X3Y5_SS4BEG),
    .W1END(Tile_X4Y6_W1BEG),
    .W2MID(Tile_X4Y6_W2BEG),
    .W2END(Tile_X4Y6_W2BEGb),
    .WW4END(Tile_X4Y6_WW4BEG),
    .W6END(Tile_X4Y6_W6BEG),
    .N1BEG(Tile_X3Y6_N1BEG),
    .N2BEG(Tile_X3Y6_N2BEG),
    .N2BEGb(Tile_X3Y6_N2BEGb),
    .N4BEG(Tile_X3Y6_N4BEG),
    .NN4BEG(Tile_X3Y6_NN4BEG),
    .Co(Tile_X3Y6_Co),
    .E1BEG(Tile_X3Y6_E1BEG),
    .E2BEG(Tile_X3Y6_E2BEG),
    .E2BEGb(Tile_X3Y6_E2BEGb),
    .EE4BEG(Tile_X3Y6_EE4BEG),
    .E6BEG(Tile_X3Y6_E6BEG),
    .S1BEG(Tile_X3Y6_S1BEG),
    .S2BEG(Tile_X3Y6_S2BEG),
    .S2BEGb(Tile_X3Y6_S2BEGb),
    .S4BEG(Tile_X3Y6_S4BEG),
    .SS4BEG(Tile_X3Y6_SS4BEG),
    .W1BEG(Tile_X3Y6_W1BEG),
    .W2BEG(Tile_X3Y6_W2BEG),
    .W2BEGb(Tile_X3Y6_W2BEGb),
    .WW4BEG(Tile_X3Y6_WW4BEG),
    .W6BEG(Tile_X3Y6_W6BEG),
    .UserCLK(Tile_X3Y7_UserCLKo),
    .UserCLKo(Tile_X3Y6_UserCLKo),
    .FrameData(Tile_X2Y6_FrameData_O),
    .FrameData_O(Tile_X3Y6_FrameData_O),
    .FrameStrobe(Tile_X3Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y6_Emulate_Bitstream)
    )
`endif
    Tile_X4Y6_LUT4AB
    (
    .N1END(Tile_X4Y7_N1BEG),
    .N2MID(Tile_X4Y7_N2BEG),
    .N2END(Tile_X4Y7_N2BEGb),
    .N4END(Tile_X4Y7_N4BEG),
    .NN4END(Tile_X4Y7_NN4BEG),
    .Ci(Tile_X4Y7_Co),
    .E1END(Tile_X3Y6_E1BEG),
    .E2MID(Tile_X3Y6_E2BEG),
    .E2END(Tile_X3Y6_E2BEGb),
    .EE4END(Tile_X3Y6_EE4BEG),
    .E6END(Tile_X3Y6_E6BEG),
    .S1END(Tile_X4Y5_S1BEG),
    .S2MID(Tile_X4Y5_S2BEG),
    .S2END(Tile_X4Y5_S2BEGb),
    .S4END(Tile_X4Y5_S4BEG),
    .SS4END(Tile_X4Y5_SS4BEG),
    .W1END(Tile_X5Y6_W1BEG),
    .W2MID(Tile_X5Y6_W2BEG),
    .W2END(Tile_X5Y6_W2BEGb),
    .WW4END(Tile_X5Y6_WW4BEG),
    .W6END(Tile_X5Y6_W6BEG),
    .N1BEG(Tile_X4Y6_N1BEG),
    .N2BEG(Tile_X4Y6_N2BEG),
    .N2BEGb(Tile_X4Y6_N2BEGb),
    .N4BEG(Tile_X4Y6_N4BEG),
    .NN4BEG(Tile_X4Y6_NN4BEG),
    .Co(Tile_X4Y6_Co),
    .E1BEG(Tile_X4Y6_E1BEG),
    .E2BEG(Tile_X4Y6_E2BEG),
    .E2BEGb(Tile_X4Y6_E2BEGb),
    .EE4BEG(Tile_X4Y6_EE4BEG),
    .E6BEG(Tile_X4Y6_E6BEG),
    .S1BEG(Tile_X4Y6_S1BEG),
    .S2BEG(Tile_X4Y6_S2BEG),
    .S2BEGb(Tile_X4Y6_S2BEGb),
    .S4BEG(Tile_X4Y6_S4BEG),
    .SS4BEG(Tile_X4Y6_SS4BEG),
    .W1BEG(Tile_X4Y6_W1BEG),
    .W2BEG(Tile_X4Y6_W2BEG),
    .W2BEGb(Tile_X4Y6_W2BEGb),
    .WW4BEG(Tile_X4Y6_WW4BEG),
    .W6BEG(Tile_X4Y6_W6BEG),
    .UserCLK(Tile_X4Y7_UserCLKo),
    .UserCLKo(Tile_X4Y6_UserCLKo),
    .FrameData(Tile_X3Y6_FrameData_O),
    .FrameData_O(Tile_X4Y6_FrameData_O),
    .FrameStrobe(Tile_X4Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y6_Emulate_Bitstream)
    )
`endif
    Tile_X5Y6_LUT4AB
    (
    .N1END(Tile_X5Y7_N1BEG),
    .N2MID(Tile_X5Y7_N2BEG),
    .N2END(Tile_X5Y7_N2BEGb),
    .N4END(Tile_X5Y7_N4BEG),
    .NN4END(Tile_X5Y7_NN4BEG),
    .Ci(Tile_X5Y7_Co),
    .E1END(Tile_X4Y6_E1BEG),
    .E2MID(Tile_X4Y6_E2BEG),
    .E2END(Tile_X4Y6_E2BEGb),
    .EE4END(Tile_X4Y6_EE4BEG),
    .E6END(Tile_X4Y6_E6BEG),
    .S1END(Tile_X5Y5_S1BEG),
    .S2MID(Tile_X5Y5_S2BEG),
    .S2END(Tile_X5Y5_S2BEGb),
    .S4END(Tile_X5Y5_S4BEG),
    .SS4END(Tile_X5Y5_SS4BEG),
    .W1END(Tile_X6Y6_W1BEG),
    .W2MID(Tile_X6Y6_W2BEG),
    .W2END(Tile_X6Y6_W2BEGb),
    .WW4END(Tile_X6Y6_WW4BEG),
    .W6END(Tile_X6Y6_W6BEG),
    .N1BEG(Tile_X5Y6_N1BEG),
    .N2BEG(Tile_X5Y6_N2BEG),
    .N2BEGb(Tile_X5Y6_N2BEGb),
    .N4BEG(Tile_X5Y6_N4BEG),
    .NN4BEG(Tile_X5Y6_NN4BEG),
    .Co(Tile_X5Y6_Co),
    .E1BEG(Tile_X5Y6_E1BEG),
    .E2BEG(Tile_X5Y6_E2BEG),
    .E2BEGb(Tile_X5Y6_E2BEGb),
    .EE4BEG(Tile_X5Y6_EE4BEG),
    .E6BEG(Tile_X5Y6_E6BEG),
    .S1BEG(Tile_X5Y6_S1BEG),
    .S2BEG(Tile_X5Y6_S2BEG),
    .S2BEGb(Tile_X5Y6_S2BEGb),
    .S4BEG(Tile_X5Y6_S4BEG),
    .SS4BEG(Tile_X5Y6_SS4BEG),
    .W1BEG(Tile_X5Y6_W1BEG),
    .W2BEG(Tile_X5Y6_W2BEG),
    .W2BEGb(Tile_X5Y6_W2BEGb),
    .WW4BEG(Tile_X5Y6_WW4BEG),
    .W6BEG(Tile_X5Y6_W6BEG),
    .UserCLK(Tile_X5Y7_UserCLKo),
    .UserCLKo(Tile_X5Y6_UserCLKo),
    .FrameData(Tile_X4Y6_FrameData_O),
    .FrameData_O(Tile_X5Y6_FrameData_O),
    .FrameStrobe(Tile_X5Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X6Y6_Emulate_Bitstream)
    )
`endif
    Tile_X6Y6_LUT4AB
    (
    .N1END(Tile_X6Y7_N1BEG),
    .N2MID(Tile_X6Y7_N2BEG),
    .N2END(Tile_X6Y7_N2BEGb),
    .N4END(Tile_X6Y7_N4BEG),
    .NN4END(Tile_X6Y7_NN4BEG),
    .Ci(Tile_X6Y7_Co),
    .E1END(Tile_X5Y6_E1BEG),
    .E2MID(Tile_X5Y6_E2BEG),
    .E2END(Tile_X5Y6_E2BEGb),
    .EE4END(Tile_X5Y6_EE4BEG),
    .E6END(Tile_X5Y6_E6BEG),
    .S1END(Tile_X6Y5_S1BEG),
    .S2MID(Tile_X6Y5_S2BEG),
    .S2END(Tile_X6Y5_S2BEGb),
    .S4END(Tile_X6Y5_S4BEG),
    .SS4END(Tile_X6Y5_SS4BEG),
    .W1END(Tile_X7Y6_W1BEG),
    .W2MID(Tile_X7Y6_W2BEG),
    .W2END(Tile_X7Y6_W2BEGb),
    .WW4END(Tile_X7Y6_WW4BEG),
    .W6END(Tile_X7Y6_W6BEG),
    .N1BEG(Tile_X6Y6_N1BEG),
    .N2BEG(Tile_X6Y6_N2BEG),
    .N2BEGb(Tile_X6Y6_N2BEGb),
    .N4BEG(Tile_X6Y6_N4BEG),
    .NN4BEG(Tile_X6Y6_NN4BEG),
    .Co(Tile_X6Y6_Co),
    .E1BEG(Tile_X6Y6_E1BEG),
    .E2BEG(Tile_X6Y6_E2BEG),
    .E2BEGb(Tile_X6Y6_E2BEGb),
    .EE4BEG(Tile_X6Y6_EE4BEG),
    .E6BEG(Tile_X6Y6_E6BEG),
    .S1BEG(Tile_X6Y6_S1BEG),
    .S2BEG(Tile_X6Y6_S2BEG),
    .S2BEGb(Tile_X6Y6_S2BEGb),
    .S4BEG(Tile_X6Y6_S4BEG),
    .SS4BEG(Tile_X6Y6_SS4BEG),
    .W1BEG(Tile_X6Y6_W1BEG),
    .W2BEG(Tile_X6Y6_W2BEG),
    .W2BEGb(Tile_X6Y6_W2BEGb),
    .WW4BEG(Tile_X6Y6_WW4BEG),
    .W6BEG(Tile_X6Y6_W6BEG),
    .UserCLK(Tile_X6Y7_UserCLKo),
    .UserCLKo(Tile_X6Y6_UserCLKo),
    .FrameData(Tile_X5Y6_FrameData_O),
    .FrameData_O(Tile_X6Y6_FrameData_O),
    .FrameStrobe(Tile_X6Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X6Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X7Y6_Emulate_Bitstream)
    )
`endif
    Tile_X7Y6_LUT4AB
    (
    .N1END(Tile_X7Y7_N1BEG),
    .N2MID(Tile_X7Y7_N2BEG),
    .N2END(Tile_X7Y7_N2BEGb),
    .N4END(Tile_X7Y7_N4BEG),
    .NN4END(Tile_X7Y7_NN4BEG),
    .Ci(Tile_X7Y7_Co),
    .E1END(Tile_X6Y6_E1BEG),
    .E2MID(Tile_X6Y6_E2BEG),
    .E2END(Tile_X6Y6_E2BEGb),
    .EE4END(Tile_X6Y6_EE4BEG),
    .E6END(Tile_X6Y6_E6BEG),
    .S1END(Tile_X7Y5_S1BEG),
    .S2MID(Tile_X7Y5_S2BEG),
    .S2END(Tile_X7Y5_S2BEGb),
    .S4END(Tile_X7Y5_S4BEG),
    .SS4END(Tile_X7Y5_SS4BEG),
    .W1END(Tile_X8Y6_W1BEG),
    .W2MID(Tile_X8Y6_W2BEG),
    .W2END(Tile_X8Y6_W2BEGb),
    .WW4END(Tile_X8Y6_WW4BEG),
    .W6END(Tile_X8Y6_W6BEG),
    .N1BEG(Tile_X7Y6_N1BEG),
    .N2BEG(Tile_X7Y6_N2BEG),
    .N2BEGb(Tile_X7Y6_N2BEGb),
    .N4BEG(Tile_X7Y6_N4BEG),
    .NN4BEG(Tile_X7Y6_NN4BEG),
    .Co(Tile_X7Y6_Co),
    .E1BEG(Tile_X7Y6_E1BEG),
    .E2BEG(Tile_X7Y6_E2BEG),
    .E2BEGb(Tile_X7Y6_E2BEGb),
    .EE4BEG(Tile_X7Y6_EE4BEG),
    .E6BEG(Tile_X7Y6_E6BEG),
    .S1BEG(Tile_X7Y6_S1BEG),
    .S2BEG(Tile_X7Y6_S2BEG),
    .S2BEGb(Tile_X7Y6_S2BEGb),
    .S4BEG(Tile_X7Y6_S4BEG),
    .SS4BEG(Tile_X7Y6_SS4BEG),
    .W1BEG(Tile_X7Y6_W1BEG),
    .W2BEG(Tile_X7Y6_W2BEG),
    .W2BEGb(Tile_X7Y6_W2BEGb),
    .WW4BEG(Tile_X7Y6_WW4BEG),
    .W6BEG(Tile_X7Y6_W6BEG),
    .UserCLK(Tile_X7Y7_UserCLKo),
    .UserCLKo(Tile_X7Y6_UserCLKo),
    .FrameData(Tile_X6Y6_FrameData_O),
    .FrameData_O(Tile_X7Y6_FrameData_O),
    .FrameStrobe(Tile_X7Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X7Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
RAM_IO
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X8Y6_Emulate_Bitstream)
    )
`endif
    Tile_X8Y6_RAM_IO
    (
    .N1END(Tile_X8Y7_N1BEG),
    .N2MID(Tile_X8Y7_N2BEG),
    .N2END(Tile_X8Y7_N2BEGb),
    .N4END(Tile_X8Y7_N4BEG),
    .E1END(Tile_X7Y6_E1BEG),
    .E2MID(Tile_X7Y6_E2BEG),
    .E2END(Tile_X7Y6_E2BEGb),
    .EE4END(Tile_X7Y6_EE4BEG),
    .E6END(Tile_X7Y6_E6BEG),
    .S1END(Tile_X8Y5_S1BEG),
    .S2MID(Tile_X8Y5_S2BEG),
    .S2END(Tile_X8Y5_S2BEGb),
    .S4END(Tile_X8Y5_S4BEG),
    .N1BEG(Tile_X8Y6_N1BEG),
    .N2BEG(Tile_X8Y6_N2BEG),
    .N2BEGb(Tile_X8Y6_N2BEGb),
    .N4BEG(Tile_X8Y6_N4BEG),
    .S1BEG(Tile_X8Y6_S1BEG),
    .S2BEG(Tile_X8Y6_S2BEG),
    .S2BEGb(Tile_X8Y6_S2BEGb),
    .S4BEG(Tile_X8Y6_S4BEG),
    .W1BEG(Tile_X8Y6_W1BEG),
    .W2BEG(Tile_X8Y6_W2BEG),
    .W2BEGb(Tile_X8Y6_W2BEGb),
    .WW4BEG(Tile_X8Y6_WW4BEG),
    .W6BEG(Tile_X8Y6_W6BEG),
    .RAM2FAB_D0_I0(Tile_X8Y6_RAM2FAB_D0_I0),
    .RAM2FAB_D0_I1(Tile_X8Y6_RAM2FAB_D0_I1),
    .RAM2FAB_D0_I2(Tile_X8Y6_RAM2FAB_D0_I2),
    .RAM2FAB_D0_I3(Tile_X8Y6_RAM2FAB_D0_I3),
    .RAM2FAB_D1_I0(Tile_X8Y6_RAM2FAB_D1_I0),
    .RAM2FAB_D1_I1(Tile_X8Y6_RAM2FAB_D1_I1),
    .RAM2FAB_D1_I2(Tile_X8Y6_RAM2FAB_D1_I2),
    .RAM2FAB_D1_I3(Tile_X8Y6_RAM2FAB_D1_I3),
    .RAM2FAB_D2_I0(Tile_X8Y6_RAM2FAB_D2_I0),
    .RAM2FAB_D2_I1(Tile_X8Y6_RAM2FAB_D2_I1),
    .RAM2FAB_D2_I2(Tile_X8Y6_RAM2FAB_D2_I2),
    .RAM2FAB_D2_I3(Tile_X8Y6_RAM2FAB_D2_I3),
    .RAM2FAB_D3_I0(Tile_X8Y6_RAM2FAB_D3_I0),
    .RAM2FAB_D3_I1(Tile_X8Y6_RAM2FAB_D3_I1),
    .RAM2FAB_D3_I2(Tile_X8Y6_RAM2FAB_D3_I2),
    .RAM2FAB_D3_I3(Tile_X8Y6_RAM2FAB_D3_I3),
    .FAB2RAM_D0_O0(Tile_X8Y6_FAB2RAM_D0_O0),
    .FAB2RAM_D0_O1(Tile_X8Y6_FAB2RAM_D0_O1),
    .FAB2RAM_D0_O2(Tile_X8Y6_FAB2RAM_D0_O2),
    .FAB2RAM_D0_O3(Tile_X8Y6_FAB2RAM_D0_O3),
    .FAB2RAM_D1_O0(Tile_X8Y6_FAB2RAM_D1_O0),
    .FAB2RAM_D1_O1(Tile_X8Y6_FAB2RAM_D1_O1),
    .FAB2RAM_D1_O2(Tile_X8Y6_FAB2RAM_D1_O2),
    .FAB2RAM_D1_O3(Tile_X8Y6_FAB2RAM_D1_O3),
    .FAB2RAM_D2_O0(Tile_X8Y6_FAB2RAM_D2_O0),
    .FAB2RAM_D2_O1(Tile_X8Y6_FAB2RAM_D2_O1),
    .FAB2RAM_D2_O2(Tile_X8Y6_FAB2RAM_D2_O2),
    .FAB2RAM_D2_O3(Tile_X8Y6_FAB2RAM_D2_O3),
    .FAB2RAM_D3_O0(Tile_X8Y6_FAB2RAM_D3_O0),
    .FAB2RAM_D3_O1(Tile_X8Y6_FAB2RAM_D3_O1),
    .FAB2RAM_D3_O2(Tile_X8Y6_FAB2RAM_D3_O2),
    .FAB2RAM_D3_O3(Tile_X8Y6_FAB2RAM_D3_O3),
    .FAB2RAM_A0_O0(Tile_X8Y6_FAB2RAM_A0_O0),
    .FAB2RAM_A0_O1(Tile_X8Y6_FAB2RAM_A0_O1),
    .FAB2RAM_A0_O2(Tile_X8Y6_FAB2RAM_A0_O2),
    .FAB2RAM_A0_O3(Tile_X8Y6_FAB2RAM_A0_O3),
    .FAB2RAM_A1_O0(Tile_X8Y6_FAB2RAM_A1_O0),
    .FAB2RAM_A1_O1(Tile_X8Y6_FAB2RAM_A1_O1),
    .FAB2RAM_A1_O2(Tile_X8Y6_FAB2RAM_A1_O2),
    .FAB2RAM_A1_O3(Tile_X8Y6_FAB2RAM_A1_O3),
    .FAB2RAM_C_O0(Tile_X8Y6_FAB2RAM_C_O0),
    .FAB2RAM_C_O1(Tile_X8Y6_FAB2RAM_C_O1),
    .FAB2RAM_C_O2(Tile_X8Y6_FAB2RAM_C_O2),
    .FAB2RAM_C_O3(Tile_X8Y6_FAB2RAM_C_O3),
    .Config_accessC_bit0(Tile_X8Y6_Config_accessC_bit0),
    .Config_accessC_bit1(Tile_X8Y6_Config_accessC_bit1),
    .Config_accessC_bit2(Tile_X8Y6_Config_accessC_bit2),
    .Config_accessC_bit3(Tile_X8Y6_Config_accessC_bit3),
    .UserCLK(Tile_X8Y7_UserCLKo),
    .UserCLKo(Tile_X8Y6_UserCLKo),
    .FrameData(Tile_X7Y6_FrameData_O),
    .FrameData_O(Tile_X8Y6_FrameData_O),
    .FrameStrobe(Tile_X8Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X8Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X1Y7_S_term_single (
    .S1END(Tile_X1Y6_S1BEG),
    .S2MID(Tile_X1Y6_S2BEG),
    .S2END(Tile_X1Y6_S2BEGb),
    .S4END(Tile_X1Y6_S4BEG),
    .SS4END(Tile_X1Y6_SS4BEG),
    .N1BEG(Tile_X1Y7_N1BEG),
    .N2BEG(Tile_X1Y7_N2BEG),
    .N2BEGb(Tile_X1Y7_N2BEGb),
    .N4BEG(Tile_X1Y7_N4BEG),
    .NN4BEG(Tile_X1Y7_NN4BEG),
    .Co(Tile_X1Y7_Co),
    .UIO_BOT_UIN0(Tile_X1Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X1Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X1Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X1Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X1Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X1Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X1Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X1Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X1Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X1Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X1Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X1Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X1Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X1Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X1Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X1Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X1Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X1Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X1Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X1Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X1Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X1Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X1Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X1Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X1Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X1Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X1Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X1Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X1Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X1Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X1Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X1Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X1Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X1Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X1Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X1Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X1Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X1Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X1Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X1Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X1Y7_UserCLKo),
    .FrameStrobe(Tile_X1_FrameStrobe),
    .FrameStrobe_O(Tile_X1Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X2Y7_S_term_single (
    .S1END(Tile_X2Y6_S1BEG),
    .S2MID(Tile_X2Y6_S2BEG),
    .S2END(Tile_X2Y6_S2BEGb),
    .S4END(Tile_X2Y6_S4BEG),
    .SS4END(Tile_X2Y6_SS4BEG),
    .N1BEG(Tile_X2Y7_N1BEG),
    .N2BEG(Tile_X2Y7_N2BEG),
    .N2BEGb(Tile_X2Y7_N2BEGb),
    .N4BEG(Tile_X2Y7_N4BEG),
    .NN4BEG(Tile_X2Y7_NN4BEG),
    .Co(Tile_X2Y7_Co),
    .UIO_BOT_UIN0(Tile_X2Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X2Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X2Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X2Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X2Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X2Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X2Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X2Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X2Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X2Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X2Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X2Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X2Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X2Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X2Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X2Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X2Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X2Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X2Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X2Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X2Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X2Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X2Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X2Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X2Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X2Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X2Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X2Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X2Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X2Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X2Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X2Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X2Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X2Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X2Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X2Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X2Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X2Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X2Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X2Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X2Y7_UserCLKo),
    .FrameStrobe(Tile_X2_FrameStrobe),
    .FrameStrobe_O(Tile_X2Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X3Y7_S_term_single (
    .S1END(Tile_X3Y6_S1BEG),
    .S2MID(Tile_X3Y6_S2BEG),
    .S2END(Tile_X3Y6_S2BEGb),
    .S4END(Tile_X3Y6_S4BEG),
    .SS4END(Tile_X3Y6_SS4BEG),
    .N1BEG(Tile_X3Y7_N1BEG),
    .N2BEG(Tile_X3Y7_N2BEG),
    .N2BEGb(Tile_X3Y7_N2BEGb),
    .N4BEG(Tile_X3Y7_N4BEG),
    .NN4BEG(Tile_X3Y7_NN4BEG),
    .Co(Tile_X3Y7_Co),
    .UIO_BOT_UIN0(Tile_X3Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X3Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X3Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X3Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X3Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X3Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X3Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X3Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X3Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X3Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X3Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X3Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X3Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X3Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X3Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X3Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X3Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X3Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X3Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X3Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X3Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X3Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X3Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X3Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X3Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X3Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X3Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X3Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X3Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X3Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X3Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X3Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X3Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X3Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X3Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X3Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X3Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X3Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X3Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X3Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X3Y7_UserCLKo),
    .FrameStrobe(Tile_X3_FrameStrobe),
    .FrameStrobe_O(Tile_X3Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X4Y7_S_term_single (
    .S1END(Tile_X4Y6_S1BEG),
    .S2MID(Tile_X4Y6_S2BEG),
    .S2END(Tile_X4Y6_S2BEGb),
    .S4END(Tile_X4Y6_S4BEG),
    .SS4END(Tile_X4Y6_SS4BEG),
    .N1BEG(Tile_X4Y7_N1BEG),
    .N2BEG(Tile_X4Y7_N2BEG),
    .N2BEGb(Tile_X4Y7_N2BEGb),
    .N4BEG(Tile_X4Y7_N4BEG),
    .NN4BEG(Tile_X4Y7_NN4BEG),
    .Co(Tile_X4Y7_Co),
    .UIO_BOT_UIN0(Tile_X4Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X4Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X4Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X4Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X4Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X4Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X4Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X4Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X4Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X4Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X4Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X4Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X4Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X4Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X4Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X4Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X4Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X4Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X4Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X4Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X4Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X4Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X4Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X4Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X4Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X4Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X4Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X4Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X4Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X4Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X4Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X4Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X4Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X4Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X4Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X4Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X4Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X4Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X4Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X4Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X4Y7_UserCLKo),
    .FrameStrobe(Tile_X4_FrameStrobe),
    .FrameStrobe_O(Tile_X4Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X5Y7_S_term_single (
    .S1END(Tile_X5Y6_S1BEG),
    .S2MID(Tile_X5Y6_S2BEG),
    .S2END(Tile_X5Y6_S2BEGb),
    .S4END(Tile_X5Y6_S4BEG),
    .SS4END(Tile_X5Y6_SS4BEG),
    .N1BEG(Tile_X5Y7_N1BEG),
    .N2BEG(Tile_X5Y7_N2BEG),
    .N2BEGb(Tile_X5Y7_N2BEGb),
    .N4BEG(Tile_X5Y7_N4BEG),
    .NN4BEG(Tile_X5Y7_NN4BEG),
    .Co(Tile_X5Y7_Co),
    .UIO_BOT_UIN0(Tile_X5Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X5Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X5Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X5Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X5Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X5Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X5Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X5Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X5Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X5Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X5Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X5Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X5Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X5Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X5Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X5Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X5Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X5Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X5Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X5Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X5Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X5Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X5Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X5Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X5Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X5Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X5Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X5Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X5Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X5Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X5Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X5Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X5Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X5Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X5Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X5Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X5Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X5Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X5Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X5Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X5Y7_UserCLKo),
    .FrameStrobe(Tile_X5_FrameStrobe),
    .FrameStrobe_O(Tile_X5Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X6Y7_S_term_single (
    .S1END(Tile_X6Y6_S1BEG),
    .S2MID(Tile_X6Y6_S2BEG),
    .S2END(Tile_X6Y6_S2BEGb),
    .S4END(Tile_X6Y6_S4BEG),
    .SS4END(Tile_X6Y6_SS4BEG),
    .N1BEG(Tile_X6Y7_N1BEG),
    .N2BEG(Tile_X6Y7_N2BEG),
    .N2BEGb(Tile_X6Y7_N2BEGb),
    .N4BEG(Tile_X6Y7_N4BEG),
    .NN4BEG(Tile_X6Y7_NN4BEG),
    .Co(Tile_X6Y7_Co),
    .UIO_BOT_UIN0(Tile_X6Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X6Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X6Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X6Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X6Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X6Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X6Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X6Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X6Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X6Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X6Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X6Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X6Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X6Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X6Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X6Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X6Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X6Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X6Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X6Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X6Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X6Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X6Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X6Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X6Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X6Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X6Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X6Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X6Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X6Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X6Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X6Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X6Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X6Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X6Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X6Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X6Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X6Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X6Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X6Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X6Y7_UserCLKo),
    .FrameStrobe(Tile_X6_FrameStrobe),
    .FrameStrobe_O(Tile_X6Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_single Tile_X7Y7_S_term_single (
    .S1END(Tile_X7Y6_S1BEG),
    .S2MID(Tile_X7Y6_S2BEG),
    .S2END(Tile_X7Y6_S2BEGb),
    .S4END(Tile_X7Y6_S4BEG),
    .SS4END(Tile_X7Y6_SS4BEG),
    .N1BEG(Tile_X7Y7_N1BEG),
    .N2BEG(Tile_X7Y7_N2BEG),
    .N2BEGb(Tile_X7Y7_N2BEGb),
    .N4BEG(Tile_X7Y7_N4BEG),
    .NN4BEG(Tile_X7Y7_NN4BEG),
    .Co(Tile_X7Y7_Co),
    .UIO_BOT_UIN0(Tile_X7Y7_UIO_BOT_UIN0),
    .UIO_BOT_UIN1(Tile_X7Y7_UIO_BOT_UIN1),
    .UIO_BOT_UIN10(Tile_X7Y7_UIO_BOT_UIN10),
    .UIO_BOT_UIN11(Tile_X7Y7_UIO_BOT_UIN11),
    .UIO_BOT_UIN12(Tile_X7Y7_UIO_BOT_UIN12),
    .UIO_BOT_UIN13(Tile_X7Y7_UIO_BOT_UIN13),
    .UIO_BOT_UIN14(Tile_X7Y7_UIO_BOT_UIN14),
    .UIO_BOT_UIN15(Tile_X7Y7_UIO_BOT_UIN15),
    .UIO_BOT_UIN16(Tile_X7Y7_UIO_BOT_UIN16),
    .UIO_BOT_UIN17(Tile_X7Y7_UIO_BOT_UIN17),
    .UIO_BOT_UIN18(Tile_X7Y7_UIO_BOT_UIN18),
    .UIO_BOT_UIN19(Tile_X7Y7_UIO_BOT_UIN19),
    .UIO_BOT_UIN2(Tile_X7Y7_UIO_BOT_UIN2),
    .UIO_BOT_UIN3(Tile_X7Y7_UIO_BOT_UIN3),
    .UIO_BOT_UIN4(Tile_X7Y7_UIO_BOT_UIN4),
    .UIO_BOT_UIN5(Tile_X7Y7_UIO_BOT_UIN5),
    .UIO_BOT_UIN6(Tile_X7Y7_UIO_BOT_UIN6),
    .UIO_BOT_UIN7(Tile_X7Y7_UIO_BOT_UIN7),
    .UIO_BOT_UIN8(Tile_X7Y7_UIO_BOT_UIN8),
    .UIO_BOT_UIN9(Tile_X7Y7_UIO_BOT_UIN9),
    .UIO_BOT_UOUT0(Tile_X7Y7_UIO_BOT_UOUT0),
    .UIO_BOT_UOUT1(Tile_X7Y7_UIO_BOT_UOUT1),
    .UIO_BOT_UOUT10(Tile_X7Y7_UIO_BOT_UOUT10),
    .UIO_BOT_UOUT11(Tile_X7Y7_UIO_BOT_UOUT11),
    .UIO_BOT_UOUT12(Tile_X7Y7_UIO_BOT_UOUT12),
    .UIO_BOT_UOUT13(Tile_X7Y7_UIO_BOT_UOUT13),
    .UIO_BOT_UOUT14(Tile_X7Y7_UIO_BOT_UOUT14),
    .UIO_BOT_UOUT15(Tile_X7Y7_UIO_BOT_UOUT15),
    .UIO_BOT_UOUT16(Tile_X7Y7_UIO_BOT_UOUT16),
    .UIO_BOT_UOUT17(Tile_X7Y7_UIO_BOT_UOUT17),
    .UIO_BOT_UOUT18(Tile_X7Y7_UIO_BOT_UOUT18),
    .UIO_BOT_UOUT19(Tile_X7Y7_UIO_BOT_UOUT19),
    .UIO_BOT_UOUT2(Tile_X7Y7_UIO_BOT_UOUT2),
    .UIO_BOT_UOUT3(Tile_X7Y7_UIO_BOT_UOUT3),
    .UIO_BOT_UOUT4(Tile_X7Y7_UIO_BOT_UOUT4),
    .UIO_BOT_UOUT5(Tile_X7Y7_UIO_BOT_UOUT5),
    .UIO_BOT_UOUT6(Tile_X7Y7_UIO_BOT_UOUT6),
    .UIO_BOT_UOUT7(Tile_X7Y7_UIO_BOT_UOUT7),
    .UIO_BOT_UOUT8(Tile_X7Y7_UIO_BOT_UOUT8),
    .UIO_BOT_UOUT9(Tile_X7Y7_UIO_BOT_UOUT9),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X7Y7_UserCLKo),
    .FrameStrobe(Tile_X7_FrameStrobe),
    .FrameStrobe_O(Tile_X7Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_term_RAM_IO Tile_X8Y7_S_term_RAM_IO (
    .S1END(Tile_X8Y6_S1BEG),
    .S2MID(Tile_X8Y6_S2BEG),
    .S2END(Tile_X8Y6_S2BEGb),
    .S4END(Tile_X8Y6_S4BEG),
    .N1BEG(Tile_X8Y7_N1BEG),
    .N2BEG(Tile_X8Y7_N2BEG),
    .N2BEGb(Tile_X8Y7_N2BEGb),
    .N4BEG(Tile_X8Y7_N4BEG),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X8Y7_UserCLKo),
    .FrameStrobe(Tile_X8_FrameStrobe),
    .FrameStrobe_O(Tile_X8Y7_FrameStrobe_O)
);

endmodule
