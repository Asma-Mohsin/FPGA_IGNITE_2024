magic
tech sky130A
magscale 1 2
timestamp 1732405367
<< viali >>
rect 5457 5321 5491 5355
rect 6745 5321 6779 5355
rect 7481 5321 7515 5355
rect 8033 5321 8067 5355
rect 8585 5321 8619 5355
rect 9505 5321 9539 5355
rect 10609 5321 10643 5355
rect 12081 5321 12115 5355
rect 12633 5321 12667 5355
rect 13737 5321 13771 5355
rect 14657 5321 14691 5355
rect 15209 5321 15243 5355
rect 15761 5321 15795 5355
rect 16313 5321 16347 5355
rect 17233 5321 17267 5355
rect 17785 5321 17819 5355
rect 18337 5321 18371 5355
rect 18889 5321 18923 5355
rect 27537 5321 27571 5355
rect 32873 5321 32907 5355
rect 34897 5321 34931 5355
rect 35449 5321 35483 5355
rect 36001 5321 36035 5355
rect 37473 5321 37507 5355
rect 39129 5321 39163 5355
rect 40601 5321 40635 5355
rect 41153 5321 41187 5355
rect 5549 5253 5583 5287
rect 7573 5253 7607 5287
rect 8125 5253 8159 5287
rect 12173 5253 12207 5287
rect 12725 5253 12759 5287
rect 15853 5253 15887 5287
rect 19349 5253 19383 5287
rect 19901 5253 19935 5287
rect 20453 5253 20487 5287
rect 20821 5253 20855 5287
rect 39957 5253 39991 5287
rect 6101 5185 6135 5219
rect 7021 5185 7055 5219
rect 8677 5185 8711 5219
rect 9597 5185 9631 5219
rect 10149 5185 10183 5219
rect 10701 5185 10735 5219
rect 11253 5185 11287 5219
rect 11713 5185 11747 5219
rect 13277 5185 13311 5219
rect 13829 5185 13863 5219
rect 14749 5185 14783 5219
rect 15301 5185 15335 5219
rect 16423 5185 16457 5219
rect 17325 5185 17359 5219
rect 17877 5185 17911 5219
rect 18429 5185 18463 5219
rect 18981 5185 19015 5219
rect 19717 5185 19751 5219
rect 20269 5185 20303 5219
rect 21373 5185 21407 5219
rect 21649 5185 21683 5219
rect 22017 5185 22051 5219
rect 22293 5185 22327 5219
rect 22569 5185 22603 5219
rect 22845 5185 22879 5219
rect 23121 5185 23155 5219
rect 23397 5185 23431 5219
rect 23673 5185 23707 5219
rect 23949 5185 23983 5219
rect 24225 5185 24259 5219
rect 24593 5185 24627 5219
rect 24869 5185 24903 5219
rect 25145 5209 25179 5243
rect 25421 5185 25455 5219
rect 25697 5185 25731 5219
rect 25789 5185 25823 5219
rect 26065 5185 26099 5219
rect 26341 5185 26375 5219
rect 26617 5185 26651 5219
rect 27169 5185 27203 5219
rect 27445 5185 27479 5219
rect 27721 5185 27755 5219
rect 27997 5185 28031 5219
rect 28273 5185 28307 5219
rect 28549 5185 28583 5219
rect 28825 5185 28859 5219
rect 29101 5185 29135 5219
rect 30113 5185 30147 5219
rect 30389 5185 30423 5219
rect 30665 5185 30699 5219
rect 30941 5185 30975 5219
rect 31217 5185 31251 5219
rect 31493 5185 31527 5219
rect 31769 5185 31803 5219
rect 32137 5185 32171 5219
rect 32413 5185 32447 5219
rect 32689 5185 32723 5219
rect 32965 5185 32999 5219
rect 33241 5185 33275 5219
rect 33517 5185 33551 5219
rect 33793 5185 33827 5219
rect 34253 5185 34287 5219
rect 34529 5185 34563 5219
rect 34805 5185 34839 5219
rect 35357 5185 35391 5219
rect 35909 5185 35943 5219
rect 36461 5185 36495 5219
rect 37381 5185 37415 5219
rect 37933 5185 37967 5219
rect 38485 5185 38519 5219
rect 39037 5185 39071 5219
rect 40509 5185 40543 5219
rect 41061 5185 41095 5219
rect 5825 5117 5859 5151
rect 9873 5117 9907 5151
rect 10977 5117 11011 5151
rect 31401 5049 31435 5083
rect 32597 5049 32631 5083
rect 33149 5049 33183 5083
rect 34069 5049 34103 5083
rect 34345 5049 34379 5083
rect 38669 5049 38703 5083
rect 11529 4981 11563 5015
rect 13185 4981 13219 5015
rect 21189 4981 21223 5015
rect 21465 4981 21499 5015
rect 21833 4981 21867 5015
rect 22109 4981 22143 5015
rect 22385 4981 22419 5015
rect 22661 4981 22695 5015
rect 22937 4981 22971 5015
rect 23213 4981 23247 5015
rect 23489 4981 23523 5015
rect 23765 4981 23799 5015
rect 24041 4981 24075 5015
rect 24409 4981 24443 5015
rect 24685 4981 24719 5015
rect 24961 4981 24995 5015
rect 25237 4981 25271 5015
rect 25513 4981 25547 5015
rect 25973 4981 26007 5015
rect 26249 4981 26283 5015
rect 26525 4981 26559 5015
rect 26801 4981 26835 5015
rect 26985 4981 27019 5015
rect 27261 4981 27295 5015
rect 27813 4981 27847 5015
rect 28089 4981 28123 5015
rect 28365 4981 28399 5015
rect 28641 4981 28675 5015
rect 28917 4981 28951 5015
rect 30297 4981 30331 5015
rect 30573 4981 30607 5015
rect 30849 4981 30883 5015
rect 31125 4981 31159 5015
rect 31677 4981 31711 5015
rect 31953 4981 31987 5015
rect 32321 4981 32355 5015
rect 33425 4981 33459 5015
rect 33701 4981 33735 5015
rect 33977 4981 34011 5015
rect 36553 4981 36587 5015
rect 38025 4981 38059 5015
rect 40049 4981 40083 5015
rect 7297 4777 7331 4811
rect 7849 4777 7883 4811
rect 8401 4777 8435 4811
rect 9321 4777 9355 4811
rect 9873 4777 9907 4811
rect 10425 4777 10459 4811
rect 11069 4777 11103 4811
rect 11437 4777 11471 4811
rect 12081 4777 12115 4811
rect 12449 4777 12483 4811
rect 13001 4777 13035 4811
rect 13553 4777 13587 4811
rect 14197 4777 14231 4811
rect 15945 4777 15979 4811
rect 17509 4777 17543 4811
rect 18153 4777 18187 4811
rect 18705 4777 18739 4811
rect 20729 4777 20763 4811
rect 21741 4777 21775 4811
rect 25789 4777 25823 4811
rect 27629 4777 27663 4811
rect 28457 4777 28491 4811
rect 29009 4777 29043 4811
rect 31677 4777 31711 4811
rect 34437 4777 34471 4811
rect 34805 4777 34839 4811
rect 35265 4777 35299 4811
rect 36093 4777 36127 4811
rect 37197 4777 37231 4811
rect 38301 4777 38335 4811
rect 38853 4777 38887 4811
rect 39405 4777 39439 4811
rect 40049 4777 40083 4811
rect 41153 4777 41187 4811
rect 5733 4709 5767 4743
rect 6285 4709 6319 4743
rect 6837 4709 6871 4743
rect 14841 4709 14875 4743
rect 15393 4709 15427 4743
rect 16497 4709 16531 4743
rect 17049 4709 17083 4743
rect 19349 4709 19383 4743
rect 20177 4709 20211 4743
rect 21373 4709 21407 4743
rect 26341 4709 26375 4743
rect 32045 4709 32079 4743
rect 33057 4709 33091 4743
rect 34161 4709 34195 4743
rect 36737 4709 36771 4743
rect 37841 4709 37875 4743
rect 40693 4709 40727 4743
rect 5917 4573 5951 4607
rect 6469 4573 6503 4607
rect 7021 4573 7055 4607
rect 8125 4573 8159 4607
rect 8677 4573 8711 4607
rect 9965 4573 9999 4607
rect 11345 4573 11379 4607
rect 13829 4573 13863 4607
rect 14473 4573 14507 4607
rect 15025 4573 15059 4607
rect 15577 4573 15611 4607
rect 15853 4573 15887 4607
rect 17785 4573 17819 4607
rect 18061 4573 18095 4607
rect 19533 4573 19567 4607
rect 19809 4573 19843 4607
rect 20077 4573 20111 4607
rect 20361 4573 20395 4607
rect 20637 4573 20671 4607
rect 20913 4573 20947 4607
rect 21189 4573 21223 4607
rect 21557 4573 21591 4607
rect 21925 4573 21959 4607
rect 22201 4573 22235 4607
rect 22477 4573 22511 4607
rect 22845 4573 22879 4607
rect 23121 4573 23155 4607
rect 23397 4573 23431 4607
rect 23673 4573 23707 4607
rect 24041 4573 24075 4607
rect 24593 4573 24627 4607
rect 24869 4573 24903 4607
rect 25145 4573 25179 4607
rect 25421 4573 25455 4607
rect 25697 4573 25731 4607
rect 25973 4573 26007 4607
rect 26157 4573 26191 4607
rect 27813 4573 27847 4607
rect 28089 4573 28123 4607
rect 28365 4573 28399 4607
rect 28641 4573 28675 4607
rect 29193 4573 29227 4607
rect 29929 4573 29963 4607
rect 30849 4573 30883 4607
rect 31217 4573 31251 4607
rect 31493 4573 31527 4607
rect 31861 4573 31895 4607
rect 32229 4573 32263 4607
rect 32873 4573 32907 4607
rect 33977 4573 34011 4607
rect 34253 4573 34287 4607
rect 35081 4573 35115 4607
rect 35357 4573 35391 4607
rect 35633 4573 35667 4607
rect 38209 4573 38243 4607
rect 41061 4573 41095 4607
rect 41521 4573 41555 4607
rect 42073 4573 42107 4607
rect 7573 4505 7607 4539
rect 9413 4505 9447 4539
rect 10517 4505 10551 4539
rect 10793 4505 10827 4539
rect 12173 4505 12207 4539
rect 12725 4505 12759 4539
rect 13277 4505 13311 4539
rect 16681 4505 16715 4539
rect 17233 4505 17267 4539
rect 18613 4505 18647 4539
rect 36001 4505 36035 4539
rect 36553 4505 36587 4539
rect 37105 4505 37139 4539
rect 37657 4505 37691 4539
rect 38761 4505 38795 4539
rect 39313 4505 39347 4539
rect 39957 4505 39991 4539
rect 40509 4505 40543 4539
rect 19625 4437 19659 4471
rect 19901 4437 19935 4471
rect 20453 4437 20487 4471
rect 21005 4437 21039 4471
rect 22017 4437 22051 4471
rect 22293 4437 22327 4471
rect 22661 4437 22695 4471
rect 22937 4437 22971 4471
rect 23213 4437 23247 4471
rect 23489 4437 23523 4471
rect 23857 4437 23891 4471
rect 24409 4437 24443 4471
rect 24685 4437 24719 4471
rect 24961 4437 24995 4471
rect 25237 4437 25271 4471
rect 25513 4437 25547 4471
rect 27905 4437 27939 4471
rect 28181 4437 28215 4471
rect 29745 4437 29779 4471
rect 31033 4437 31067 4471
rect 31401 4437 31435 4471
rect 32413 4437 32447 4471
rect 35541 4437 35575 4471
rect 35817 4437 35851 4471
rect 41705 4437 41739 4471
rect 42257 4437 42291 4471
rect 10885 4233 10919 4267
rect 11161 4233 11195 4267
rect 12173 4233 12207 4267
rect 12633 4233 12667 4267
rect 13553 4233 13587 4267
rect 16037 4233 16071 4267
rect 17049 4233 17083 4267
rect 17785 4233 17819 4267
rect 18061 4233 18095 4267
rect 18613 4233 18647 4267
rect 18889 4233 18923 4267
rect 19165 4233 19199 4267
rect 19533 4233 19567 4267
rect 35909 4233 35943 4267
rect 36185 4233 36219 4267
rect 9229 4165 9263 4199
rect 11805 4165 11839 4199
rect 12541 4165 12575 4199
rect 13277 4165 13311 4199
rect 14013 4165 14047 4199
rect 14381 4165 14415 4199
rect 15025 4165 15059 4199
rect 15485 4165 15519 4199
rect 8861 4097 8895 4131
rect 9689 4097 9723 4131
rect 10057 4097 10091 4131
rect 11069 4097 11103 4131
rect 11345 4097 11379 4131
rect 12357 4097 12391 4131
rect 13001 4097 13035 4131
rect 13737 4097 13771 4131
rect 14657 4097 14691 4131
rect 15669 4097 15703 4131
rect 15945 4097 15979 4131
rect 16221 4097 16255 4131
rect 17233 4097 17267 4131
rect 17969 4097 18003 4131
rect 18245 4097 18279 4131
rect 18521 4097 18555 4131
rect 18797 4097 18831 4131
rect 19073 4097 19107 4131
rect 19349 4097 19383 4131
rect 19717 4097 19751 4131
rect 20453 4097 20487 4131
rect 21005 4097 21039 4131
rect 26433 4097 26467 4131
rect 35449 4097 35483 4131
rect 35725 4097 35759 4131
rect 36001 4097 36035 4131
rect 36277 4097 36311 4131
rect 36553 4097 36587 4131
rect 39129 4097 39163 4131
rect 39865 4097 39899 4131
rect 40601 4097 40635 4131
rect 11989 3961 12023 3995
rect 12817 3961 12851 3995
rect 13461 3961 13495 3995
rect 14197 3961 14231 3995
rect 14565 3961 14599 3995
rect 18337 3961 18371 3995
rect 35633 3961 35667 3995
rect 36461 3961 36495 3995
rect 15761 3893 15795 3927
rect 20269 3893 20303 3927
rect 20821 3893 20855 3927
rect 26617 3893 26651 3927
rect 36737 3893 36771 3927
rect 39313 3893 39347 3927
rect 40049 3893 40083 3927
rect 40785 3893 40819 3927
rect 16129 3689 16163 3723
rect 33793 3689 33827 3723
rect 26893 3621 26927 3655
rect 16313 3485 16347 3519
rect 26709 3485 26743 3519
rect 31677 3485 31711 3519
rect 33609 3485 33643 3519
rect 31493 3349 31527 3383
rect 2605 3145 2639 3179
rect 12725 3145 12759 3179
rect 15577 3145 15611 3179
rect 15853 3145 15887 3179
rect 16313 3145 16347 3179
rect 16865 3145 16899 3179
rect 17141 3145 17175 3179
rect 24225 3145 24259 3179
rect 25329 3145 25363 3179
rect 26985 3145 27019 3179
rect 32413 3145 32447 3179
rect 32965 3145 32999 3179
rect 33241 3145 33275 3179
rect 1501 3009 1535 3043
rect 2513 3009 2547 3043
rect 4169 3009 4203 3043
rect 5457 3009 5491 3043
rect 10333 3009 10367 3043
rect 11069 3009 11103 3043
rect 11253 3009 11287 3043
rect 12909 3009 12943 3043
rect 15761 3009 15795 3043
rect 16037 3009 16071 3043
rect 16221 3009 16255 3043
rect 17049 3009 17083 3043
rect 17325 3009 17359 3043
rect 24041 3009 24075 3043
rect 25513 3009 25547 3043
rect 26249 3009 26283 3043
rect 27169 3009 27203 3043
rect 27721 3009 27755 3043
rect 32229 3009 32263 3043
rect 32689 3009 32723 3043
rect 32781 3009 32815 3043
rect 33057 3009 33091 3043
rect 34805 3009 34839 3043
rect 43637 3009 43671 3043
rect 44189 3009 44223 3043
rect 3893 2941 3927 2975
rect 1685 2873 1719 2907
rect 5641 2873 5675 2907
rect 10517 2873 10551 2907
rect 26065 2805 26099 2839
rect 27537 2805 27571 2839
rect 32505 2805 32539 2839
rect 34989 2805 35023 2839
rect 43913 2805 43947 2839
rect 44281 2805 44315 2839
rect 1869 2601 1903 2635
rect 9965 2601 9999 2635
rect 10701 2601 10735 2635
rect 11713 2601 11747 2635
rect 12173 2601 12207 2635
rect 12909 2601 12943 2635
rect 13645 2601 13679 2635
rect 14381 2601 14415 2635
rect 15117 2601 15151 2635
rect 15853 2601 15887 2635
rect 16681 2601 16715 2635
rect 17141 2601 17175 2635
rect 18613 2601 18647 2635
rect 23029 2601 23063 2635
rect 25973 2601 26007 2635
rect 26985 2601 27019 2635
rect 27445 2601 27479 2635
rect 28181 2601 28215 2635
rect 28917 2601 28951 2635
rect 29653 2601 29687 2635
rect 30389 2601 30423 2635
rect 19349 2533 19383 2567
rect 22293 2533 22327 2567
rect 25237 2533 25271 2567
rect 4721 2465 4755 2499
rect 4445 2397 4479 2431
rect 5917 2397 5951 2431
rect 6193 2397 6227 2431
rect 6837 2397 6871 2431
rect 7113 2397 7147 2431
rect 7757 2397 7791 2431
rect 8309 2397 8343 2431
rect 9045 2397 9079 2431
rect 9781 2397 9815 2431
rect 10517 2397 10551 2431
rect 11529 2397 11563 2431
rect 11989 2397 12023 2431
rect 12725 2397 12759 2431
rect 13461 2397 13495 2431
rect 14197 2397 14231 2431
rect 14933 2397 14967 2431
rect 15669 2397 15703 2431
rect 16865 2397 16899 2431
rect 17325 2397 17359 2431
rect 18061 2397 18095 2431
rect 18797 2397 18831 2431
rect 19533 2397 19567 2431
rect 20269 2397 20303 2431
rect 21005 2397 21039 2431
rect 22017 2397 22051 2431
rect 22477 2397 22511 2431
rect 23213 2397 23247 2431
rect 23949 2397 23983 2431
rect 24685 2397 24719 2431
rect 25421 2397 25455 2431
rect 26157 2397 26191 2431
rect 27169 2397 27203 2431
rect 27629 2397 27663 2431
rect 28365 2397 28399 2431
rect 29101 2397 29135 2431
rect 29837 2397 29871 2431
rect 30573 2397 30607 2431
rect 31493 2397 31527 2431
rect 32505 2397 32539 2431
rect 33425 2397 33459 2431
rect 34161 2397 34195 2431
rect 34897 2397 34931 2431
rect 36369 2397 36403 2431
rect 37381 2397 37415 2431
rect 37933 2397 37967 2431
rect 38577 2397 38611 2431
rect 39313 2397 39347 2431
rect 40049 2397 40083 2431
rect 40785 2397 40819 2431
rect 41521 2397 41555 2431
rect 42533 2397 42567 2431
rect 43085 2397 43119 2431
rect 43729 2397 43763 2431
rect 1777 2329 1811 2363
rect 3433 2329 3467 2363
rect 3617 2329 3651 2363
rect 31125 2329 31159 2363
rect 32137 2329 32171 2363
rect 32781 2329 32815 2363
rect 35633 2329 35667 2363
rect 7941 2261 7975 2295
rect 8493 2261 8527 2295
rect 9229 2261 9263 2295
rect 17877 2261 17911 2295
rect 20085 2261 20119 2295
rect 20821 2261 20855 2295
rect 21833 2261 21867 2295
rect 23765 2261 23799 2295
rect 24501 2261 24535 2295
rect 32873 2261 32907 2295
rect 33517 2261 33551 2295
rect 34253 2261 34287 2295
rect 34989 2261 35023 2295
rect 35909 2261 35943 2295
rect 36461 2261 36495 2295
rect 37473 2261 37507 2295
rect 38025 2261 38059 2295
rect 38669 2261 38703 2295
rect 39405 2261 39439 2295
rect 40141 2261 40175 2295
rect 40877 2261 40911 2295
rect 41613 2261 41647 2295
rect 42809 2261 42843 2295
rect 43177 2261 43211 2295
rect 43821 2261 43855 2295
<< metal1 >>
rect 28074 6536 28080 6588
rect 28132 6576 28138 6588
rect 28534 6576 28540 6588
rect 28132 6548 28540 6576
rect 28132 6536 28138 6548
rect 28534 6536 28540 6548
rect 28592 6536 28598 6588
rect 5902 6468 5908 6520
rect 5960 6508 5966 6520
rect 19978 6508 19984 6520
rect 5960 6480 19984 6508
rect 5960 6468 5966 6480
rect 19978 6468 19984 6480
rect 20036 6468 20042 6520
rect 9490 6400 9496 6452
rect 9548 6440 9554 6452
rect 23566 6440 23572 6452
rect 9548 6412 23572 6440
rect 9548 6400 9554 6412
rect 23566 6400 23572 6412
rect 23624 6400 23630 6452
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 25222 6372 25228 6384
rect 7708 6344 25228 6372
rect 7708 6332 7714 6344
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 35158 6304 35164 6316
rect 4212 6276 35164 6304
rect 4212 6264 4218 6276
rect 35158 6264 35164 6276
rect 35216 6264 35222 6316
rect 1946 6196 1952 6248
rect 2004 6236 2010 6248
rect 33226 6236 33232 6248
rect 2004 6208 33232 6236
rect 2004 6196 2010 6208
rect 33226 6196 33232 6208
rect 33284 6196 33290 6248
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 35066 6168 35072 6180
rect 2740 6140 35072 6168
rect 2740 6128 2746 6140
rect 35066 6128 35072 6140
rect 35124 6128 35130 6180
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 28994 6100 29000 6112
rect 13688 6072 29000 6100
rect 13688 6060 13694 6072
rect 28994 6060 29000 6072
rect 29052 6060 29058 6112
rect 8110 5992 8116 6044
rect 8168 6032 8174 6044
rect 24118 6032 24124 6044
rect 8168 6004 24124 6032
rect 8168 5992 8174 6004
rect 24118 5992 24124 6004
rect 24176 5992 24182 6044
rect 8018 5924 8024 5976
rect 8076 5964 8082 5976
rect 25130 5964 25136 5976
rect 8076 5936 25136 5964
rect 8076 5924 8082 5936
rect 25130 5924 25136 5936
rect 25188 5924 25194 5976
rect 16390 5856 16396 5908
rect 16448 5896 16454 5908
rect 40310 5896 40316 5908
rect 16448 5868 40316 5896
rect 16448 5856 16454 5868
rect 40310 5856 40316 5868
rect 40368 5856 40374 5908
rect 15746 5788 15752 5840
rect 15804 5828 15810 5840
rect 40586 5828 40592 5840
rect 15804 5800 40592 5828
rect 15804 5788 15810 5800
rect 40586 5788 40592 5800
rect 40644 5788 40650 5840
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 38654 5760 38660 5772
rect 12676 5732 38660 5760
rect 12676 5720 12682 5732
rect 38654 5720 38660 5732
rect 38712 5720 38718 5772
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 22186 5692 22192 5704
rect 9456 5664 22192 5692
rect 9456 5652 9462 5664
rect 22186 5652 22192 5664
rect 22244 5652 22250 5704
rect 7742 5584 7748 5636
rect 7800 5624 7806 5636
rect 23842 5624 23848 5636
rect 7800 5596 23848 5624
rect 7800 5584 7806 5596
rect 23842 5584 23848 5596
rect 23900 5584 23906 5636
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 25406 5556 25412 5568
rect 14976 5528 25412 5556
rect 14976 5516 14982 5528
rect 25406 5516 25412 5528
rect 25464 5516 25470 5568
rect 1104 5466 45051 5488
rect 1104 5414 11896 5466
rect 11948 5414 11960 5466
rect 12012 5414 12024 5466
rect 12076 5414 12088 5466
rect 12140 5414 12152 5466
rect 12204 5414 22843 5466
rect 22895 5414 22907 5466
rect 22959 5414 22971 5466
rect 23023 5414 23035 5466
rect 23087 5414 23099 5466
rect 23151 5414 33790 5466
rect 33842 5414 33854 5466
rect 33906 5414 33918 5466
rect 33970 5414 33982 5466
rect 34034 5414 34046 5466
rect 34098 5414 44737 5466
rect 44789 5414 44801 5466
rect 44853 5414 44865 5466
rect 44917 5414 44929 5466
rect 44981 5414 44993 5466
rect 45045 5414 45051 5466
rect 1104 5392 45051 5414
rect 5445 5355 5503 5361
rect 5445 5321 5457 5355
rect 5491 5352 5503 5355
rect 5994 5352 6000 5364
rect 5491 5324 6000 5352
rect 5491 5321 5503 5324
rect 5445 5315 5503 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6733 5355 6791 5361
rect 6733 5321 6745 5355
rect 6779 5352 6791 5355
rect 7374 5352 7380 5364
rect 6779 5324 7380 5352
rect 6779 5321 6791 5324
rect 6733 5315 6791 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5352 7527 5355
rect 7926 5352 7932 5364
rect 7515 5324 7932 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8478 5352 8484 5364
rect 8067 5324 8484 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 9030 5352 9036 5364
rect 8619 5324 9036 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 10134 5352 10140 5364
rect 9539 5324 10140 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 11238 5352 11244 5364
rect 10643 5324 11244 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 12069 5355 12127 5361
rect 12069 5321 12081 5355
rect 12115 5352 12127 5355
rect 12526 5352 12532 5364
rect 12115 5324 12532 5352
rect 12115 5321 12127 5324
rect 12069 5315 12127 5321
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 12621 5355 12679 5361
rect 12621 5321 12633 5355
rect 12667 5352 12679 5355
rect 13170 5352 13176 5364
rect 12667 5324 13176 5352
rect 12667 5321 12679 5324
rect 12621 5315 12679 5321
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 13725 5355 13783 5361
rect 13725 5321 13737 5355
rect 13771 5352 13783 5355
rect 14274 5352 14280 5364
rect 13771 5324 14280 5352
rect 13771 5321 13783 5324
rect 13725 5315 13783 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 14645 5355 14703 5361
rect 14645 5321 14657 5355
rect 14691 5352 14703 5355
rect 15102 5352 15108 5364
rect 14691 5324 15108 5352
rect 14691 5321 14703 5324
rect 14645 5315 14703 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 15197 5355 15255 5361
rect 15197 5321 15209 5355
rect 15243 5352 15255 5355
rect 15654 5352 15660 5364
rect 15243 5324 15660 5352
rect 15243 5321 15255 5324
rect 15197 5315 15255 5321
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 16206 5352 16212 5364
rect 15795 5324 16212 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 16301 5355 16359 5361
rect 16301 5321 16313 5355
rect 16347 5352 16359 5355
rect 16758 5352 16764 5364
rect 16347 5324 16764 5352
rect 16347 5321 16359 5324
rect 16301 5315 16359 5321
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 17221 5355 17279 5361
rect 17221 5321 17233 5355
rect 17267 5352 17279 5355
rect 17586 5352 17592 5364
rect 17267 5324 17592 5352
rect 17267 5321 17279 5324
rect 17221 5315 17279 5321
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 17773 5355 17831 5361
rect 17773 5321 17785 5355
rect 17819 5352 17831 5355
rect 18138 5352 18144 5364
rect 17819 5324 18144 5352
rect 17819 5321 17831 5324
rect 17773 5315 17831 5321
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 18325 5355 18383 5361
rect 18325 5321 18337 5355
rect 18371 5352 18383 5355
rect 18690 5352 18696 5364
rect 18371 5324 18696 5352
rect 18371 5321 18383 5324
rect 18325 5315 18383 5321
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 18874 5312 18880 5364
rect 18932 5312 18938 5364
rect 18984 5324 19472 5352
rect 5537 5287 5595 5293
rect 5537 5253 5549 5287
rect 5583 5284 5595 5287
rect 7561 5287 7619 5293
rect 5583 5256 6776 5284
rect 5583 5253 5595 5256
rect 5537 5247 5595 5253
rect 6748 5228 6776 5256
rect 7561 5253 7573 5287
rect 7607 5284 7619 5287
rect 7742 5284 7748 5296
rect 7607 5256 7748 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 7742 5244 7748 5256
rect 7800 5244 7806 5296
rect 8113 5287 8171 5293
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 9398 5284 9404 5296
rect 8159 5256 9404 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 12161 5287 12219 5293
rect 10152 5256 12020 5284
rect 6086 5176 6092 5228
rect 6144 5176 6150 5228
rect 6730 5176 6736 5228
rect 6788 5176 6794 5228
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 10152 5225 10180 5256
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5185 9643 5219
rect 9585 5179 9643 5185
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6546 5148 6552 5160
rect 5859 5120 6552 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 8680 5012 8708 5179
rect 9600 5080 9628 5179
rect 10502 5176 10508 5228
rect 10560 5176 10566 5228
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 11146 5216 11152 5228
rect 10735 5188 11152 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11330 5216 11336 5228
rect 11287 5188 11336 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 11606 5176 11612 5228
rect 11664 5176 11670 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 11747 5188 11928 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 10520 5148 10548 5176
rect 9907 5120 10548 5148
rect 10965 5151 11023 5157
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 10965 5117 10977 5151
rect 11011 5148 11023 5151
rect 11624 5148 11652 5176
rect 11011 5120 11652 5148
rect 11011 5117 11023 5120
rect 10965 5111 11023 5117
rect 11900 5080 11928 5188
rect 11992 5148 12020 5256
rect 12161 5253 12173 5287
rect 12207 5284 12219 5287
rect 12713 5287 12771 5293
rect 12207 5256 12664 5284
rect 12207 5253 12219 5256
rect 12161 5247 12219 5253
rect 12636 5216 12664 5256
rect 12713 5253 12725 5287
rect 12759 5284 12771 5287
rect 13630 5284 13636 5296
rect 12759 5256 13636 5284
rect 12759 5253 12771 5256
rect 12713 5247 12771 5253
rect 13630 5244 13636 5256
rect 13688 5244 13694 5296
rect 15841 5287 15899 5293
rect 13832 5256 15240 5284
rect 13078 5216 13084 5228
rect 12636 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 13832 5225 13860 5256
rect 15212 5228 15240 5256
rect 15841 5253 15853 5287
rect 15887 5284 15899 5287
rect 16942 5284 16948 5296
rect 15887 5256 16948 5284
rect 15887 5253 15899 5256
rect 15841 5247 15899 5253
rect 16942 5244 16948 5256
rect 17000 5244 17006 5296
rect 17126 5244 17132 5296
rect 17184 5284 17190 5296
rect 18984 5284 19012 5324
rect 17184 5256 19012 5284
rect 17184 5244 17190 5256
rect 19242 5244 19248 5296
rect 19300 5284 19306 5296
rect 19337 5287 19395 5293
rect 19337 5284 19349 5287
rect 19300 5256 19349 5284
rect 19300 5244 19306 5256
rect 19337 5253 19349 5256
rect 19383 5253 19395 5287
rect 19444 5284 19472 5324
rect 19518 5312 19524 5364
rect 19576 5352 19582 5364
rect 21910 5352 21916 5364
rect 19576 5324 20484 5352
rect 19576 5312 19582 5324
rect 19444 5256 19840 5284
rect 19337 5247 19395 5253
rect 13265 5219 13323 5225
rect 13265 5216 13277 5219
rect 13228 5188 13277 5216
rect 13228 5176 13234 5188
rect 13265 5185 13277 5188
rect 13311 5185 13323 5219
rect 13265 5179 13323 5185
rect 13817 5219 13875 5225
rect 13817 5185 13829 5219
rect 13863 5185 13875 5219
rect 13817 5179 13875 5185
rect 14734 5176 14740 5228
rect 14792 5176 14798 5228
rect 15194 5176 15200 5228
rect 15252 5176 15258 5228
rect 15286 5176 15292 5228
rect 15344 5176 15350 5228
rect 16411 5219 16469 5225
rect 16411 5216 16423 5219
rect 16316 5188 16423 5216
rect 11992 5120 12434 5148
rect 12406 5080 12434 5120
rect 13262 5080 13268 5092
rect 9600 5052 11836 5080
rect 11900 5052 12112 5080
rect 12406 5052 13268 5080
rect 11238 5012 11244 5024
rect 8680 4984 11244 5012
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 11808 5012 11836 5052
rect 11882 5012 11888 5024
rect 11808 4984 11888 5012
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12084 5012 12112 5052
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 16316 5080 16344 5188
rect 16411 5185 16423 5188
rect 16457 5185 16469 5219
rect 16411 5179 16469 5185
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5216 17371 5219
rect 17770 5216 17776 5228
rect 17359 5188 17776 5216
rect 17359 5185 17371 5188
rect 17313 5179 17371 5185
rect 17770 5176 17776 5188
rect 17828 5176 17834 5228
rect 17865 5219 17923 5225
rect 17865 5185 17877 5219
rect 17911 5216 17923 5219
rect 17954 5216 17960 5228
rect 17911 5188 17960 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5216 18475 5219
rect 18874 5216 18880 5228
rect 18463 5188 18880 5216
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 18966 5176 18972 5228
rect 19024 5176 19030 5228
rect 19702 5176 19708 5228
rect 19760 5176 19766 5228
rect 19812 5216 19840 5256
rect 19886 5244 19892 5296
rect 19944 5244 19950 5296
rect 20456 5293 20484 5324
rect 20732 5324 21916 5352
rect 20441 5287 20499 5293
rect 20441 5253 20453 5287
rect 20487 5253 20499 5287
rect 20441 5247 20499 5253
rect 20162 5216 20168 5228
rect 19812 5188 20168 5216
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20732 5216 20760 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 24762 5312 24768 5364
rect 24820 5352 24826 5364
rect 27525 5355 27583 5361
rect 27525 5352 27537 5355
rect 24820 5324 25176 5352
rect 24820 5312 24826 5324
rect 20809 5287 20867 5293
rect 20809 5253 20821 5287
rect 20855 5284 20867 5287
rect 24946 5284 24952 5296
rect 20855 5256 24952 5284
rect 20855 5253 20867 5256
rect 20809 5247 20867 5253
rect 24946 5244 24952 5256
rect 25004 5244 25010 5296
rect 25148 5249 25176 5324
rect 26896 5324 27537 5352
rect 25133 5243 25191 5249
rect 25314 5244 25320 5296
rect 25372 5284 25378 5296
rect 25372 5256 25728 5284
rect 25372 5244 25378 5256
rect 20303 5188 20760 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 21358 5176 21364 5228
rect 21416 5176 21422 5228
rect 21634 5176 21640 5228
rect 21692 5176 21698 5228
rect 21726 5176 21732 5228
rect 21784 5216 21790 5228
rect 22005 5219 22063 5225
rect 22005 5216 22017 5219
rect 21784 5188 22017 5216
rect 21784 5176 21790 5188
rect 22005 5185 22017 5188
rect 22051 5185 22063 5219
rect 22005 5179 22063 5185
rect 22094 5176 22100 5228
rect 22152 5216 22158 5228
rect 22281 5219 22339 5225
rect 22281 5216 22293 5219
rect 22152 5188 22293 5216
rect 22152 5176 22158 5188
rect 22281 5185 22293 5188
rect 22327 5185 22339 5219
rect 22281 5179 22339 5185
rect 22554 5176 22560 5228
rect 22612 5176 22618 5228
rect 22830 5176 22836 5228
rect 22888 5176 22894 5228
rect 23106 5176 23112 5228
rect 23164 5176 23170 5228
rect 23382 5176 23388 5228
rect 23440 5176 23446 5228
rect 23474 5176 23480 5228
rect 23532 5216 23538 5228
rect 23661 5219 23719 5225
rect 23661 5216 23673 5219
rect 23532 5188 23673 5216
rect 23532 5176 23538 5188
rect 23661 5185 23673 5188
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23937 5219 23995 5225
rect 23937 5216 23949 5219
rect 23808 5188 23949 5216
rect 23808 5176 23814 5188
rect 23937 5185 23949 5188
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 24026 5176 24032 5228
rect 24084 5216 24090 5228
rect 24213 5219 24271 5225
rect 24213 5216 24225 5219
rect 24084 5188 24225 5216
rect 24084 5176 24090 5188
rect 24213 5185 24225 5188
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 24302 5176 24308 5228
rect 24360 5216 24366 5228
rect 24581 5219 24639 5225
rect 24581 5216 24593 5219
rect 24360 5188 24593 5216
rect 24360 5176 24366 5188
rect 24581 5185 24593 5188
rect 24627 5185 24639 5219
rect 24581 5179 24639 5185
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 25133 5209 25145 5243
rect 25179 5209 25191 5243
rect 25700 5225 25728 5256
rect 25866 5244 25872 5296
rect 25924 5284 25930 5296
rect 26896 5284 26924 5324
rect 27525 5321 27537 5324
rect 27571 5321 27583 5355
rect 27525 5315 27583 5321
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 32861 5355 32919 5361
rect 27672 5324 28028 5352
rect 27672 5312 27678 5324
rect 25924 5256 26924 5284
rect 25924 5244 25930 5256
rect 26970 5244 26976 5296
rect 27028 5284 27034 5296
rect 27028 5256 27476 5284
rect 27028 5244 27034 5256
rect 25133 5203 25191 5209
rect 25409 5219 25467 5225
rect 25409 5185 25421 5219
rect 25455 5185 25467 5219
rect 25409 5179 25467 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5185 25743 5219
rect 25685 5179 25743 5185
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 23014 5148 23020 5160
rect 18380 5120 23020 5148
rect 18380 5108 18386 5120
rect 23014 5108 23020 5120
rect 23072 5108 23078 5160
rect 25038 5108 25044 5160
rect 25096 5148 25102 5160
rect 25424 5148 25452 5179
rect 25774 5176 25780 5228
rect 25832 5176 25838 5228
rect 26050 5176 26056 5228
rect 26108 5176 26114 5228
rect 26326 5176 26332 5228
rect 26384 5176 26390 5228
rect 26602 5176 26608 5228
rect 26660 5176 26666 5228
rect 26694 5176 26700 5228
rect 26752 5216 26758 5228
rect 27448 5225 27476 5256
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26752 5188 27169 5216
rect 26752 5176 26758 5188
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27433 5219 27491 5225
rect 27433 5185 27445 5219
rect 27479 5185 27491 5219
rect 27433 5179 27491 5185
rect 27706 5176 27712 5228
rect 27764 5176 27770 5228
rect 28000 5225 28028 5324
rect 32861 5321 32873 5355
rect 32907 5352 32919 5355
rect 34514 5352 34520 5364
rect 32907 5324 34520 5352
rect 32907 5321 32919 5324
rect 32861 5315 32919 5321
rect 34514 5312 34520 5324
rect 34572 5312 34578 5364
rect 34606 5312 34612 5364
rect 34664 5352 34670 5364
rect 34885 5355 34943 5361
rect 34885 5352 34897 5355
rect 34664 5324 34897 5352
rect 34664 5312 34670 5324
rect 34885 5321 34897 5324
rect 34931 5321 34943 5355
rect 34885 5315 34943 5321
rect 34974 5312 34980 5364
rect 35032 5352 35038 5364
rect 35437 5355 35495 5361
rect 35437 5352 35449 5355
rect 35032 5324 35449 5352
rect 35032 5312 35038 5324
rect 35437 5321 35449 5324
rect 35483 5321 35495 5355
rect 35437 5315 35495 5321
rect 35526 5312 35532 5364
rect 35584 5352 35590 5364
rect 35989 5355 36047 5361
rect 35989 5352 36001 5355
rect 35584 5324 36001 5352
rect 35584 5312 35590 5324
rect 35989 5321 36001 5324
rect 36035 5321 36047 5355
rect 35989 5315 36047 5321
rect 36538 5312 36544 5364
rect 36596 5352 36602 5364
rect 37461 5355 37519 5361
rect 37461 5352 37473 5355
rect 36596 5324 37473 5352
rect 36596 5312 36602 5324
rect 37461 5321 37473 5324
rect 37507 5321 37519 5355
rect 37461 5315 37519 5321
rect 38194 5312 38200 5364
rect 38252 5352 38258 5364
rect 39117 5355 39175 5361
rect 39117 5352 39129 5355
rect 38252 5324 39129 5352
rect 38252 5312 38258 5324
rect 39117 5321 39129 5324
rect 39163 5321 39175 5355
rect 39117 5315 39175 5321
rect 39666 5312 39672 5364
rect 39724 5352 39730 5364
rect 40589 5355 40647 5361
rect 40589 5352 40601 5355
rect 39724 5324 40601 5352
rect 39724 5312 39730 5324
rect 40589 5321 40601 5324
rect 40635 5321 40647 5355
rect 40589 5315 40647 5321
rect 41141 5355 41199 5361
rect 41141 5321 41153 5355
rect 41187 5321 41199 5355
rect 41141 5315 41199 5321
rect 28350 5244 28356 5296
rect 28408 5284 28414 5296
rect 28408 5256 28672 5284
rect 28408 5244 28414 5256
rect 27985 5219 28043 5225
rect 27985 5185 27997 5219
rect 28031 5185 28043 5219
rect 27985 5179 28043 5185
rect 28261 5219 28319 5225
rect 28261 5185 28273 5219
rect 28307 5185 28319 5219
rect 28261 5179 28319 5185
rect 25096 5120 25452 5148
rect 25096 5108 25102 5120
rect 27798 5108 27804 5160
rect 27856 5148 27862 5160
rect 28276 5148 28304 5179
rect 28534 5176 28540 5228
rect 28592 5176 28598 5228
rect 28644 5216 28672 5256
rect 28718 5244 28724 5296
rect 28776 5284 28782 5296
rect 28776 5256 29132 5284
rect 28776 5244 28782 5256
rect 29104 5225 29132 5256
rect 36648 5256 38516 5284
rect 28813 5219 28871 5225
rect 28813 5216 28825 5219
rect 28644 5188 28825 5216
rect 28813 5185 28825 5188
rect 28859 5185 28871 5219
rect 28813 5179 28871 5185
rect 29089 5219 29147 5225
rect 29089 5185 29101 5219
rect 29135 5185 29147 5219
rect 29089 5179 29147 5185
rect 30098 5176 30104 5228
rect 30156 5176 30162 5228
rect 30374 5176 30380 5228
rect 30432 5176 30438 5228
rect 30650 5176 30656 5228
rect 30708 5176 30714 5228
rect 30926 5176 30932 5228
rect 30984 5176 30990 5228
rect 31202 5176 31208 5228
rect 31260 5176 31266 5228
rect 31478 5176 31484 5228
rect 31536 5176 31542 5228
rect 31754 5176 31760 5228
rect 31812 5176 31818 5228
rect 32122 5176 32128 5228
rect 32180 5176 32186 5228
rect 32398 5176 32404 5228
rect 32456 5176 32462 5228
rect 32674 5176 32680 5228
rect 32732 5176 32738 5228
rect 32950 5176 32956 5228
rect 33008 5176 33014 5228
rect 33042 5176 33048 5228
rect 33100 5216 33106 5228
rect 33229 5219 33287 5225
rect 33229 5216 33241 5219
rect 33100 5188 33241 5216
rect 33100 5176 33106 5188
rect 33229 5185 33241 5188
rect 33275 5185 33287 5219
rect 33229 5179 33287 5185
rect 33502 5176 33508 5228
rect 33560 5176 33566 5228
rect 33778 5176 33784 5228
rect 33836 5176 33842 5228
rect 34238 5176 34244 5228
rect 34296 5176 34302 5228
rect 34330 5176 34336 5228
rect 34388 5216 34394 5228
rect 34517 5219 34575 5225
rect 34517 5216 34529 5219
rect 34388 5188 34529 5216
rect 34388 5176 34394 5188
rect 34517 5185 34529 5188
rect 34563 5185 34575 5219
rect 34517 5179 34575 5185
rect 34606 5176 34612 5228
rect 34664 5216 34670 5228
rect 34793 5219 34851 5225
rect 34793 5216 34805 5219
rect 34664 5188 34805 5216
rect 34664 5176 34670 5188
rect 34793 5185 34805 5188
rect 34839 5185 34851 5219
rect 34793 5179 34851 5185
rect 35342 5176 35348 5228
rect 35400 5176 35406 5228
rect 35897 5219 35955 5225
rect 35897 5216 35909 5219
rect 35452 5188 35909 5216
rect 27856 5120 28304 5148
rect 32508 5120 34376 5148
rect 27856 5108 27862 5120
rect 32508 5092 32536 5120
rect 22002 5080 22008 5092
rect 16316 5052 22008 5080
rect 22002 5040 22008 5052
rect 22060 5040 22066 5092
rect 27982 5080 27988 5092
rect 22204 5052 27988 5080
rect 22204 5024 22232 5052
rect 27982 5040 27988 5052
rect 28040 5040 28046 5092
rect 31389 5083 31447 5089
rect 31389 5049 31401 5083
rect 31435 5080 31447 5083
rect 31846 5080 31852 5092
rect 31435 5052 31852 5080
rect 31435 5049 31447 5052
rect 31389 5043 31447 5049
rect 31846 5040 31852 5052
rect 31904 5040 31910 5092
rect 32490 5040 32496 5092
rect 32548 5040 32554 5092
rect 32585 5083 32643 5089
rect 32585 5049 32597 5083
rect 32631 5080 32643 5083
rect 33042 5080 33048 5092
rect 32631 5052 33048 5080
rect 32631 5049 32643 5052
rect 32585 5043 32643 5049
rect 33042 5040 33048 5052
rect 33100 5040 33106 5092
rect 33134 5040 33140 5092
rect 33192 5040 33198 5092
rect 33318 5040 33324 5092
rect 33376 5080 33382 5092
rect 34348 5089 34376 5120
rect 35250 5108 35256 5160
rect 35308 5148 35314 5160
rect 35452 5148 35480 5188
rect 35897 5185 35909 5188
rect 35943 5185 35955 5219
rect 35897 5179 35955 5185
rect 36449 5219 36507 5225
rect 36449 5185 36461 5219
rect 36495 5185 36507 5219
rect 36449 5179 36507 5185
rect 35308 5120 35480 5148
rect 35308 5108 35314 5120
rect 35526 5108 35532 5160
rect 35584 5148 35590 5160
rect 36464 5148 36492 5179
rect 35584 5120 36492 5148
rect 35584 5108 35590 5120
rect 34057 5083 34115 5089
rect 34057 5080 34069 5083
rect 33376 5052 34069 5080
rect 33376 5040 33382 5052
rect 34057 5049 34069 5052
rect 34103 5049 34115 5083
rect 34057 5043 34115 5049
rect 34333 5083 34391 5089
rect 34333 5049 34345 5083
rect 34379 5049 34391 5083
rect 34333 5043 34391 5049
rect 34422 5040 34428 5092
rect 34480 5080 34486 5092
rect 36648 5080 36676 5256
rect 36722 5176 36728 5228
rect 36780 5216 36786 5228
rect 38488 5225 38516 5256
rect 38654 5244 38660 5296
rect 38712 5284 38718 5296
rect 39945 5287 40003 5293
rect 39945 5284 39957 5287
rect 38712 5256 39957 5284
rect 38712 5244 38718 5256
rect 39945 5253 39957 5256
rect 39991 5253 40003 5287
rect 39945 5247 40003 5253
rect 40034 5244 40040 5296
rect 40092 5284 40098 5296
rect 41156 5284 41184 5315
rect 40092 5256 41184 5284
rect 40092 5244 40098 5256
rect 37369 5219 37427 5225
rect 37369 5216 37381 5219
rect 36780 5188 37381 5216
rect 36780 5176 36786 5188
rect 37369 5185 37381 5188
rect 37415 5185 37427 5219
rect 37369 5179 37427 5185
rect 37921 5219 37979 5225
rect 37921 5185 37933 5219
rect 37967 5185 37979 5219
rect 37921 5179 37979 5185
rect 38473 5219 38531 5225
rect 38473 5185 38485 5219
rect 38519 5185 38531 5219
rect 38473 5179 38531 5185
rect 39025 5219 39083 5225
rect 39025 5185 39037 5219
rect 39071 5185 39083 5219
rect 39025 5179 39083 5185
rect 37182 5108 37188 5160
rect 37240 5148 37246 5160
rect 37936 5148 37964 5179
rect 37240 5120 37964 5148
rect 37240 5108 37246 5120
rect 38010 5108 38016 5160
rect 38068 5148 38074 5160
rect 39040 5148 39068 5179
rect 40494 5176 40500 5228
rect 40552 5176 40558 5228
rect 40586 5176 40592 5228
rect 40644 5216 40650 5228
rect 41049 5219 41107 5225
rect 41049 5216 41061 5219
rect 40644 5188 41061 5216
rect 40644 5176 40650 5188
rect 41049 5185 41061 5188
rect 41095 5185 41107 5219
rect 41049 5179 41107 5185
rect 38068 5120 39068 5148
rect 38068 5108 38074 5120
rect 34480 5052 36676 5080
rect 34480 5040 34486 5052
rect 37642 5040 37648 5092
rect 37700 5080 37706 5092
rect 38657 5083 38715 5089
rect 38657 5080 38669 5083
rect 37700 5052 38669 5080
rect 37700 5040 37706 5052
rect 38657 5049 38669 5052
rect 38703 5049 38715 5083
rect 38657 5043 38715 5049
rect 12802 5012 12808 5024
rect 12084 4984 12808 5012
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 13173 5015 13231 5021
rect 13173 4981 13185 5015
rect 13219 5012 13231 5015
rect 13722 5012 13728 5024
rect 13219 4984 13728 5012
rect 13219 4981 13231 4984
rect 13173 4975 13231 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 20530 5012 20536 5024
rect 13872 4984 20536 5012
rect 13872 4972 13878 4984
rect 20530 4972 20536 4984
rect 20588 4972 20594 5024
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 21177 5015 21235 5021
rect 21177 5012 21189 5015
rect 20772 4984 21189 5012
rect 20772 4972 20778 4984
rect 21177 4981 21189 4984
rect 21223 4981 21235 5015
rect 21177 4975 21235 4981
rect 21266 4972 21272 5024
rect 21324 5012 21330 5024
rect 21453 5015 21511 5021
rect 21453 5012 21465 5015
rect 21324 4984 21465 5012
rect 21324 4972 21330 4984
rect 21453 4981 21465 4984
rect 21499 4981 21511 5015
rect 21453 4975 21511 4981
rect 21818 4972 21824 5024
rect 21876 4972 21882 5024
rect 22094 4972 22100 5024
rect 22152 4972 22158 5024
rect 22186 4972 22192 5024
rect 22244 4972 22250 5024
rect 22370 4972 22376 5024
rect 22428 4972 22434 5024
rect 22646 4972 22652 5024
rect 22704 4972 22710 5024
rect 22922 4972 22928 5024
rect 22980 4972 22986 5024
rect 23198 4972 23204 5024
rect 23256 4972 23262 5024
rect 23474 4972 23480 5024
rect 23532 4972 23538 5024
rect 23750 4972 23756 5024
rect 23808 4972 23814 5024
rect 24026 4972 24032 5024
rect 24084 4972 24090 5024
rect 24394 4972 24400 5024
rect 24452 4972 24458 5024
rect 24670 4972 24676 5024
rect 24728 4972 24734 5024
rect 24946 4972 24952 5024
rect 25004 4972 25010 5024
rect 25222 4972 25228 5024
rect 25280 4972 25286 5024
rect 25498 4972 25504 5024
rect 25556 4972 25562 5024
rect 25958 4972 25964 5024
rect 26016 4972 26022 5024
rect 26234 4972 26240 5024
rect 26292 4972 26298 5024
rect 26510 4972 26516 5024
rect 26568 4972 26574 5024
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 26789 5015 26847 5021
rect 26789 5012 26801 5015
rect 26752 4984 26801 5012
rect 26752 4972 26758 4984
rect 26789 4981 26801 4984
rect 26835 4981 26847 5015
rect 26789 4975 26847 4981
rect 26970 4972 26976 5024
rect 27028 4972 27034 5024
rect 27246 4972 27252 5024
rect 27304 4972 27310 5024
rect 27798 4972 27804 5024
rect 27856 4972 27862 5024
rect 27890 4972 27896 5024
rect 27948 5012 27954 5024
rect 28077 5015 28135 5021
rect 28077 5012 28089 5015
rect 27948 4984 28089 5012
rect 27948 4972 27954 4984
rect 28077 4981 28089 4984
rect 28123 4981 28135 5015
rect 28077 4975 28135 4981
rect 28258 4972 28264 5024
rect 28316 5012 28322 5024
rect 28353 5015 28411 5021
rect 28353 5012 28365 5015
rect 28316 4984 28365 5012
rect 28316 4972 28322 4984
rect 28353 4981 28365 4984
rect 28399 4981 28411 5015
rect 28353 4975 28411 4981
rect 28629 5015 28687 5021
rect 28629 4981 28641 5015
rect 28675 5012 28687 5015
rect 28718 5012 28724 5024
rect 28675 4984 28724 5012
rect 28675 4981 28687 4984
rect 28629 4975 28687 4981
rect 28718 4972 28724 4984
rect 28776 4972 28782 5024
rect 28902 4972 28908 5024
rect 28960 4972 28966 5024
rect 30285 5015 30343 5021
rect 30285 4981 30297 5015
rect 30331 5012 30343 5015
rect 30466 5012 30472 5024
rect 30331 4984 30472 5012
rect 30331 4981 30343 4984
rect 30285 4975 30343 4981
rect 30466 4972 30472 4984
rect 30524 4972 30530 5024
rect 30558 4972 30564 5024
rect 30616 4972 30622 5024
rect 30834 4972 30840 5024
rect 30892 4972 30898 5024
rect 31110 4972 31116 5024
rect 31168 4972 31174 5024
rect 31665 5015 31723 5021
rect 31665 4981 31677 5015
rect 31711 5012 31723 5015
rect 31754 5012 31760 5024
rect 31711 4984 31760 5012
rect 31711 4981 31723 4984
rect 31665 4975 31723 4981
rect 31754 4972 31760 4984
rect 31812 4972 31818 5024
rect 31938 4972 31944 5024
rect 31996 4972 32002 5024
rect 32306 4972 32312 5024
rect 32364 4972 32370 5024
rect 33410 4972 33416 5024
rect 33468 4972 33474 5024
rect 33686 4972 33692 5024
rect 33744 4972 33750 5024
rect 33965 5015 34023 5021
rect 33965 4981 33977 5015
rect 34011 5012 34023 5015
rect 34146 5012 34152 5024
rect 34011 4984 34152 5012
rect 34011 4981 34023 4984
rect 33965 4975 34023 4981
rect 34146 4972 34152 4984
rect 34204 4972 34210 5024
rect 35710 4972 35716 5024
rect 35768 5012 35774 5024
rect 36541 5015 36599 5021
rect 36541 5012 36553 5015
rect 35768 4984 36553 5012
rect 35768 4972 35774 4984
rect 36541 4981 36553 4984
rect 36587 4981 36599 5015
rect 36541 4975 36599 4981
rect 36906 4972 36912 5024
rect 36964 5012 36970 5024
rect 38013 5015 38071 5021
rect 38013 5012 38025 5015
rect 36964 4984 38025 5012
rect 36964 4972 36970 4984
rect 38013 4981 38025 4984
rect 38059 4981 38071 5015
rect 38013 4975 38071 4981
rect 39298 4972 39304 5024
rect 39356 5012 39362 5024
rect 40037 5015 40095 5021
rect 40037 5012 40049 5015
rect 39356 4984 40049 5012
rect 39356 4972 39362 4984
rect 40037 4981 40049 4984
rect 40083 4981 40095 5015
rect 40037 4975 40095 4981
rect 1104 4922 44896 4944
rect 1104 4870 6423 4922
rect 6475 4870 6487 4922
rect 6539 4870 6551 4922
rect 6603 4870 6615 4922
rect 6667 4870 6679 4922
rect 6731 4870 17370 4922
rect 17422 4870 17434 4922
rect 17486 4870 17498 4922
rect 17550 4870 17562 4922
rect 17614 4870 17626 4922
rect 17678 4870 28317 4922
rect 28369 4870 28381 4922
rect 28433 4870 28445 4922
rect 28497 4870 28509 4922
rect 28561 4870 28573 4922
rect 28625 4870 39264 4922
rect 39316 4870 39328 4922
rect 39380 4870 39392 4922
rect 39444 4870 39456 4922
rect 39508 4870 39520 4922
rect 39572 4870 44896 4922
rect 1104 4848 44896 4870
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 6144 4780 7236 4808
rect 6144 4768 6150 4780
rect 5718 4700 5724 4752
rect 5776 4700 5782 4752
rect 6270 4700 6276 4752
rect 6328 4700 6334 4752
rect 6822 4700 6828 4752
rect 6880 4700 6886 4752
rect 7208 4740 7236 4780
rect 7282 4768 7288 4820
rect 7340 4768 7346 4820
rect 7834 4768 7840 4820
rect 7892 4768 7898 4820
rect 8386 4768 8392 4820
rect 8444 4768 8450 4820
rect 9306 4768 9312 4820
rect 9364 4768 9370 4820
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 10410 4768 10416 4820
rect 10468 4768 10474 4820
rect 11054 4768 11060 4820
rect 11112 4768 11118 4820
rect 11422 4768 11428 4820
rect 11480 4768 11486 4820
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 12434 4768 12440 4820
rect 12492 4768 12498 4820
rect 12986 4768 12992 4820
rect 13044 4768 13050 4820
rect 13538 4768 13544 4820
rect 13596 4768 13602 4820
rect 14182 4768 14188 4820
rect 14240 4768 14246 4820
rect 14292 4780 15516 4808
rect 11698 4740 11704 4752
rect 7208 4712 11704 4740
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 14292 4740 14320 4780
rect 13740 4712 14320 4740
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6236 4576 6469 4604
rect 6236 4564 6242 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 7009 4607 7067 4613
rect 7009 4573 7021 4607
rect 7055 4604 7067 4607
rect 8018 4604 8024 4616
rect 7055 4576 8024 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8110 4564 8116 4616
rect 8168 4564 8174 4616
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9490 4604 9496 4616
rect 8711 4576 9496 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 9490 4564 9496 4576
rect 9548 4564 9554 4616
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4604 10011 4607
rect 11333 4607 11391 4613
rect 9999 4576 11284 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 7561 4539 7619 4545
rect 7561 4505 7573 4539
rect 7607 4536 7619 4539
rect 7650 4536 7656 4548
rect 7607 4508 7656 4536
rect 7607 4505 7619 4508
rect 7561 4499 7619 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 9398 4496 9404 4548
rect 9456 4496 9462 4548
rect 10505 4539 10563 4545
rect 10505 4505 10517 4539
rect 10551 4505 10563 4539
rect 10505 4499 10563 4505
rect 10520 4468 10548 4499
rect 10778 4496 10784 4548
rect 10836 4496 10842 4548
rect 11256 4536 11284 4576
rect 11333 4573 11345 4607
rect 11379 4604 11391 4607
rect 11422 4604 11428 4616
rect 11379 4576 11428 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 13740 4604 13768 4712
rect 14826 4700 14832 4752
rect 14884 4700 14890 4752
rect 15378 4700 15384 4752
rect 15436 4700 15442 4752
rect 15488 4740 15516 4780
rect 15930 4768 15936 4820
rect 15988 4768 15994 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16080 4780 17172 4808
rect 16080 4768 16086 4780
rect 15488 4712 15976 4740
rect 15102 4672 15108 4684
rect 13832 4644 15108 4672
rect 13832 4613 13860 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 15948 4672 15976 4712
rect 16482 4700 16488 4752
rect 16540 4700 16546 4752
rect 17034 4700 17040 4752
rect 17092 4700 17098 4752
rect 17144 4740 17172 4780
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 17497 4811 17555 4817
rect 17497 4808 17509 4811
rect 17368 4780 17509 4808
rect 17368 4768 17374 4780
rect 17497 4777 17509 4780
rect 17543 4777 17555 4811
rect 17497 4771 17555 4777
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 17920 4780 18153 4808
rect 17920 4768 17926 4780
rect 18141 4777 18153 4780
rect 18187 4777 18199 4811
rect 18141 4771 18199 4777
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18693 4811 18751 4817
rect 18693 4808 18705 4811
rect 18472 4780 18705 4808
rect 18472 4768 18478 4780
rect 18693 4777 18705 4780
rect 18739 4777 18751 4811
rect 18693 4771 18751 4777
rect 18782 4768 18788 4820
rect 18840 4808 18846 4820
rect 19794 4808 19800 4820
rect 18840 4780 19800 4808
rect 18840 4768 18846 4780
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 19996 4780 20208 4808
rect 17144 4712 18276 4740
rect 17126 4672 17132 4684
rect 15712 4644 15884 4672
rect 15948 4644 17132 4672
rect 15712 4632 15718 4644
rect 12084 4576 13768 4604
rect 13817 4607 13875 4613
rect 12084 4536 12112 4576
rect 13817 4573 13829 4607
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 14918 4604 14924 4616
rect 14507 4576 14924 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4604 15071 4607
rect 15378 4604 15384 4616
rect 15059 4576 15384 4604
rect 15059 4573 15071 4576
rect 15013 4567 15071 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15562 4564 15568 4616
rect 15620 4564 15626 4616
rect 15856 4613 15884 4644
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 18248 4672 18276 4712
rect 19334 4700 19340 4752
rect 19392 4700 19398 4752
rect 19886 4740 19892 4752
rect 19444 4712 19892 4740
rect 19444 4672 19472 4712
rect 19886 4700 19892 4712
rect 19944 4700 19950 4752
rect 19996 4672 20024 4780
rect 20180 4749 20208 4780
rect 20438 4768 20444 4820
rect 20496 4808 20502 4820
rect 20717 4811 20775 4817
rect 20717 4808 20729 4811
rect 20496 4780 20729 4808
rect 20496 4768 20502 4780
rect 20717 4777 20729 4780
rect 20763 4777 20775 4811
rect 21729 4811 21787 4817
rect 21729 4808 21741 4811
rect 20717 4771 20775 4777
rect 20824 4780 21741 4808
rect 20165 4743 20223 4749
rect 20165 4709 20177 4743
rect 20211 4709 20223 4743
rect 20165 4703 20223 4709
rect 17788 4644 18184 4672
rect 18248 4644 19472 4672
rect 19536 4644 20024 4672
rect 17788 4613 17816 4644
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 17773 4607 17831 4613
rect 15841 4567 15899 4573
rect 16592 4576 17724 4604
rect 11256 4508 12112 4536
rect 12161 4539 12219 4545
rect 12161 4505 12173 4539
rect 12207 4536 12219 4539
rect 12250 4536 12256 4548
rect 12207 4508 12256 4536
rect 12207 4505 12219 4508
rect 12161 4499 12219 4505
rect 12250 4496 12256 4508
rect 12308 4496 12314 4548
rect 12710 4496 12716 4548
rect 12768 4496 12774 4548
rect 13262 4496 13268 4548
rect 13320 4496 13326 4548
rect 13354 4496 13360 4548
rect 13412 4536 13418 4548
rect 16592 4536 16620 4576
rect 13412 4508 16620 4536
rect 13412 4496 13418 4508
rect 16666 4496 16672 4548
rect 16724 4496 16730 4548
rect 17218 4496 17224 4548
rect 17276 4496 17282 4548
rect 17696 4536 17724 4576
rect 17773 4573 17785 4607
rect 17819 4573 17831 4607
rect 17773 4567 17831 4573
rect 18046 4564 18052 4616
rect 18104 4564 18110 4616
rect 18156 4604 18184 4644
rect 18322 4604 18328 4616
rect 18156 4576 18328 4604
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 19536 4613 19564 4644
rect 20254 4632 20260 4684
rect 20312 4672 20318 4684
rect 20824 4672 20852 4780
rect 21729 4777 21741 4780
rect 21775 4777 21787 4811
rect 22094 4808 22100 4820
rect 21729 4771 21787 4777
rect 22066 4768 22100 4808
rect 22152 4768 22158 4820
rect 22646 4768 22652 4820
rect 22704 4768 22710 4820
rect 22922 4808 22928 4820
rect 22756 4780 22928 4808
rect 21361 4743 21419 4749
rect 21361 4709 21373 4743
rect 21407 4740 21419 4743
rect 21450 4740 21456 4752
rect 21407 4712 21456 4740
rect 21407 4709 21419 4712
rect 21361 4703 21419 4709
rect 21450 4700 21456 4712
rect 21508 4700 21514 4752
rect 22066 4740 22094 4768
rect 21560 4712 22094 4740
rect 20312 4644 20852 4672
rect 20312 4632 20318 4644
rect 19521 4607 19579 4613
rect 18524 4576 19472 4604
rect 18524 4536 18552 4576
rect 17696 4508 18552 4536
rect 18598 4496 18604 4548
rect 18656 4496 18662 4548
rect 18782 4496 18788 4548
rect 18840 4496 18846 4548
rect 18800 4468 18828 4496
rect 10520 4440 18828 4468
rect 19444 4468 19472 4576
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 20070 4613 20076 4616
rect 19797 4607 19855 4613
rect 19668 4576 19748 4604
rect 19668 4564 19674 4576
rect 19518 4468 19524 4480
rect 19444 4440 19524 4468
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19613 4471 19671 4477
rect 19613 4437 19625 4471
rect 19659 4468 19671 4471
rect 19720 4468 19748 4576
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 19843 4576 20024 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 19659 4440 19748 4468
rect 19659 4437 19671 4440
rect 19613 4431 19671 4437
rect 19886 4428 19892 4480
rect 19944 4428 19950 4480
rect 19996 4468 20024 4576
rect 20065 4567 20076 4613
rect 20070 4564 20076 4567
rect 20128 4564 20134 4616
rect 20346 4564 20352 4616
rect 20404 4564 20410 4616
rect 20530 4564 20536 4616
rect 20588 4564 20594 4616
rect 20622 4564 20628 4616
rect 20680 4564 20686 4616
rect 20901 4607 20959 4613
rect 20901 4573 20913 4607
rect 20947 4604 20959 4607
rect 21177 4607 21235 4613
rect 20947 4576 21128 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 20548 4536 20576 4564
rect 20806 4536 20812 4548
rect 20548 4508 20812 4536
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 21100 4536 21128 4576
rect 21177 4573 21189 4607
rect 21223 4604 21235 4607
rect 21358 4604 21364 4616
rect 21223 4576 21364 4604
rect 21223 4573 21235 4576
rect 21177 4567 21235 4573
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 21560 4613 21588 4712
rect 21818 4632 21824 4684
rect 21876 4632 21882 4684
rect 22664 4672 22692 4768
rect 22204 4644 22692 4672
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 21836 4536 21864 4632
rect 22204 4613 22232 4644
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4604 21971 4607
rect 22189 4607 22247 4613
rect 21959 4576 22094 4604
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 21100 4508 21864 4536
rect 22066 4536 22094 4576
rect 22189 4573 22201 4607
rect 22235 4573 22247 4607
rect 22189 4567 22247 4573
rect 22370 4564 22376 4616
rect 22428 4564 22434 4616
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4604 22523 4607
rect 22756 4604 22784 4780
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 23198 4768 23204 4820
rect 23256 4768 23262 4820
rect 23474 4808 23480 4820
rect 23308 4780 23480 4808
rect 23216 4672 23244 4768
rect 22848 4644 23244 4672
rect 22848 4613 22876 4644
rect 22511 4576 22784 4604
rect 22833 4607 22891 4613
rect 22511 4573 22523 4576
rect 22465 4567 22523 4573
rect 22833 4573 22845 4607
rect 22879 4573 22891 4607
rect 22833 4567 22891 4573
rect 23109 4607 23167 4613
rect 23109 4573 23121 4607
rect 23155 4604 23167 4607
rect 23308 4604 23336 4780
rect 23474 4768 23480 4780
rect 23532 4768 23538 4820
rect 23750 4768 23756 4820
rect 23808 4768 23814 4820
rect 24026 4808 24032 4820
rect 23860 4780 24032 4808
rect 23768 4672 23796 4768
rect 23400 4644 23796 4672
rect 23400 4613 23428 4644
rect 23155 4576 23336 4604
rect 23385 4607 23443 4613
rect 23155 4573 23167 4576
rect 23109 4567 23167 4573
rect 23385 4573 23397 4607
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 23566 4564 23572 4616
rect 23624 4564 23630 4616
rect 23661 4607 23719 4613
rect 23661 4573 23673 4607
rect 23707 4604 23719 4607
rect 23860 4604 23888 4780
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 24394 4768 24400 4820
rect 24452 4768 24458 4820
rect 24670 4768 24676 4820
rect 24728 4768 24734 4820
rect 24854 4768 24860 4820
rect 24912 4808 24918 4820
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 24912 4780 25789 4808
rect 24912 4768 24918 4780
rect 25777 4777 25789 4780
rect 25823 4777 25835 4811
rect 25777 4771 25835 4777
rect 25958 4768 25964 4820
rect 26016 4768 26022 4820
rect 27614 4768 27620 4820
rect 27672 4768 27678 4820
rect 28166 4808 28172 4820
rect 27816 4780 28172 4808
rect 23707 4576 23888 4604
rect 24029 4607 24087 4613
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 24029 4573 24041 4607
rect 24075 4604 24087 4607
rect 24412 4604 24440 4768
rect 24075 4576 24440 4604
rect 24075 4573 24087 4576
rect 24029 4567 24087 4573
rect 24486 4564 24492 4616
rect 24544 4564 24550 4616
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 24688 4604 24716 4768
rect 24946 4700 24952 4752
rect 25004 4700 25010 4752
rect 25222 4700 25228 4752
rect 25280 4700 25286 4752
rect 25498 4700 25504 4752
rect 25556 4700 25562 4752
rect 24627 4576 24716 4604
rect 24857 4607 24915 4613
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 24857 4573 24869 4607
rect 24903 4604 24915 4607
rect 24964 4604 24992 4700
rect 24903 4576 24992 4604
rect 25133 4607 25191 4613
rect 24903 4573 24915 4576
rect 24857 4567 24915 4573
rect 25133 4573 25145 4607
rect 25179 4604 25191 4607
rect 25240 4604 25268 4700
rect 25179 4576 25268 4604
rect 25409 4607 25467 4613
rect 25179 4573 25191 4576
rect 25133 4567 25191 4573
rect 25409 4573 25421 4607
rect 25455 4604 25467 4607
rect 25516 4604 25544 4700
rect 25976 4672 26004 4768
rect 26326 4700 26332 4752
rect 26384 4700 26390 4752
rect 25700 4644 26188 4672
rect 25700 4613 25728 4644
rect 26160 4613 26188 4644
rect 26234 4632 26240 4684
rect 26292 4632 26298 4684
rect 25455 4576 25544 4604
rect 25685 4607 25743 4613
rect 25455 4573 25467 4576
rect 25409 4567 25467 4573
rect 25685 4573 25697 4607
rect 25731 4573 25743 4607
rect 25685 4567 25743 4573
rect 25961 4607 26019 4613
rect 25961 4573 25973 4607
rect 26007 4573 26019 4607
rect 25961 4567 26019 4573
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4573 26203 4607
rect 26145 4567 26203 4573
rect 22388 4536 22416 4564
rect 22066 4508 22416 4536
rect 22480 4508 23244 4536
rect 22480 4480 22508 4508
rect 20070 4468 20076 4480
rect 19996 4440 20076 4468
rect 20070 4428 20076 4440
rect 20128 4428 20134 4480
rect 20254 4428 20260 4480
rect 20312 4468 20318 4480
rect 20441 4471 20499 4477
rect 20441 4468 20453 4471
rect 20312 4440 20453 4468
rect 20312 4428 20318 4440
rect 20441 4437 20453 4440
rect 20487 4437 20499 4471
rect 20441 4431 20499 4437
rect 20898 4428 20904 4480
rect 20956 4468 20962 4480
rect 20993 4471 21051 4477
rect 20993 4468 21005 4471
rect 20956 4440 21005 4468
rect 20956 4428 20962 4440
rect 20993 4437 21005 4440
rect 21039 4437 21051 4471
rect 20993 4431 21051 4437
rect 21082 4428 21088 4480
rect 21140 4468 21146 4480
rect 22005 4471 22063 4477
rect 22005 4468 22017 4471
rect 21140 4440 22017 4468
rect 21140 4428 21146 4440
rect 22005 4437 22017 4440
rect 22051 4437 22063 4471
rect 22005 4431 22063 4437
rect 22278 4428 22284 4480
rect 22336 4428 22342 4480
rect 22462 4428 22468 4480
rect 22520 4428 22526 4480
rect 22646 4428 22652 4480
rect 22704 4428 22710 4480
rect 22738 4428 22744 4480
rect 22796 4468 22802 4480
rect 23216 4477 23244 4508
rect 22925 4471 22983 4477
rect 22925 4468 22937 4471
rect 22796 4440 22937 4468
rect 22796 4428 22802 4440
rect 22925 4437 22937 4440
rect 22971 4437 22983 4471
rect 22925 4431 22983 4437
rect 23201 4471 23259 4477
rect 23201 4437 23213 4471
rect 23247 4437 23259 4471
rect 23201 4431 23259 4437
rect 23477 4471 23535 4477
rect 23477 4437 23489 4471
rect 23523 4468 23535 4471
rect 23584 4468 23612 4564
rect 24118 4496 24124 4548
rect 24176 4536 24182 4548
rect 24176 4508 24440 4536
rect 24176 4496 24182 4508
rect 23523 4440 23612 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 23842 4428 23848 4480
rect 23900 4428 23906 4480
rect 24412 4477 24440 4508
rect 24397 4471 24455 4477
rect 24397 4437 24409 4471
rect 24443 4437 24455 4471
rect 24504 4468 24532 4564
rect 25038 4496 25044 4548
rect 25096 4536 25102 4548
rect 25976 4536 26004 4567
rect 26252 4536 26280 4632
rect 27816 4613 27844 4780
rect 28166 4768 28172 4780
rect 28224 4768 28230 4820
rect 28442 4768 28448 4820
rect 28500 4768 28506 4820
rect 28718 4768 28724 4820
rect 28776 4768 28782 4820
rect 28902 4768 28908 4820
rect 28960 4768 28966 4820
rect 28994 4768 29000 4820
rect 29052 4768 29058 4820
rect 30558 4768 30564 4820
rect 30616 4768 30622 4820
rect 30834 4768 30840 4820
rect 30892 4768 30898 4820
rect 31110 4768 31116 4820
rect 31168 4768 31174 4820
rect 31665 4811 31723 4817
rect 31665 4777 31677 4811
rect 31711 4808 31723 4811
rect 33502 4808 33508 4820
rect 31711 4780 33508 4808
rect 31711 4777 31723 4780
rect 31665 4771 31723 4777
rect 33502 4768 33508 4780
rect 33560 4768 33566 4820
rect 34422 4768 34428 4820
rect 34480 4768 34486 4820
rect 34790 4768 34796 4820
rect 34848 4768 34854 4820
rect 35250 4768 35256 4820
rect 35308 4768 35314 4820
rect 35342 4768 35348 4820
rect 35400 4768 35406 4820
rect 35802 4768 35808 4820
rect 35860 4808 35866 4820
rect 36081 4811 36139 4817
rect 36081 4808 36093 4811
rect 35860 4780 36093 4808
rect 35860 4768 35866 4780
rect 36081 4777 36093 4780
rect 36127 4777 36139 4811
rect 36081 4771 36139 4777
rect 36630 4768 36636 4820
rect 36688 4808 36694 4820
rect 37185 4811 37243 4817
rect 37185 4808 37197 4811
rect 36688 4780 37197 4808
rect 36688 4768 36694 4780
rect 37185 4777 37197 4780
rect 37231 4777 37243 4811
rect 37185 4771 37243 4777
rect 37734 4768 37740 4820
rect 37792 4808 37798 4820
rect 38289 4811 38347 4817
rect 38289 4808 38301 4811
rect 37792 4780 38301 4808
rect 37792 4768 37798 4780
rect 38289 4777 38301 4780
rect 38335 4777 38347 4811
rect 38289 4771 38347 4777
rect 38378 4768 38384 4820
rect 38436 4808 38442 4820
rect 38841 4811 38899 4817
rect 38841 4808 38853 4811
rect 38436 4780 38853 4808
rect 38436 4768 38442 4780
rect 38841 4777 38853 4780
rect 38887 4777 38899 4811
rect 38841 4771 38899 4777
rect 39393 4811 39451 4817
rect 39393 4777 39405 4811
rect 39439 4777 39451 4811
rect 39393 4771 39451 4777
rect 28736 4740 28764 4768
rect 28092 4712 28764 4740
rect 28092 4613 28120 4712
rect 28920 4672 28948 4768
rect 28368 4644 28948 4672
rect 28368 4613 28396 4644
rect 27801 4607 27859 4613
rect 27801 4573 27813 4607
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 28077 4607 28135 4613
rect 28077 4573 28089 4607
rect 28123 4573 28135 4607
rect 28077 4567 28135 4573
rect 28353 4607 28411 4613
rect 28353 4573 28365 4607
rect 28399 4573 28411 4607
rect 28353 4567 28411 4573
rect 28629 4607 28687 4613
rect 28629 4573 28641 4607
rect 28675 4604 28687 4607
rect 28902 4604 28908 4616
rect 28675 4576 28908 4604
rect 28675 4573 28687 4576
rect 28629 4567 28687 4573
rect 28902 4564 28908 4576
rect 28960 4564 28966 4616
rect 29178 4564 29184 4616
rect 29236 4564 29242 4616
rect 29914 4564 29920 4616
rect 29972 4564 29978 4616
rect 30576 4604 30604 4768
rect 30852 4672 30880 4768
rect 31128 4740 31156 4768
rect 31128 4712 31524 4740
rect 30852 4644 31248 4672
rect 31220 4613 31248 4644
rect 31496 4613 31524 4712
rect 31754 4700 31760 4752
rect 31812 4700 31818 4752
rect 31846 4700 31852 4752
rect 31904 4700 31910 4752
rect 32030 4700 32036 4752
rect 32088 4700 32094 4752
rect 33045 4743 33103 4749
rect 33045 4709 33057 4743
rect 33091 4709 33103 4743
rect 33045 4703 33103 4709
rect 34149 4743 34207 4749
rect 34149 4709 34161 4743
rect 34195 4740 34207 4743
rect 35360 4740 35388 4768
rect 34195 4712 35388 4740
rect 34195 4709 34207 4712
rect 34149 4703 34207 4709
rect 30837 4607 30895 4613
rect 30837 4604 30849 4607
rect 30576 4576 30849 4604
rect 30837 4573 30849 4576
rect 30883 4573 30895 4607
rect 30837 4567 30895 4573
rect 31205 4607 31263 4613
rect 31205 4573 31217 4607
rect 31251 4573 31263 4607
rect 31205 4567 31263 4573
rect 31481 4607 31539 4613
rect 31481 4573 31493 4607
rect 31527 4573 31539 4607
rect 31772 4604 31800 4700
rect 31864 4672 31892 4700
rect 33060 4672 33088 4703
rect 36170 4700 36176 4752
rect 36228 4740 36234 4752
rect 36725 4743 36783 4749
rect 36725 4740 36737 4743
rect 36228 4712 36737 4740
rect 36228 4700 36234 4712
rect 36725 4709 36737 4712
rect 36771 4709 36783 4743
rect 36725 4703 36783 4709
rect 37274 4700 37280 4752
rect 37332 4740 37338 4752
rect 37829 4743 37887 4749
rect 37829 4740 37841 4743
rect 37332 4712 37841 4740
rect 37332 4700 37338 4712
rect 37829 4709 37841 4712
rect 37875 4709 37887 4743
rect 37829 4703 37887 4709
rect 38562 4700 38568 4752
rect 38620 4740 38626 4752
rect 39408 4740 39436 4771
rect 39666 4768 39672 4820
rect 39724 4808 39730 4820
rect 40037 4811 40095 4817
rect 40037 4808 40049 4811
rect 39724 4780 40049 4808
rect 39724 4768 39730 4780
rect 40037 4777 40049 4780
rect 40083 4777 40095 4811
rect 40037 4771 40095 4777
rect 40218 4768 40224 4820
rect 40276 4808 40282 4820
rect 41141 4811 41199 4817
rect 41141 4808 41153 4811
rect 40276 4780 41153 4808
rect 40276 4768 40282 4780
rect 41141 4777 41153 4780
rect 41187 4777 41199 4811
rect 41141 4771 41199 4777
rect 38620 4712 39436 4740
rect 38620 4700 38626 4712
rect 39942 4700 39948 4752
rect 40000 4740 40006 4752
rect 40681 4743 40739 4749
rect 40681 4740 40693 4743
rect 40000 4712 40693 4740
rect 40000 4700 40006 4712
rect 40681 4709 40693 4712
rect 40727 4709 40739 4743
rect 40681 4703 40739 4709
rect 31864 4644 32260 4672
rect 33060 4644 35894 4672
rect 32232 4613 32260 4644
rect 31849 4607 31907 4613
rect 31849 4604 31861 4607
rect 31772 4576 31861 4604
rect 31481 4567 31539 4573
rect 31849 4573 31861 4576
rect 31895 4573 31907 4607
rect 31849 4567 31907 4573
rect 32217 4607 32275 4613
rect 32217 4573 32229 4607
rect 32263 4573 32275 4607
rect 32861 4607 32919 4613
rect 32861 4604 32873 4607
rect 32217 4567 32275 4573
rect 32324 4576 32873 4604
rect 25096 4508 25912 4536
rect 25976 4508 26280 4536
rect 26344 4508 27936 4536
rect 25096 4496 25102 4508
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 24504 4440 24685 4468
rect 24397 4431 24455 4437
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 24673 4431 24731 4437
rect 24946 4428 24952 4480
rect 25004 4428 25010 4480
rect 25130 4428 25136 4480
rect 25188 4468 25194 4480
rect 25225 4471 25283 4477
rect 25225 4468 25237 4471
rect 25188 4440 25237 4468
rect 25188 4428 25194 4440
rect 25225 4437 25237 4440
rect 25271 4437 25283 4471
rect 25225 4431 25283 4437
rect 25498 4428 25504 4480
rect 25556 4428 25562 4480
rect 25884 4468 25912 4508
rect 26344 4468 26372 4508
rect 27908 4477 27936 4508
rect 27982 4496 27988 4548
rect 28040 4536 28046 4548
rect 28040 4508 31754 4536
rect 28040 4496 28046 4508
rect 25884 4440 26372 4468
rect 27893 4471 27951 4477
rect 27893 4437 27905 4471
rect 27939 4437 27951 4471
rect 27893 4431 27951 4437
rect 28074 4428 28080 4480
rect 28132 4468 28138 4480
rect 28169 4471 28227 4477
rect 28169 4468 28181 4471
rect 28132 4440 28181 4468
rect 28132 4428 28138 4440
rect 28169 4437 28181 4440
rect 28215 4437 28227 4471
rect 28169 4431 28227 4437
rect 29730 4428 29736 4480
rect 29788 4428 29794 4480
rect 31018 4428 31024 4480
rect 31076 4428 31082 4480
rect 31386 4428 31392 4480
rect 31444 4428 31450 4480
rect 31726 4468 31754 4508
rect 32324 4468 32352 4576
rect 32861 4573 32873 4576
rect 32907 4573 32919 4607
rect 32861 4567 32919 4573
rect 33226 4564 33232 4616
rect 33284 4604 33290 4616
rect 33965 4607 34023 4613
rect 33965 4604 33977 4607
rect 33284 4576 33977 4604
rect 33284 4564 33290 4576
rect 33965 4573 33977 4576
rect 34011 4573 34023 4607
rect 33965 4567 34023 4573
rect 34241 4607 34299 4613
rect 34241 4573 34253 4607
rect 34287 4604 34299 4607
rect 34422 4604 34428 4616
rect 34287 4576 34428 4604
rect 34287 4573 34299 4576
rect 34241 4567 34299 4573
rect 34422 4564 34428 4576
rect 34480 4564 34486 4616
rect 35066 4564 35072 4616
rect 35124 4564 35130 4616
rect 35158 4564 35164 4616
rect 35216 4604 35222 4616
rect 35345 4607 35403 4613
rect 35345 4604 35357 4607
rect 35216 4576 35357 4604
rect 35216 4564 35222 4576
rect 35345 4573 35357 4576
rect 35391 4573 35403 4607
rect 35345 4567 35403 4573
rect 35618 4564 35624 4616
rect 35676 4564 35682 4616
rect 35866 4604 35894 4644
rect 40126 4632 40132 4684
rect 40184 4672 40190 4684
rect 40184 4644 42104 4672
rect 40184 4632 40190 4644
rect 38197 4607 38255 4613
rect 38197 4604 38209 4607
rect 35866 4576 38209 4604
rect 38197 4573 38209 4576
rect 38243 4573 38255 4607
rect 38197 4567 38255 4573
rect 40310 4564 40316 4616
rect 40368 4604 40374 4616
rect 41049 4607 41107 4613
rect 41049 4604 41061 4607
rect 40368 4576 41061 4604
rect 40368 4564 40374 4576
rect 41049 4573 41061 4576
rect 41095 4573 41107 4607
rect 41049 4567 41107 4573
rect 41506 4564 41512 4616
rect 41564 4564 41570 4616
rect 42076 4613 42104 4644
rect 42061 4607 42119 4613
rect 42061 4573 42073 4607
rect 42107 4573 42119 4607
rect 42061 4567 42119 4573
rect 35989 4539 36047 4545
rect 35989 4536 36001 4539
rect 35544 4508 36001 4536
rect 31726 4440 32352 4468
rect 32401 4471 32459 4477
rect 32401 4437 32413 4471
rect 32447 4468 32459 4471
rect 32950 4468 32956 4480
rect 32447 4440 32956 4468
rect 32447 4437 32459 4440
rect 32401 4431 32459 4437
rect 32950 4428 32956 4440
rect 33008 4428 33014 4480
rect 35544 4477 35572 4508
rect 35989 4505 36001 4508
rect 36035 4505 36047 4539
rect 35989 4499 36047 4505
rect 36541 4539 36599 4545
rect 36541 4505 36553 4539
rect 36587 4505 36599 4539
rect 36541 4499 36599 4505
rect 35529 4471 35587 4477
rect 35529 4437 35541 4471
rect 35575 4437 35587 4471
rect 35529 4431 35587 4437
rect 35805 4471 35863 4477
rect 35805 4437 35817 4471
rect 35851 4468 35863 4471
rect 36556 4468 36584 4499
rect 37090 4496 37096 4548
rect 37148 4496 37154 4548
rect 37642 4496 37648 4548
rect 37700 4496 37706 4548
rect 37734 4496 37740 4548
rect 37792 4536 37798 4548
rect 38749 4539 38807 4545
rect 38749 4536 38761 4539
rect 37792 4508 38761 4536
rect 37792 4496 37798 4508
rect 38749 4505 38761 4508
rect 38795 4505 38807 4539
rect 38749 4499 38807 4505
rect 39298 4496 39304 4548
rect 39356 4496 39362 4548
rect 39942 4496 39948 4548
rect 40000 4496 40006 4548
rect 40497 4539 40555 4545
rect 40497 4505 40509 4539
rect 40543 4505 40555 4539
rect 40497 4499 40555 4505
rect 35851 4440 36584 4468
rect 35851 4437 35863 4440
rect 35805 4431 35863 4437
rect 38654 4428 38660 4480
rect 38712 4468 38718 4480
rect 40512 4468 40540 4499
rect 38712 4440 40540 4468
rect 38712 4428 38718 4440
rect 41690 4428 41696 4480
rect 41748 4428 41754 4480
rect 42245 4471 42303 4477
rect 42245 4437 42257 4471
rect 42291 4468 42303 4471
rect 42702 4468 42708 4480
rect 42291 4440 42708 4468
rect 42291 4437 42303 4440
rect 42245 4431 42303 4437
rect 42702 4428 42708 4440
rect 42760 4428 42766 4480
rect 1104 4378 45051 4400
rect 1104 4326 11896 4378
rect 11948 4326 11960 4378
rect 12012 4326 12024 4378
rect 12076 4326 12088 4378
rect 12140 4326 12152 4378
rect 12204 4326 22843 4378
rect 22895 4326 22907 4378
rect 22959 4326 22971 4378
rect 23023 4326 23035 4378
rect 23087 4326 23099 4378
rect 23151 4326 33790 4378
rect 33842 4326 33854 4378
rect 33906 4326 33918 4378
rect 33970 4326 33982 4378
rect 34034 4326 34046 4378
rect 34098 4326 44737 4378
rect 44789 4326 44801 4378
rect 44853 4326 44865 4378
rect 44917 4326 44929 4378
rect 44981 4326 44993 4378
rect 45045 4326 45051 4378
rect 1104 4304 45051 4326
rect 10778 4224 10784 4276
rect 10836 4264 10842 4276
rect 10873 4267 10931 4273
rect 10873 4264 10885 4267
rect 10836 4236 10885 4264
rect 10836 4224 10842 4236
rect 10873 4233 10885 4236
rect 10919 4233 10931 4267
rect 10873 4227 10931 4233
rect 11146 4224 11152 4276
rect 11204 4224 11210 4276
rect 11330 4224 11336 4276
rect 11388 4264 11394 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11388 4236 12173 4264
rect 11388 4224 11394 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 12618 4224 12624 4276
rect 12676 4224 12682 4276
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13541 4267 13599 4273
rect 13541 4264 13553 4267
rect 13136 4236 13553 4264
rect 13136 4224 13142 4236
rect 13541 4233 13553 4236
rect 13587 4233 13599 4267
rect 13541 4227 13599 4233
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 16025 4267 16083 4273
rect 16025 4264 16037 4267
rect 15436 4236 16037 4264
rect 15436 4224 15442 4236
rect 16025 4233 16037 4236
rect 16071 4233 16083 4267
rect 16025 4227 16083 4233
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 17037 4267 17095 4273
rect 17037 4264 17049 4267
rect 16632 4236 17049 4264
rect 16632 4224 16638 4236
rect 17037 4233 17049 4236
rect 17083 4233 17095 4267
rect 17037 4227 17095 4233
rect 17218 4224 17224 4276
rect 17276 4224 17282 4276
rect 17770 4224 17776 4276
rect 17828 4224 17834 4276
rect 18046 4224 18052 4276
rect 18104 4224 18110 4276
rect 18598 4224 18604 4276
rect 18656 4224 18662 4276
rect 18874 4224 18880 4276
rect 18932 4224 18938 4276
rect 18966 4224 18972 4276
rect 19024 4264 19030 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 19024 4236 19165 4264
rect 19024 4224 19030 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19153 4227 19211 4233
rect 19521 4267 19579 4273
rect 19521 4233 19533 4267
rect 19567 4264 19579 4267
rect 19702 4264 19708 4276
rect 19567 4236 19708 4264
rect 19567 4233 19579 4236
rect 19521 4227 19579 4233
rect 19702 4224 19708 4236
rect 19760 4224 19766 4276
rect 25038 4264 25044 4276
rect 19812 4236 21404 4264
rect 9217 4199 9275 4205
rect 9217 4165 9229 4199
rect 9263 4196 9275 4199
rect 11238 4196 11244 4208
rect 9263 4168 11244 4196
rect 9263 4165 9275 4168
rect 9217 4159 9275 4165
rect 11238 4156 11244 4168
rect 11296 4156 11302 4208
rect 11790 4156 11796 4208
rect 11848 4156 11854 4208
rect 12526 4156 12532 4208
rect 12584 4156 12590 4208
rect 13262 4156 13268 4208
rect 13320 4156 13326 4208
rect 13648 4168 13860 4196
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9677 4131 9735 4137
rect 9677 4128 9689 4131
rect 9640 4100 9689 4128
rect 9640 4088 9646 4100
rect 9677 4097 9689 4100
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 11057 4131 11115 4137
rect 10091 4100 11008 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 10980 3924 11008 4100
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11072 4060 11100 4091
rect 11330 4088 11336 4140
rect 11388 4088 11394 4140
rect 12345 4131 12403 4137
rect 12345 4097 12357 4131
rect 12391 4128 12403 4131
rect 12391 4100 12940 4128
rect 12391 4097 12403 4100
rect 12345 4091 12403 4097
rect 12618 4060 12624 4072
rect 11072 4032 12624 4060
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12912 4060 12940 4100
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 13648 4060 13676 4168
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 12912 4032 13676 4060
rect 11974 3952 11980 4004
rect 12032 3952 12038 4004
rect 12250 3952 12256 4004
rect 12308 3992 12314 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 12308 3964 12817 3992
rect 12308 3952 12314 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 12805 3955 12863 3961
rect 13446 3952 13452 4004
rect 13504 3952 13510 4004
rect 13630 3952 13636 4004
rect 13688 3952 13694 4004
rect 13648 3924 13676 3952
rect 10980 3896 13676 3924
rect 13740 3924 13768 4091
rect 13832 4060 13860 4168
rect 13998 4156 14004 4208
rect 14056 4156 14062 4208
rect 14366 4156 14372 4208
rect 14424 4156 14430 4208
rect 15010 4156 15016 4208
rect 15068 4156 15074 4208
rect 15470 4156 15476 4208
rect 15528 4156 15534 4208
rect 17236 4196 17264 4224
rect 19812 4196 19840 4236
rect 20806 4196 20812 4208
rect 17236 4168 19840 4196
rect 19904 4168 20812 4196
rect 14642 4088 14648 4140
rect 14700 4088 14706 4140
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 15657 4131 15715 4137
rect 15657 4097 15669 4131
rect 15703 4128 15715 4131
rect 15746 4128 15752 4140
rect 15703 4100 15752 4128
rect 15703 4097 15715 4100
rect 15657 4091 15715 4097
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 15396 4060 15424 4088
rect 13832 4032 15424 4060
rect 15948 4060 15976 4091
rect 16206 4088 16212 4140
rect 16264 4088 16270 4140
rect 17221 4131 17279 4137
rect 17221 4097 17233 4131
rect 17267 4097 17279 4131
rect 17221 4091 17279 4097
rect 16574 4060 16580 4072
rect 15948 4032 16580 4060
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 14182 3952 14188 4004
rect 14240 3952 14246 4004
rect 14550 3952 14556 4004
rect 14608 3952 14614 4004
rect 16758 3992 16764 4004
rect 15488 3964 16764 3992
rect 15488 3924 15516 3964
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 13740 3896 15516 3924
rect 15562 3884 15568 3936
rect 15620 3924 15626 3936
rect 15749 3927 15807 3933
rect 15749 3924 15761 3927
rect 15620 3896 15761 3924
rect 15620 3884 15626 3896
rect 15749 3893 15761 3896
rect 15795 3893 15807 3927
rect 17236 3924 17264 4091
rect 17954 4088 17960 4140
rect 18012 4088 18018 4140
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4097 18291 4131
rect 18233 4091 18291 4097
rect 17862 4020 17868 4072
rect 17920 4020 17926 4072
rect 18248 4060 18276 4091
rect 18506 4088 18512 4140
rect 18564 4088 18570 4140
rect 18782 4088 18788 4140
rect 18840 4088 18846 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4097 19119 4131
rect 19061 4091 19119 4097
rect 19076 4060 19104 4091
rect 19334 4088 19340 4140
rect 19392 4088 19398 4140
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4097 19763 4131
rect 19705 4091 19763 4097
rect 19426 4060 19432 4072
rect 18248 4032 19012 4060
rect 19076 4032 19432 4060
rect 17880 3992 17908 4020
rect 18325 3995 18383 4001
rect 18325 3992 18337 3995
rect 17880 3964 18337 3992
rect 18325 3961 18337 3964
rect 18371 3961 18383 3995
rect 18984 3992 19012 4032
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 19518 3992 19524 4004
rect 18984 3964 19524 3992
rect 18325 3955 18383 3961
rect 19518 3952 19524 3964
rect 19576 3952 19582 4004
rect 19720 3992 19748 4091
rect 19794 4088 19800 4140
rect 19852 4128 19858 4140
rect 19904 4128 19932 4168
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 20898 4156 20904 4208
rect 20956 4156 20962 4208
rect 21266 4156 21272 4208
rect 21324 4156 21330 4208
rect 21376 4196 21404 4236
rect 21560 4236 25044 4264
rect 21560 4196 21588 4236
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 25498 4224 25504 4276
rect 25556 4224 25562 4276
rect 25866 4264 25872 4276
rect 25608 4236 25872 4264
rect 21376 4168 21588 4196
rect 21910 4156 21916 4208
rect 21968 4196 21974 4208
rect 25516 4196 25544 4224
rect 21968 4168 25544 4196
rect 21968 4156 21974 4168
rect 19852 4100 19932 4128
rect 20441 4131 20499 4137
rect 19852 4088 19858 4100
rect 20441 4097 20453 4131
rect 20487 4128 20499 4131
rect 20916 4128 20944 4156
rect 20487 4100 20944 4128
rect 20993 4131 21051 4137
rect 20487 4097 20499 4100
rect 20441 4091 20499 4097
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21284 4128 21312 4156
rect 21039 4100 21312 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 23934 4088 23940 4140
rect 23992 4128 23998 4140
rect 25608 4128 25636 4236
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 26234 4224 26240 4276
rect 26292 4224 26298 4276
rect 31018 4224 31024 4276
rect 31076 4224 31082 4276
rect 31386 4224 31392 4276
rect 31444 4264 31450 4276
rect 34514 4264 34520 4276
rect 31444 4236 34520 4264
rect 31444 4224 31450 4236
rect 34514 4224 34520 4236
rect 34572 4224 34578 4276
rect 35897 4267 35955 4273
rect 35897 4233 35909 4267
rect 35943 4233 35955 4267
rect 35897 4227 35955 4233
rect 36173 4267 36231 4273
rect 36173 4233 36185 4267
rect 36219 4264 36231 4267
rect 37090 4264 37096 4276
rect 36219 4236 37096 4264
rect 36219 4233 36231 4236
rect 36173 4227 36231 4233
rect 23992 4100 25636 4128
rect 26252 4128 26280 4224
rect 31036 4196 31064 4224
rect 34330 4196 34336 4208
rect 31036 4168 34336 4196
rect 34330 4156 34336 4168
rect 34388 4156 34394 4208
rect 35912 4196 35940 4227
rect 37090 4224 37096 4236
rect 37148 4224 37154 4276
rect 36722 4196 36728 4208
rect 35912 4168 36728 4196
rect 36722 4156 36728 4168
rect 36780 4156 36786 4208
rect 26421 4131 26479 4137
rect 26421 4128 26433 4131
rect 26252 4100 26433 4128
rect 23992 4088 23998 4100
rect 26421 4097 26433 4100
rect 26467 4097 26479 4131
rect 26421 4091 26479 4097
rect 30466 4088 30472 4140
rect 30524 4128 30530 4140
rect 35437 4131 35495 4137
rect 35437 4128 35449 4131
rect 30524 4100 35449 4128
rect 30524 4088 30530 4100
rect 35437 4097 35449 4100
rect 35483 4097 35495 4131
rect 35437 4091 35495 4097
rect 35710 4088 35716 4140
rect 35768 4088 35774 4140
rect 35986 4088 35992 4140
rect 36044 4088 36050 4140
rect 36262 4088 36268 4140
rect 36320 4088 36326 4140
rect 36538 4088 36544 4140
rect 36596 4088 36602 4140
rect 39114 4088 39120 4140
rect 39172 4088 39178 4140
rect 39853 4131 39911 4137
rect 39853 4097 39865 4131
rect 39899 4097 39911 4131
rect 39853 4091 39911 4097
rect 40589 4131 40647 4137
rect 40589 4097 40601 4131
rect 40635 4097 40647 4131
rect 40589 4091 40647 4097
rect 24394 4020 24400 4072
rect 24452 4060 24458 4072
rect 26694 4060 26700 4072
rect 24452 4032 26700 4060
rect 24452 4020 24458 4032
rect 26694 4020 26700 4032
rect 26752 4060 26758 4072
rect 27338 4060 27344 4072
rect 26752 4032 27344 4060
rect 26752 4020 26758 4032
rect 27338 4020 27344 4032
rect 27396 4020 27402 4072
rect 33686 4020 33692 4072
rect 33744 4060 33750 4072
rect 39868 4060 39896 4091
rect 33744 4032 39896 4060
rect 33744 4020 33750 4032
rect 26234 3992 26240 4004
rect 19720 3964 26240 3992
rect 26234 3952 26240 3964
rect 26292 3992 26298 4004
rect 26510 3992 26516 4004
rect 26292 3964 26516 3992
rect 26292 3952 26298 3964
rect 26510 3952 26516 3964
rect 26568 3952 26574 4004
rect 35621 3995 35679 4001
rect 35621 3961 35633 3995
rect 35667 3992 35679 3995
rect 36078 3992 36084 4004
rect 35667 3964 36084 3992
rect 35667 3961 35679 3964
rect 35621 3955 35679 3961
rect 36078 3952 36084 3964
rect 36136 3952 36142 4004
rect 36449 3995 36507 4001
rect 36449 3961 36461 3995
rect 36495 3992 36507 3995
rect 37182 3992 37188 4004
rect 36495 3964 37188 3992
rect 36495 3961 36507 3964
rect 36449 3955 36507 3961
rect 37182 3952 37188 3964
rect 37240 3952 37246 4004
rect 38194 3952 38200 4004
rect 38252 3992 38258 4004
rect 40604 3992 40632 4091
rect 38252 3964 40632 3992
rect 38252 3952 38258 3964
rect 19886 3924 19892 3936
rect 17236 3896 19892 3924
rect 15749 3887 15807 3893
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 19978 3884 19984 3936
rect 20036 3924 20042 3936
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 20036 3896 20269 3924
rect 20036 3884 20042 3896
rect 20257 3893 20269 3896
rect 20303 3893 20315 3927
rect 20257 3887 20315 3893
rect 20806 3884 20812 3936
rect 20864 3884 20870 3936
rect 26605 3927 26663 3933
rect 26605 3893 26617 3927
rect 26651 3924 26663 3927
rect 33134 3924 33140 3936
rect 26651 3896 33140 3924
rect 26651 3893 26663 3896
rect 26605 3887 26663 3893
rect 33134 3884 33140 3896
rect 33192 3884 33198 3936
rect 36725 3927 36783 3933
rect 36725 3893 36737 3927
rect 36771 3924 36783 3927
rect 37274 3924 37280 3936
rect 36771 3896 37280 3924
rect 36771 3893 36783 3896
rect 36725 3887 36783 3893
rect 37274 3884 37280 3896
rect 37332 3884 37338 3936
rect 39301 3927 39359 3933
rect 39301 3893 39313 3927
rect 39347 3924 39359 3927
rect 39666 3924 39672 3936
rect 39347 3896 39672 3924
rect 39347 3893 39359 3896
rect 39301 3887 39359 3893
rect 39666 3884 39672 3896
rect 39724 3884 39730 3936
rect 40037 3927 40095 3933
rect 40037 3893 40049 3927
rect 40083 3924 40095 3927
rect 40402 3924 40408 3936
rect 40083 3896 40408 3924
rect 40083 3893 40095 3896
rect 40037 3887 40095 3893
rect 40402 3884 40408 3896
rect 40460 3884 40466 3936
rect 40773 3927 40831 3933
rect 40773 3893 40785 3927
rect 40819 3924 40831 3927
rect 41414 3924 41420 3936
rect 40819 3896 41420 3924
rect 40819 3893 40831 3896
rect 40773 3887 40831 3893
rect 41414 3884 41420 3896
rect 41472 3884 41478 3936
rect 1104 3834 44896 3856
rect 1104 3782 6423 3834
rect 6475 3782 6487 3834
rect 6539 3782 6551 3834
rect 6603 3782 6615 3834
rect 6667 3782 6679 3834
rect 6731 3782 17370 3834
rect 17422 3782 17434 3834
rect 17486 3782 17498 3834
rect 17550 3782 17562 3834
rect 17614 3782 17626 3834
rect 17678 3782 28317 3834
rect 28369 3782 28381 3834
rect 28433 3782 28445 3834
rect 28497 3782 28509 3834
rect 28561 3782 28573 3834
rect 28625 3782 39264 3834
rect 39316 3782 39328 3834
rect 39380 3782 39392 3834
rect 39444 3782 39456 3834
rect 39508 3782 39520 3834
rect 39572 3782 44896 3834
rect 1104 3760 44896 3782
rect 11330 3680 11336 3732
rect 11388 3720 11394 3732
rect 11388 3692 12434 3720
rect 11388 3680 11394 3692
rect 12406 3448 12434 3692
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 16117 3723 16175 3729
rect 16117 3720 16129 3723
rect 14792 3692 16129 3720
rect 14792 3680 14798 3692
rect 16117 3689 16129 3692
rect 16163 3689 16175 3723
rect 16117 3683 16175 3689
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 27246 3720 27252 3732
rect 18840 3692 27252 3720
rect 18840 3680 18846 3692
rect 27246 3680 27252 3692
rect 27304 3680 27310 3732
rect 27338 3680 27344 3732
rect 27396 3720 27402 3732
rect 33781 3723 33839 3729
rect 27396 3692 31754 3720
rect 27396 3680 27402 3692
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 17218 3652 17224 3664
rect 13044 3624 17224 3652
rect 13044 3612 13050 3624
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 19334 3612 19340 3664
rect 19392 3612 19398 3664
rect 19426 3612 19432 3664
rect 19484 3612 19490 3664
rect 26881 3655 26939 3661
rect 26881 3652 26893 3655
rect 26804 3624 26893 3652
rect 12618 3476 12624 3528
rect 12676 3516 12682 3528
rect 16301 3519 16359 3525
rect 12676 3488 15884 3516
rect 12676 3476 12682 3488
rect 15746 3448 15752 3460
rect 12406 3420 15752 3448
rect 15746 3408 15752 3420
rect 15804 3408 15810 3460
rect 15856 3448 15884 3488
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 17126 3516 17132 3528
rect 16347 3488 17132 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 19352 3516 19380 3612
rect 19444 3584 19472 3612
rect 19444 3556 24532 3584
rect 24394 3516 24400 3528
rect 19352 3488 24400 3516
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 20714 3448 20720 3460
rect 15856 3420 20720 3448
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 24504 3448 24532 3556
rect 26234 3544 26240 3596
rect 26292 3544 26298 3596
rect 26252 3516 26280 3544
rect 26697 3519 26755 3525
rect 26697 3516 26709 3519
rect 26252 3488 26709 3516
rect 26697 3485 26709 3488
rect 26743 3485 26755 3519
rect 26804 3516 26832 3624
rect 26881 3621 26893 3624
rect 26927 3621 26939 3655
rect 31726 3652 31754 3692
rect 33781 3689 33793 3723
rect 33827 3720 33839 3723
rect 34606 3720 34612 3732
rect 33827 3692 34612 3720
rect 33827 3689 33839 3692
rect 33781 3683 33839 3689
rect 34606 3680 34612 3692
rect 34664 3680 34670 3732
rect 36538 3720 36544 3732
rect 35866 3692 36544 3720
rect 35866 3652 35894 3692
rect 36538 3680 36544 3692
rect 36596 3680 36602 3732
rect 38194 3680 38200 3732
rect 38252 3680 38258 3732
rect 39114 3680 39120 3732
rect 39172 3680 39178 3732
rect 31726 3624 35894 3652
rect 26881 3615 26939 3621
rect 33410 3544 33416 3596
rect 33468 3584 33474 3596
rect 38212 3584 38240 3680
rect 33468 3556 38240 3584
rect 33468 3544 33474 3556
rect 31665 3519 31723 3525
rect 26804 3488 29316 3516
rect 26697 3479 26755 3485
rect 26970 3448 26976 3460
rect 24504 3420 26976 3448
rect 26970 3408 26976 3420
rect 27028 3408 27034 3460
rect 29288 3448 29316 3488
rect 31665 3485 31677 3519
rect 31711 3516 31723 3519
rect 32490 3516 32496 3528
rect 31711 3488 32496 3516
rect 31711 3485 31723 3488
rect 31665 3479 31723 3485
rect 32490 3476 32496 3488
rect 32548 3476 32554 3528
rect 33594 3476 33600 3528
rect 33652 3476 33658 3528
rect 34146 3476 34152 3528
rect 34204 3516 34210 3528
rect 39132 3516 39160 3680
rect 34204 3488 39160 3516
rect 34204 3476 34210 3488
rect 34238 3448 34244 3460
rect 29288 3420 34244 3448
rect 34238 3408 34244 3420
rect 34296 3408 34302 3460
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 27890 3380 27896 3392
rect 18012 3352 27896 3380
rect 18012 3340 18018 3352
rect 27890 3340 27896 3352
rect 27948 3340 27954 3392
rect 31478 3340 31484 3392
rect 31536 3340 31542 3392
rect 1104 3290 45051 3312
rect 1104 3238 11896 3290
rect 11948 3238 11960 3290
rect 12012 3238 12024 3290
rect 12076 3238 12088 3290
rect 12140 3238 12152 3290
rect 12204 3238 22843 3290
rect 22895 3238 22907 3290
rect 22959 3238 22971 3290
rect 23023 3238 23035 3290
rect 23087 3238 23099 3290
rect 23151 3238 33790 3290
rect 33842 3238 33854 3290
rect 33906 3238 33918 3290
rect 33970 3238 33982 3290
rect 34034 3238 34046 3290
rect 34098 3238 44737 3290
rect 44789 3238 44801 3290
rect 44853 3238 44865 3290
rect 44917 3238 44929 3290
rect 44981 3238 44993 3290
rect 45045 3238 45051 3290
rect 1104 3216 45051 3238
rect 2593 3179 2651 3185
rect 2593 3145 2605 3179
rect 2639 3176 2651 3179
rect 2682 3176 2688 3188
rect 2639 3148 2688 3176
rect 2639 3145 2651 3148
rect 2593 3139 2651 3145
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 12710 3136 12716 3188
rect 12768 3136 12774 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15565 3179 15623 3185
rect 15565 3176 15577 3179
rect 15344 3148 15577 3176
rect 15344 3136 15350 3148
rect 15565 3145 15577 3148
rect 15611 3145 15623 3179
rect 15565 3139 15623 3145
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 15841 3179 15899 3185
rect 15841 3176 15853 3179
rect 15712 3148 15853 3176
rect 15712 3136 15718 3148
rect 15841 3145 15853 3148
rect 15887 3145 15899 3179
rect 15841 3139 15899 3145
rect 16301 3179 16359 3185
rect 16301 3145 16313 3179
rect 16347 3176 16359 3179
rect 16482 3176 16488 3188
rect 16347 3148 16488 3176
rect 16347 3145 16359 3148
rect 16301 3139 16359 3145
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 16853 3179 16911 3185
rect 16853 3176 16865 3179
rect 16724 3148 16865 3176
rect 16724 3136 16730 3148
rect 16853 3145 16865 3148
rect 16899 3145 16911 3179
rect 16853 3139 16911 3145
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 17129 3179 17187 3185
rect 17129 3176 17141 3179
rect 17000 3148 17141 3176
rect 17000 3136 17006 3148
rect 17129 3145 17141 3148
rect 17175 3145 17187 3179
rect 17129 3139 17187 3145
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 18564 3148 22094 3176
rect 18564 3136 18570 3148
rect 17770 3108 17776 3120
rect 12912 3080 17776 3108
rect 842 3000 848 3052
rect 900 3040 906 3052
rect 1489 3043 1547 3049
rect 1489 3040 1501 3043
rect 900 3012 1501 3040
rect 900 3000 906 3012
rect 1489 3009 1501 3012
rect 1535 3009 1547 3043
rect 1489 3003 1547 3009
rect 2498 3000 2504 3052
rect 2556 3000 2562 3052
rect 4154 3000 4160 3052
rect 4212 3000 4218 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 10318 3000 10324 3052
rect 10376 3000 10382 3052
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 11238 3000 11244 3052
rect 11296 3000 11302 3052
rect 12912 3049 12940 3080
rect 17770 3068 17776 3080
rect 17828 3068 17834 3120
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 12897 3003 12955 3009
rect 15749 3043 15807 3049
rect 15749 3009 15761 3043
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3009 16083 3043
rect 16025 3003 16083 3009
rect 3878 2932 3884 2984
rect 3936 2932 3942 2984
rect 1670 2864 1676 2916
rect 1728 2864 1734 2916
rect 5626 2864 5632 2916
rect 5684 2864 5690 2916
rect 10502 2864 10508 2916
rect 10560 2864 10566 2916
rect 13170 2864 13176 2916
rect 13228 2864 13234 2916
rect 15764 2904 15792 3003
rect 16040 2972 16068 3003
rect 16206 3000 16212 3052
rect 16264 3000 16270 3052
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17313 3043 17371 3049
rect 17313 3009 17325 3043
rect 17359 3040 17371 3043
rect 20162 3040 20168 3052
rect 17359 3012 20168 3040
rect 17359 3009 17371 3012
rect 17313 3003 17371 3009
rect 16758 2972 16764 2984
rect 16040 2944 16764 2972
rect 16758 2932 16764 2944
rect 16816 2932 16822 2984
rect 17052 2972 17080 3003
rect 20162 3000 20168 3012
rect 20220 3000 20226 3052
rect 22066 3040 22094 3148
rect 23382 3136 23388 3188
rect 23440 3136 23446 3188
rect 24210 3136 24216 3188
rect 24268 3136 24274 3188
rect 25317 3179 25375 3185
rect 25317 3145 25329 3179
rect 25363 3145 25375 3179
rect 25317 3139 25375 3145
rect 23400 3108 23428 3136
rect 25332 3108 25360 3139
rect 25406 3136 25412 3188
rect 25464 3176 25470 3188
rect 26973 3179 27031 3185
rect 26973 3176 26985 3179
rect 25464 3148 26985 3176
rect 25464 3136 25470 3148
rect 26973 3145 26985 3148
rect 27019 3145 27031 3179
rect 26973 3139 27031 3145
rect 31938 3136 31944 3188
rect 31996 3136 32002 3188
rect 32306 3136 32312 3188
rect 32364 3136 32370 3188
rect 32401 3179 32459 3185
rect 32401 3145 32413 3179
rect 32447 3176 32459 3179
rect 32953 3179 33011 3185
rect 32447 3148 32904 3176
rect 32447 3145 32459 3148
rect 32401 3139 32459 3145
rect 23400 3080 25360 3108
rect 23934 3040 23940 3052
rect 22066 3012 23940 3040
rect 23934 3000 23940 3012
rect 23992 3000 23998 3052
rect 24026 3000 24032 3052
rect 24084 3000 24090 3052
rect 25498 3000 25504 3052
rect 25556 3000 25562 3052
rect 26234 3000 26240 3052
rect 26292 3000 26298 3052
rect 27154 3000 27160 3052
rect 27212 3000 27218 3052
rect 27706 3000 27712 3052
rect 27764 3000 27770 3052
rect 31956 3040 31984 3136
rect 32324 3108 32352 3136
rect 32324 3080 32812 3108
rect 32784 3049 32812 3080
rect 32217 3043 32275 3049
rect 32217 3040 32229 3043
rect 31956 3012 32229 3040
rect 32217 3009 32229 3012
rect 32263 3009 32275 3043
rect 32217 3003 32275 3009
rect 32677 3043 32735 3049
rect 32677 3009 32689 3043
rect 32723 3009 32735 3043
rect 32677 3003 32735 3009
rect 32769 3043 32827 3049
rect 32769 3009 32781 3043
rect 32815 3009 32827 3043
rect 32769 3003 32827 3009
rect 19702 2972 19708 2984
rect 17052 2944 19708 2972
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 16850 2904 16856 2916
rect 15764 2876 16856 2904
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 22066 2876 27568 2904
rect 13188 2836 13216 2864
rect 22066 2836 22094 2876
rect 13188 2808 22094 2836
rect 26050 2796 26056 2848
rect 26108 2796 26114 2848
rect 27540 2845 27568 2876
rect 27525 2839 27583 2845
rect 27525 2805 27537 2839
rect 27571 2805 27583 2839
rect 27525 2799 27583 2805
rect 32490 2796 32496 2848
rect 32548 2796 32554 2848
rect 32692 2836 32720 3003
rect 32876 2904 32904 3148
rect 32953 3145 32965 3179
rect 32999 3145 33011 3179
rect 32953 3139 33011 3145
rect 32968 2972 32996 3139
rect 33042 3136 33048 3188
rect 33100 3136 33106 3188
rect 33229 3179 33287 3185
rect 33229 3145 33241 3179
rect 33275 3176 33287 3179
rect 43162 3176 43168 3188
rect 33275 3148 43168 3176
rect 33275 3145 33287 3148
rect 33229 3139 33287 3145
rect 43162 3136 43168 3148
rect 43220 3136 43226 3188
rect 33060 3049 33088 3136
rect 35912 3080 44220 3108
rect 33045 3043 33103 3049
rect 33045 3009 33057 3043
rect 33091 3009 33103 3043
rect 33045 3003 33103 3009
rect 34790 3000 34796 3052
rect 34848 3000 34854 3052
rect 35912 2972 35940 3080
rect 44192 3049 44220 3080
rect 43625 3043 43683 3049
rect 43625 3040 43637 3043
rect 32968 2944 35940 2972
rect 39776 3012 43637 3040
rect 39776 2904 39804 3012
rect 43625 3009 43637 3012
rect 43671 3009 43683 3043
rect 43625 3003 43683 3009
rect 44177 3043 44235 3049
rect 44177 3009 44189 3043
rect 44223 3009 44235 3043
rect 44177 3003 44235 3009
rect 44634 2904 44640 2916
rect 32876 2876 39804 2904
rect 43916 2876 44640 2904
rect 33318 2836 33324 2848
rect 32692 2808 33324 2836
rect 33318 2796 33324 2808
rect 33376 2796 33382 2848
rect 34977 2839 35035 2845
rect 34977 2805 34989 2839
rect 35023 2836 35035 2839
rect 35526 2836 35532 2848
rect 35023 2808 35532 2836
rect 35023 2805 35035 2808
rect 34977 2799 35035 2805
rect 35526 2796 35532 2808
rect 35584 2796 35590 2848
rect 43916 2845 43944 2876
rect 44634 2864 44640 2876
rect 44692 2864 44698 2916
rect 43901 2839 43959 2845
rect 43901 2805 43913 2839
rect 43947 2805 43959 2839
rect 43901 2799 43959 2805
rect 44266 2796 44272 2848
rect 44324 2796 44330 2848
rect 1104 2746 44896 2768
rect 1104 2694 6423 2746
rect 6475 2694 6487 2746
rect 6539 2694 6551 2746
rect 6603 2694 6615 2746
rect 6667 2694 6679 2746
rect 6731 2694 17370 2746
rect 17422 2694 17434 2746
rect 17486 2694 17498 2746
rect 17550 2694 17562 2746
rect 17614 2694 17626 2746
rect 17678 2694 28317 2746
rect 28369 2694 28381 2746
rect 28433 2694 28445 2746
rect 28497 2694 28509 2746
rect 28561 2694 28573 2746
rect 28625 2694 39264 2746
rect 39316 2694 39328 2746
rect 39380 2694 39392 2746
rect 39444 2694 39456 2746
rect 39508 2694 39520 2746
rect 39572 2694 44896 2746
rect 1104 2672 44896 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 1946 2632 1952 2644
rect 1903 2604 1952 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10318 2632 10324 2644
rect 9999 2604 10324 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 10689 2635 10747 2641
rect 10689 2601 10701 2635
rect 10735 2632 10747 2635
rect 11054 2632 11060 2644
rect 10735 2604 11060 2632
rect 10735 2601 10747 2604
rect 10689 2595 10747 2601
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 11790 2632 11796 2644
rect 11747 2604 11796 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 12161 2635 12219 2641
rect 12161 2601 12173 2635
rect 12207 2632 12219 2635
rect 12526 2632 12532 2644
rect 12207 2604 12532 2632
rect 12207 2601 12219 2604
rect 12161 2595 12219 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 13262 2632 13268 2644
rect 12943 2604 13268 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13633 2635 13691 2641
rect 13633 2601 13645 2635
rect 13679 2632 13691 2635
rect 13998 2632 14004 2644
rect 13679 2604 14004 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14366 2592 14372 2644
rect 14424 2592 14430 2644
rect 15105 2635 15163 2641
rect 15105 2601 15117 2635
rect 15151 2632 15163 2635
rect 15470 2632 15476 2644
rect 15151 2604 15476 2632
rect 15151 2601 15163 2604
rect 15105 2595 15163 2601
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 16206 2632 16212 2644
rect 15887 2604 16212 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 16669 2635 16727 2641
rect 16669 2632 16681 2635
rect 16632 2604 16681 2632
rect 16632 2592 16638 2604
rect 16669 2601 16681 2604
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 17126 2592 17132 2644
rect 17184 2592 17190 2644
rect 17218 2592 17224 2644
rect 17276 2592 17282 2644
rect 17770 2592 17776 2644
rect 17828 2632 17834 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 17828 2604 18613 2632
rect 17828 2592 17834 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 18601 2595 18659 2601
rect 19702 2592 19708 2644
rect 19760 2592 19766 2644
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 23017 2635 23075 2641
rect 23017 2632 23029 2635
rect 20220 2604 23029 2632
rect 20220 2592 20226 2604
rect 23017 2601 23029 2604
rect 23063 2601 23075 2635
rect 23017 2595 23075 2601
rect 25498 2592 25504 2644
rect 25556 2632 25562 2644
rect 25961 2635 26019 2641
rect 25961 2632 25973 2635
rect 25556 2604 25973 2632
rect 25556 2592 25562 2604
rect 25961 2601 25973 2604
rect 26007 2601 26019 2635
rect 25961 2595 26019 2601
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 26973 2635 27031 2641
rect 26973 2632 26985 2635
rect 26292 2604 26985 2632
rect 26292 2592 26298 2604
rect 26973 2601 26985 2604
rect 27019 2601 27031 2635
rect 26973 2595 27031 2601
rect 27154 2592 27160 2644
rect 27212 2632 27218 2644
rect 27433 2635 27491 2641
rect 27433 2632 27445 2635
rect 27212 2604 27445 2632
rect 27212 2592 27218 2604
rect 27433 2601 27445 2604
rect 27479 2601 27491 2635
rect 27433 2595 27491 2601
rect 27706 2592 27712 2644
rect 27764 2632 27770 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27764 2604 28181 2632
rect 27764 2592 27770 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 28902 2592 28908 2644
rect 28960 2592 28966 2644
rect 29178 2592 29184 2644
rect 29236 2632 29242 2644
rect 29641 2635 29699 2641
rect 29641 2632 29653 2635
rect 29236 2604 29653 2632
rect 29236 2592 29242 2604
rect 29641 2601 29653 2604
rect 29687 2601 29699 2635
rect 29641 2595 29699 2601
rect 29914 2592 29920 2644
rect 29972 2632 29978 2644
rect 30377 2635 30435 2641
rect 30377 2632 30389 2635
rect 29972 2604 30389 2632
rect 29972 2592 29978 2604
rect 30377 2601 30389 2604
rect 30423 2601 30435 2635
rect 30377 2595 30435 2601
rect 33134 2592 33140 2644
rect 33192 2632 33198 2644
rect 33192 2604 38608 2632
rect 33192 2592 33198 2604
rect 17236 2564 17264 2592
rect 19337 2567 19395 2573
rect 19337 2564 19349 2567
rect 17236 2536 19349 2564
rect 19337 2533 19349 2536
rect 19383 2533 19395 2567
rect 19720 2564 19748 2592
rect 22281 2567 22339 2573
rect 22281 2564 22293 2567
rect 19720 2536 22293 2564
rect 19337 2527 19395 2533
rect 22281 2533 22293 2536
rect 22327 2533 22339 2567
rect 22281 2527 22339 2533
rect 25225 2567 25283 2573
rect 25225 2533 25237 2567
rect 25271 2533 25283 2567
rect 25225 2527 25283 2533
rect 26344 2536 38056 2564
rect 4706 2456 4712 2508
rect 4764 2456 4770 2508
rect 16390 2456 16396 2508
rect 16448 2496 16454 2508
rect 25240 2496 25268 2527
rect 26344 2508 26372 2536
rect 16448 2468 25268 2496
rect 16448 2456 16454 2468
rect 26326 2456 26332 2508
rect 26384 2456 26390 2508
rect 34256 2468 37964 2496
rect 34256 2440 34284 2468
rect 4430 2388 4436 2440
rect 4488 2388 4494 2440
rect 5902 2388 5908 2440
rect 5960 2388 5966 2440
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 10502 2388 10508 2440
rect 10560 2388 10566 2440
rect 11514 2388 11520 2440
rect 11572 2388 11578 2440
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12710 2388 12716 2440
rect 12768 2388 12774 2440
rect 13446 2388 13452 2440
rect 13504 2388 13510 2440
rect 14182 2388 14188 2440
rect 14240 2388 14246 2440
rect 14918 2388 14924 2440
rect 14976 2388 14982 2440
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16632 2400 16865 2428
rect 16632 2388 16638 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17034 2388 17040 2440
rect 17092 2428 17098 2440
rect 17313 2431 17371 2437
rect 17313 2428 17325 2431
rect 17092 2400 17325 2428
rect 17092 2388 17098 2400
rect 17313 2397 17325 2400
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 17828 2400 18061 2428
rect 17828 2388 17834 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 18564 2400 18797 2428
rect 18564 2388 18570 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 19242 2388 19248 2440
rect 19300 2428 19306 2440
rect 19521 2431 19579 2437
rect 19521 2428 19533 2431
rect 19300 2400 19533 2428
rect 19300 2388 19306 2400
rect 19521 2397 19533 2400
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 20990 2388 20996 2440
rect 21048 2388 21054 2440
rect 21450 2388 21456 2440
rect 21508 2428 21514 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21508 2400 22017 2428
rect 21508 2388 21514 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 22186 2388 22192 2440
rect 22244 2428 22250 2440
rect 22465 2431 22523 2437
rect 22465 2428 22477 2431
rect 22244 2400 22477 2428
rect 22244 2388 22250 2400
rect 22465 2397 22477 2400
rect 22511 2397 22523 2431
rect 22465 2391 22523 2397
rect 23198 2388 23204 2440
rect 23256 2388 23262 2440
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 23937 2431 23995 2437
rect 23937 2428 23949 2431
rect 23716 2400 23949 2428
rect 23716 2388 23722 2400
rect 23937 2397 23949 2400
rect 23983 2397 23995 2431
rect 23937 2391 23995 2397
rect 24670 2388 24676 2440
rect 24728 2388 24734 2440
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25409 2431 25467 2437
rect 25409 2428 25421 2431
rect 25188 2400 25421 2428
rect 25188 2388 25194 2400
rect 25409 2397 25421 2400
rect 25455 2397 25467 2431
rect 25409 2391 25467 2397
rect 26142 2388 26148 2440
rect 26200 2388 26206 2440
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 27157 2431 27215 2437
rect 27157 2428 27169 2431
rect 26660 2400 27169 2428
rect 26660 2388 26666 2400
rect 27157 2397 27169 2400
rect 27203 2397 27215 2431
rect 27157 2391 27215 2397
rect 27614 2388 27620 2440
rect 27672 2388 27678 2440
rect 28074 2388 28080 2440
rect 28132 2428 28138 2440
rect 28353 2431 28411 2437
rect 28353 2428 28365 2431
rect 28132 2400 28365 2428
rect 28132 2388 28138 2400
rect 28353 2397 28365 2400
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 28810 2388 28816 2440
rect 28868 2428 28874 2440
rect 29089 2431 29147 2437
rect 29089 2428 29101 2431
rect 28868 2400 29101 2428
rect 28868 2388 28874 2400
rect 29089 2397 29101 2400
rect 29135 2397 29147 2431
rect 29089 2391 29147 2397
rect 29822 2388 29828 2440
rect 29880 2388 29886 2440
rect 30282 2388 30288 2440
rect 30340 2428 30346 2440
rect 30561 2431 30619 2437
rect 30561 2428 30573 2431
rect 30340 2400 30573 2428
rect 30340 2388 30346 2400
rect 30561 2397 30573 2400
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 31478 2388 31484 2440
rect 31536 2388 31542 2440
rect 32030 2388 32036 2440
rect 32088 2428 32094 2440
rect 32088 2400 32444 2428
rect 32088 2388 32094 2400
rect 1762 2320 1768 2372
rect 1820 2320 1826 2372
rect 3418 2320 3424 2372
rect 3476 2320 3482 2372
rect 3602 2320 3608 2372
rect 3660 2320 3666 2372
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 16816 2332 23796 2360
rect 16816 2320 16822 2332
rect 7926 2252 7932 2304
rect 7984 2252 7990 2304
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 9214 2252 9220 2304
rect 9272 2252 9278 2304
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17865 2295 17923 2301
rect 17865 2292 17877 2295
rect 17000 2264 17877 2292
rect 17000 2252 17006 2264
rect 17865 2261 17877 2264
rect 17911 2261 17923 2295
rect 17865 2255 17923 2261
rect 20070 2252 20076 2304
rect 20128 2252 20134 2304
rect 20806 2252 20812 2304
rect 20864 2252 20870 2304
rect 21818 2252 21824 2304
rect 21876 2252 21882 2304
rect 23768 2301 23796 2332
rect 31110 2320 31116 2372
rect 31168 2320 31174 2372
rect 32122 2320 32128 2372
rect 32180 2320 32186 2372
rect 32416 2360 32444 2400
rect 32490 2388 32496 2440
rect 32548 2388 32554 2440
rect 32950 2388 32956 2440
rect 33008 2428 33014 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 33008 2400 33425 2428
rect 33008 2388 33014 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 33502 2388 33508 2440
rect 33560 2428 33566 2440
rect 34149 2431 34207 2437
rect 34149 2428 34161 2431
rect 33560 2400 34161 2428
rect 33560 2388 33566 2400
rect 34149 2397 34161 2400
rect 34195 2397 34207 2431
rect 34149 2391 34207 2397
rect 34238 2388 34244 2440
rect 34296 2388 34302 2440
rect 34330 2388 34336 2440
rect 34388 2388 34394 2440
rect 34514 2388 34520 2440
rect 34572 2428 34578 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34572 2400 34897 2428
rect 34572 2388 34578 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36136 2400 36369 2428
rect 36136 2388 36142 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 37274 2388 37280 2440
rect 37332 2428 37338 2440
rect 37936 2437 37964 2468
rect 37369 2431 37427 2437
rect 37369 2428 37381 2431
rect 37332 2400 37381 2428
rect 37332 2388 37338 2400
rect 37369 2397 37381 2400
rect 37415 2397 37427 2431
rect 37369 2391 37427 2397
rect 37921 2431 37979 2437
rect 37921 2397 37933 2431
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 32769 2363 32827 2369
rect 32769 2360 32781 2363
rect 32416 2332 32781 2360
rect 32769 2329 32781 2332
rect 32815 2329 32827 2363
rect 34348 2360 34376 2388
rect 35621 2363 35679 2369
rect 35621 2360 35633 2363
rect 34348 2332 35633 2360
rect 32769 2323 32827 2329
rect 35621 2329 35633 2332
rect 35667 2329 35679 2363
rect 38028 2360 38056 2536
rect 38580 2437 38608 2604
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 39301 2431 39359 2437
rect 39301 2397 39313 2431
rect 39347 2397 39359 2431
rect 39301 2391 39359 2397
rect 39316 2360 39344 2391
rect 39666 2388 39672 2440
rect 39724 2428 39730 2440
rect 40037 2431 40095 2437
rect 40037 2428 40049 2431
rect 39724 2400 40049 2428
rect 39724 2388 39730 2400
rect 40037 2397 40049 2400
rect 40083 2397 40095 2431
rect 40037 2391 40095 2397
rect 40402 2388 40408 2440
rect 40460 2428 40466 2440
rect 40773 2431 40831 2437
rect 40773 2428 40785 2431
rect 40460 2400 40785 2428
rect 40460 2388 40466 2400
rect 40773 2397 40785 2400
rect 40819 2397 40831 2431
rect 40773 2391 40831 2397
rect 41414 2388 41420 2440
rect 41472 2428 41478 2440
rect 41509 2431 41567 2437
rect 41509 2428 41521 2431
rect 41472 2400 41521 2428
rect 41472 2388 41478 2400
rect 41509 2397 41521 2400
rect 41555 2397 41567 2431
rect 41509 2391 41567 2397
rect 41690 2388 41696 2440
rect 41748 2428 41754 2440
rect 42521 2431 42579 2437
rect 42521 2428 42533 2431
rect 41748 2400 42533 2428
rect 41748 2388 41754 2400
rect 42521 2397 42533 2400
rect 42567 2397 42579 2431
rect 42521 2391 42579 2397
rect 42702 2388 42708 2440
rect 42760 2428 42766 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 42760 2400 43085 2428
rect 42760 2388 42766 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 43162 2388 43168 2440
rect 43220 2428 43226 2440
rect 43717 2431 43775 2437
rect 43717 2428 43729 2431
rect 43220 2400 43729 2428
rect 43220 2388 43226 2400
rect 43717 2397 43729 2400
rect 43763 2397 43775 2431
rect 43717 2391 43775 2397
rect 38028 2332 39344 2360
rect 35621 2323 35679 2329
rect 23753 2295 23811 2301
rect 23753 2261 23765 2295
rect 23799 2261 23811 2295
rect 23753 2255 23811 2261
rect 24486 2252 24492 2304
rect 24544 2252 24550 2304
rect 32490 2252 32496 2304
rect 32548 2292 32554 2304
rect 32861 2295 32919 2301
rect 32861 2292 32873 2295
rect 32548 2264 32873 2292
rect 32548 2252 32554 2264
rect 32861 2261 32873 2264
rect 32907 2261 32919 2295
rect 32861 2255 32919 2261
rect 33502 2252 33508 2304
rect 33560 2252 33566 2304
rect 34238 2252 34244 2304
rect 34296 2252 34302 2304
rect 34974 2252 34980 2304
rect 35032 2252 35038 2304
rect 35894 2252 35900 2304
rect 35952 2252 35958 2304
rect 36446 2252 36452 2304
rect 36504 2252 36510 2304
rect 37182 2252 37188 2304
rect 37240 2292 37246 2304
rect 37461 2295 37519 2301
rect 37461 2292 37473 2295
rect 37240 2264 37473 2292
rect 37240 2252 37246 2264
rect 37461 2261 37473 2264
rect 37507 2261 37519 2295
rect 37461 2255 37519 2261
rect 38010 2252 38016 2304
rect 38068 2252 38074 2304
rect 38378 2252 38384 2304
rect 38436 2292 38442 2304
rect 38657 2295 38715 2301
rect 38657 2292 38669 2295
rect 38436 2264 38669 2292
rect 38436 2252 38442 2264
rect 38657 2261 38669 2264
rect 38703 2261 38715 2295
rect 38657 2255 38715 2261
rect 39390 2252 39396 2304
rect 39448 2252 39454 2304
rect 39850 2252 39856 2304
rect 39908 2292 39914 2304
rect 40129 2295 40187 2301
rect 40129 2292 40141 2295
rect 39908 2264 40141 2292
rect 39908 2252 39914 2264
rect 40129 2261 40141 2264
rect 40175 2261 40187 2295
rect 40129 2255 40187 2261
rect 40862 2252 40868 2304
rect 40920 2252 40926 2304
rect 41322 2252 41328 2304
rect 41380 2292 41386 2304
rect 41601 2295 41659 2301
rect 41601 2292 41613 2295
rect 41380 2264 41613 2292
rect 41380 2252 41386 2264
rect 41601 2261 41613 2264
rect 41647 2261 41659 2295
rect 41601 2255 41659 2261
rect 42426 2252 42432 2304
rect 42484 2292 42490 2304
rect 42797 2295 42855 2301
rect 42797 2292 42809 2295
rect 42484 2264 42809 2292
rect 42484 2252 42490 2264
rect 42797 2261 42809 2264
rect 42843 2261 42855 2295
rect 42797 2255 42855 2261
rect 43162 2252 43168 2304
rect 43220 2252 43226 2304
rect 43806 2252 43812 2304
rect 43864 2252 43870 2304
rect 1104 2202 45051 2224
rect 1104 2150 11896 2202
rect 11948 2150 11960 2202
rect 12012 2150 12024 2202
rect 12076 2150 12088 2202
rect 12140 2150 12152 2202
rect 12204 2150 22843 2202
rect 22895 2150 22907 2202
rect 22959 2150 22971 2202
rect 23023 2150 23035 2202
rect 23087 2150 23099 2202
rect 23151 2150 33790 2202
rect 33842 2150 33854 2202
rect 33906 2150 33918 2202
rect 33970 2150 33982 2202
rect 34034 2150 34046 2202
rect 34098 2150 44737 2202
rect 44789 2150 44801 2202
rect 44853 2150 44865 2202
rect 44917 2150 44929 2202
rect 44981 2150 44993 2202
rect 45045 2150 45051 2202
rect 1104 2128 45051 2150
rect 7926 2048 7932 2100
rect 7984 2048 7990 2100
rect 15378 2048 15384 2100
rect 15436 2088 15442 2100
rect 20070 2088 20076 2100
rect 15436 2060 20076 2088
rect 15436 2048 15442 2060
rect 20070 2048 20076 2060
rect 20128 2048 20134 2100
rect 20272 2060 24072 2088
rect 7944 2020 7972 2048
rect 20272 2020 20300 2060
rect 24044 2032 24072 2060
rect 7944 1992 20300 2020
rect 24026 1980 24032 2032
rect 24084 1980 24090 2032
rect 15746 1912 15752 1964
rect 15804 1952 15810 1964
rect 21818 1952 21824 1964
rect 15804 1924 21824 1952
rect 15804 1912 15810 1924
rect 21818 1912 21824 1924
rect 21876 1912 21882 1964
rect 12802 1844 12808 1896
rect 12860 1884 12866 1896
rect 20806 1884 20812 1896
rect 12860 1856 20812 1884
rect 12860 1844 12866 1856
rect 20806 1844 20812 1856
rect 20864 1844 20870 1896
rect 16850 1776 16856 1828
rect 16908 1816 16914 1828
rect 24486 1816 24492 1828
rect 16908 1788 24492 1816
rect 16908 1776 16914 1788
rect 24486 1776 24492 1788
rect 24544 1776 24550 1828
rect 1670 1300 1676 1352
rect 1728 1340 1734 1352
rect 33594 1340 33600 1352
rect 1728 1312 33600 1340
rect 1728 1300 1734 1312
rect 33594 1300 33600 1312
rect 33652 1300 33658 1352
rect 3602 1232 3608 1284
rect 3660 1272 3666 1284
rect 34790 1272 34796 1284
rect 3660 1244 34796 1272
rect 3660 1232 3666 1244
rect 34790 1232 34796 1244
rect 34848 1232 34854 1284
rect 5626 1164 5632 1216
rect 5684 1204 5690 1216
rect 35710 1204 35716 1216
rect 5684 1176 35716 1204
rect 5684 1164 5690 1176
rect 35710 1164 35716 1176
rect 35768 1164 35774 1216
<< via1 >>
rect 28080 6536 28132 6588
rect 28540 6536 28592 6588
rect 5908 6468 5960 6520
rect 19984 6468 20036 6520
rect 9496 6400 9548 6452
rect 23572 6400 23624 6452
rect 7656 6332 7708 6384
rect 25228 6332 25280 6384
rect 4160 6264 4212 6316
rect 35164 6264 35216 6316
rect 1952 6196 2004 6248
rect 33232 6196 33284 6248
rect 2688 6128 2740 6180
rect 35072 6128 35124 6180
rect 13636 6060 13688 6112
rect 29000 6060 29052 6112
rect 8116 5992 8168 6044
rect 24124 5992 24176 6044
rect 8024 5924 8076 5976
rect 25136 5924 25188 5976
rect 16396 5856 16448 5908
rect 40316 5856 40368 5908
rect 15752 5788 15804 5840
rect 40592 5788 40644 5840
rect 12624 5720 12676 5772
rect 38660 5720 38712 5772
rect 9404 5652 9456 5704
rect 22192 5652 22244 5704
rect 7748 5584 7800 5636
rect 23848 5584 23900 5636
rect 14924 5516 14976 5568
rect 25412 5516 25464 5568
rect 11896 5414 11948 5466
rect 11960 5414 12012 5466
rect 12024 5414 12076 5466
rect 12088 5414 12140 5466
rect 12152 5414 12204 5466
rect 22843 5414 22895 5466
rect 22907 5414 22959 5466
rect 22971 5414 23023 5466
rect 23035 5414 23087 5466
rect 23099 5414 23151 5466
rect 33790 5414 33842 5466
rect 33854 5414 33906 5466
rect 33918 5414 33970 5466
rect 33982 5414 34034 5466
rect 34046 5414 34098 5466
rect 44737 5414 44789 5466
rect 44801 5414 44853 5466
rect 44865 5414 44917 5466
rect 44929 5414 44981 5466
rect 44993 5414 45045 5466
rect 6000 5312 6052 5364
rect 7380 5312 7432 5364
rect 7932 5312 7984 5364
rect 8484 5312 8536 5364
rect 9036 5312 9088 5364
rect 10140 5312 10192 5364
rect 11244 5312 11296 5364
rect 12532 5312 12584 5364
rect 13176 5312 13228 5364
rect 14280 5312 14332 5364
rect 15108 5312 15160 5364
rect 15660 5312 15712 5364
rect 16212 5312 16264 5364
rect 16764 5312 16816 5364
rect 17592 5312 17644 5364
rect 18144 5312 18196 5364
rect 18696 5312 18748 5364
rect 18880 5355 18932 5364
rect 18880 5321 18889 5355
rect 18889 5321 18923 5355
rect 18923 5321 18932 5355
rect 18880 5312 18932 5321
rect 7748 5244 7800 5296
rect 9404 5244 9456 5296
rect 6092 5219 6144 5228
rect 6092 5185 6101 5219
rect 6101 5185 6135 5219
rect 6135 5185 6144 5219
rect 6092 5176 6144 5185
rect 6736 5176 6788 5228
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 6552 5108 6604 5160
rect 10508 5176 10560 5228
rect 11152 5176 11204 5228
rect 11336 5176 11388 5228
rect 11612 5176 11664 5228
rect 13636 5244 13688 5296
rect 13084 5176 13136 5228
rect 13176 5176 13228 5228
rect 16948 5244 17000 5296
rect 17132 5244 17184 5296
rect 19248 5244 19300 5296
rect 19524 5312 19576 5364
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 15200 5176 15252 5228
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 11244 4972 11296 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 11888 4972 11940 5024
rect 13268 5040 13320 5092
rect 17776 5176 17828 5228
rect 17960 5176 18012 5228
rect 18880 5176 18932 5228
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 19708 5219 19760 5228
rect 19708 5185 19717 5219
rect 19717 5185 19751 5219
rect 19751 5185 19760 5219
rect 19708 5176 19760 5185
rect 19892 5287 19944 5296
rect 19892 5253 19901 5287
rect 19901 5253 19935 5287
rect 19935 5253 19944 5287
rect 19892 5244 19944 5253
rect 20168 5176 20220 5228
rect 21916 5312 21968 5364
rect 24768 5312 24820 5364
rect 24952 5244 25004 5296
rect 25320 5244 25372 5296
rect 21364 5219 21416 5228
rect 21364 5185 21373 5219
rect 21373 5185 21407 5219
rect 21407 5185 21416 5219
rect 21364 5176 21416 5185
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 21732 5176 21784 5228
rect 22100 5176 22152 5228
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 23112 5219 23164 5228
rect 23112 5185 23121 5219
rect 23121 5185 23155 5219
rect 23155 5185 23164 5219
rect 23112 5176 23164 5185
rect 23388 5219 23440 5228
rect 23388 5185 23397 5219
rect 23397 5185 23431 5219
rect 23431 5185 23440 5219
rect 23388 5176 23440 5185
rect 23480 5176 23532 5228
rect 23756 5176 23808 5228
rect 24032 5176 24084 5228
rect 24308 5176 24360 5228
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 25872 5244 25924 5296
rect 27620 5312 27672 5364
rect 26976 5244 27028 5296
rect 18328 5108 18380 5160
rect 23020 5108 23072 5160
rect 25044 5108 25096 5160
rect 25780 5219 25832 5228
rect 25780 5185 25789 5219
rect 25789 5185 25823 5219
rect 25823 5185 25832 5219
rect 25780 5176 25832 5185
rect 26056 5219 26108 5228
rect 26056 5185 26065 5219
rect 26065 5185 26099 5219
rect 26099 5185 26108 5219
rect 26056 5176 26108 5185
rect 26332 5219 26384 5228
rect 26332 5185 26341 5219
rect 26341 5185 26375 5219
rect 26375 5185 26384 5219
rect 26332 5176 26384 5185
rect 26608 5219 26660 5228
rect 26608 5185 26617 5219
rect 26617 5185 26651 5219
rect 26651 5185 26660 5219
rect 26608 5176 26660 5185
rect 26700 5176 26752 5228
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 34520 5312 34572 5364
rect 34612 5312 34664 5364
rect 34980 5312 35032 5364
rect 35532 5312 35584 5364
rect 36544 5312 36596 5364
rect 38200 5312 38252 5364
rect 39672 5312 39724 5364
rect 28356 5244 28408 5296
rect 27804 5108 27856 5160
rect 28540 5219 28592 5228
rect 28540 5185 28549 5219
rect 28549 5185 28583 5219
rect 28583 5185 28592 5219
rect 28540 5176 28592 5185
rect 28724 5244 28776 5296
rect 30104 5219 30156 5228
rect 30104 5185 30113 5219
rect 30113 5185 30147 5219
rect 30147 5185 30156 5219
rect 30104 5176 30156 5185
rect 30380 5219 30432 5228
rect 30380 5185 30389 5219
rect 30389 5185 30423 5219
rect 30423 5185 30432 5219
rect 30380 5176 30432 5185
rect 30656 5219 30708 5228
rect 30656 5185 30665 5219
rect 30665 5185 30699 5219
rect 30699 5185 30708 5219
rect 30656 5176 30708 5185
rect 30932 5219 30984 5228
rect 30932 5185 30941 5219
rect 30941 5185 30975 5219
rect 30975 5185 30984 5219
rect 30932 5176 30984 5185
rect 31208 5219 31260 5228
rect 31208 5185 31217 5219
rect 31217 5185 31251 5219
rect 31251 5185 31260 5219
rect 31208 5176 31260 5185
rect 31484 5219 31536 5228
rect 31484 5185 31493 5219
rect 31493 5185 31527 5219
rect 31527 5185 31536 5219
rect 31484 5176 31536 5185
rect 31760 5219 31812 5228
rect 31760 5185 31769 5219
rect 31769 5185 31803 5219
rect 31803 5185 31812 5219
rect 31760 5176 31812 5185
rect 32128 5219 32180 5228
rect 32128 5185 32137 5219
rect 32137 5185 32171 5219
rect 32171 5185 32180 5219
rect 32128 5176 32180 5185
rect 32404 5219 32456 5228
rect 32404 5185 32413 5219
rect 32413 5185 32447 5219
rect 32447 5185 32456 5219
rect 32404 5176 32456 5185
rect 32680 5219 32732 5228
rect 32680 5185 32689 5219
rect 32689 5185 32723 5219
rect 32723 5185 32732 5219
rect 32680 5176 32732 5185
rect 32956 5219 33008 5228
rect 32956 5185 32965 5219
rect 32965 5185 32999 5219
rect 32999 5185 33008 5219
rect 32956 5176 33008 5185
rect 33048 5176 33100 5228
rect 33508 5219 33560 5228
rect 33508 5185 33517 5219
rect 33517 5185 33551 5219
rect 33551 5185 33560 5219
rect 33508 5176 33560 5185
rect 33784 5219 33836 5228
rect 33784 5185 33793 5219
rect 33793 5185 33827 5219
rect 33827 5185 33836 5219
rect 33784 5176 33836 5185
rect 34244 5219 34296 5228
rect 34244 5185 34253 5219
rect 34253 5185 34287 5219
rect 34287 5185 34296 5219
rect 34244 5176 34296 5185
rect 34336 5176 34388 5228
rect 34612 5176 34664 5228
rect 35348 5219 35400 5228
rect 35348 5185 35357 5219
rect 35357 5185 35391 5219
rect 35391 5185 35400 5219
rect 35348 5176 35400 5185
rect 22008 5040 22060 5092
rect 27988 5040 28040 5092
rect 31852 5040 31904 5092
rect 32496 5040 32548 5092
rect 33048 5040 33100 5092
rect 33140 5083 33192 5092
rect 33140 5049 33149 5083
rect 33149 5049 33183 5083
rect 33183 5049 33192 5083
rect 33140 5040 33192 5049
rect 33324 5040 33376 5092
rect 35256 5108 35308 5160
rect 35532 5108 35584 5160
rect 34428 5040 34480 5092
rect 36728 5176 36780 5228
rect 38660 5244 38712 5296
rect 40040 5244 40092 5296
rect 37188 5108 37240 5160
rect 38016 5108 38068 5160
rect 40500 5219 40552 5228
rect 40500 5185 40509 5219
rect 40509 5185 40543 5219
rect 40543 5185 40552 5219
rect 40500 5176 40552 5185
rect 40592 5176 40644 5228
rect 37648 5040 37700 5092
rect 12808 4972 12860 5024
rect 13728 4972 13780 5024
rect 13820 4972 13872 5024
rect 20536 4972 20588 5024
rect 20720 4972 20772 5024
rect 21272 4972 21324 5024
rect 21824 5015 21876 5024
rect 21824 4981 21833 5015
rect 21833 4981 21867 5015
rect 21867 4981 21876 5015
rect 21824 4972 21876 4981
rect 22100 5015 22152 5024
rect 22100 4981 22109 5015
rect 22109 4981 22143 5015
rect 22143 4981 22152 5015
rect 22100 4972 22152 4981
rect 22192 4972 22244 5024
rect 22376 5015 22428 5024
rect 22376 4981 22385 5015
rect 22385 4981 22419 5015
rect 22419 4981 22428 5015
rect 22376 4972 22428 4981
rect 22652 5015 22704 5024
rect 22652 4981 22661 5015
rect 22661 4981 22695 5015
rect 22695 4981 22704 5015
rect 22652 4972 22704 4981
rect 22928 5015 22980 5024
rect 22928 4981 22937 5015
rect 22937 4981 22971 5015
rect 22971 4981 22980 5015
rect 22928 4972 22980 4981
rect 23204 5015 23256 5024
rect 23204 4981 23213 5015
rect 23213 4981 23247 5015
rect 23247 4981 23256 5015
rect 23204 4972 23256 4981
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 23756 5015 23808 5024
rect 23756 4981 23765 5015
rect 23765 4981 23799 5015
rect 23799 4981 23808 5015
rect 23756 4972 23808 4981
rect 24032 5015 24084 5024
rect 24032 4981 24041 5015
rect 24041 4981 24075 5015
rect 24075 4981 24084 5015
rect 24032 4972 24084 4981
rect 24400 5015 24452 5024
rect 24400 4981 24409 5015
rect 24409 4981 24443 5015
rect 24443 4981 24452 5015
rect 24400 4972 24452 4981
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 24952 5015 25004 5024
rect 24952 4981 24961 5015
rect 24961 4981 24995 5015
rect 24995 4981 25004 5015
rect 24952 4972 25004 4981
rect 25228 5015 25280 5024
rect 25228 4981 25237 5015
rect 25237 4981 25271 5015
rect 25271 4981 25280 5015
rect 25228 4972 25280 4981
rect 25504 5015 25556 5024
rect 25504 4981 25513 5015
rect 25513 4981 25547 5015
rect 25547 4981 25556 5015
rect 25504 4972 25556 4981
rect 25964 5015 26016 5024
rect 25964 4981 25973 5015
rect 25973 4981 26007 5015
rect 26007 4981 26016 5015
rect 25964 4972 26016 4981
rect 26240 5015 26292 5024
rect 26240 4981 26249 5015
rect 26249 4981 26283 5015
rect 26283 4981 26292 5015
rect 26240 4972 26292 4981
rect 26516 5015 26568 5024
rect 26516 4981 26525 5015
rect 26525 4981 26559 5015
rect 26559 4981 26568 5015
rect 26516 4972 26568 4981
rect 26700 4972 26752 5024
rect 26976 5015 27028 5024
rect 26976 4981 26985 5015
rect 26985 4981 27019 5015
rect 27019 4981 27028 5015
rect 26976 4972 27028 4981
rect 27252 5015 27304 5024
rect 27252 4981 27261 5015
rect 27261 4981 27295 5015
rect 27295 4981 27304 5015
rect 27252 4972 27304 4981
rect 27804 5015 27856 5024
rect 27804 4981 27813 5015
rect 27813 4981 27847 5015
rect 27847 4981 27856 5015
rect 27804 4972 27856 4981
rect 27896 4972 27948 5024
rect 28264 4972 28316 5024
rect 28724 4972 28776 5024
rect 28908 5015 28960 5024
rect 28908 4981 28917 5015
rect 28917 4981 28951 5015
rect 28951 4981 28960 5015
rect 28908 4972 28960 4981
rect 30472 4972 30524 5024
rect 30564 5015 30616 5024
rect 30564 4981 30573 5015
rect 30573 4981 30607 5015
rect 30607 4981 30616 5015
rect 30564 4972 30616 4981
rect 30840 5015 30892 5024
rect 30840 4981 30849 5015
rect 30849 4981 30883 5015
rect 30883 4981 30892 5015
rect 30840 4972 30892 4981
rect 31116 5015 31168 5024
rect 31116 4981 31125 5015
rect 31125 4981 31159 5015
rect 31159 4981 31168 5015
rect 31116 4972 31168 4981
rect 31760 4972 31812 5024
rect 31944 5015 31996 5024
rect 31944 4981 31953 5015
rect 31953 4981 31987 5015
rect 31987 4981 31996 5015
rect 31944 4972 31996 4981
rect 32312 5015 32364 5024
rect 32312 4981 32321 5015
rect 32321 4981 32355 5015
rect 32355 4981 32364 5015
rect 32312 4972 32364 4981
rect 33416 5015 33468 5024
rect 33416 4981 33425 5015
rect 33425 4981 33459 5015
rect 33459 4981 33468 5015
rect 33416 4972 33468 4981
rect 33692 5015 33744 5024
rect 33692 4981 33701 5015
rect 33701 4981 33735 5015
rect 33735 4981 33744 5015
rect 33692 4972 33744 4981
rect 34152 4972 34204 5024
rect 35716 4972 35768 5024
rect 36912 4972 36964 5024
rect 39304 4972 39356 5024
rect 6423 4870 6475 4922
rect 6487 4870 6539 4922
rect 6551 4870 6603 4922
rect 6615 4870 6667 4922
rect 6679 4870 6731 4922
rect 17370 4870 17422 4922
rect 17434 4870 17486 4922
rect 17498 4870 17550 4922
rect 17562 4870 17614 4922
rect 17626 4870 17678 4922
rect 28317 4870 28369 4922
rect 28381 4870 28433 4922
rect 28445 4870 28497 4922
rect 28509 4870 28561 4922
rect 28573 4870 28625 4922
rect 39264 4870 39316 4922
rect 39328 4870 39380 4922
rect 39392 4870 39444 4922
rect 39456 4870 39508 4922
rect 39520 4870 39572 4922
rect 6092 4768 6144 4820
rect 5724 4743 5776 4752
rect 5724 4709 5733 4743
rect 5733 4709 5767 4743
rect 5767 4709 5776 4743
rect 5724 4700 5776 4709
rect 6276 4743 6328 4752
rect 6276 4709 6285 4743
rect 6285 4709 6319 4743
rect 6319 4709 6328 4743
rect 6276 4700 6328 4709
rect 6828 4743 6880 4752
rect 6828 4709 6837 4743
rect 6837 4709 6871 4743
rect 6871 4709 6880 4743
rect 6828 4700 6880 4709
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 9312 4811 9364 4820
rect 9312 4777 9321 4811
rect 9321 4777 9355 4811
rect 9355 4777 9364 4811
rect 9312 4768 9364 4777
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10416 4811 10468 4820
rect 10416 4777 10425 4811
rect 10425 4777 10459 4811
rect 10459 4777 10468 4811
rect 10416 4768 10468 4777
rect 11060 4811 11112 4820
rect 11060 4777 11069 4811
rect 11069 4777 11103 4811
rect 11103 4777 11112 4811
rect 11060 4768 11112 4777
rect 11428 4811 11480 4820
rect 11428 4777 11437 4811
rect 11437 4777 11471 4811
rect 11471 4777 11480 4811
rect 11428 4768 11480 4777
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14188 4811 14240 4820
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 11704 4700 11756 4752
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 6184 4564 6236 4616
rect 8024 4564 8076 4616
rect 8116 4607 8168 4616
rect 8116 4573 8125 4607
rect 8125 4573 8159 4607
rect 8159 4573 8168 4607
rect 8116 4564 8168 4573
rect 9496 4564 9548 4616
rect 7656 4496 7708 4548
rect 9404 4539 9456 4548
rect 9404 4505 9413 4539
rect 9413 4505 9447 4539
rect 9447 4505 9456 4539
rect 9404 4496 9456 4505
rect 10784 4539 10836 4548
rect 10784 4505 10793 4539
rect 10793 4505 10827 4539
rect 10827 4505 10836 4539
rect 10784 4496 10836 4505
rect 11428 4564 11480 4616
rect 14832 4743 14884 4752
rect 14832 4709 14841 4743
rect 14841 4709 14875 4743
rect 14875 4709 14884 4743
rect 14832 4700 14884 4709
rect 15384 4743 15436 4752
rect 15384 4709 15393 4743
rect 15393 4709 15427 4743
rect 15427 4709 15436 4743
rect 15384 4700 15436 4709
rect 15936 4811 15988 4820
rect 15936 4777 15945 4811
rect 15945 4777 15979 4811
rect 15979 4777 15988 4811
rect 15936 4768 15988 4777
rect 16028 4768 16080 4820
rect 15108 4632 15160 4684
rect 15660 4632 15712 4684
rect 16488 4743 16540 4752
rect 16488 4709 16497 4743
rect 16497 4709 16531 4743
rect 16531 4709 16540 4743
rect 16488 4700 16540 4709
rect 17040 4743 17092 4752
rect 17040 4709 17049 4743
rect 17049 4709 17083 4743
rect 17083 4709 17092 4743
rect 17040 4700 17092 4709
rect 17316 4768 17368 4820
rect 17868 4768 17920 4820
rect 18420 4768 18472 4820
rect 18788 4768 18840 4820
rect 19800 4768 19852 4820
rect 14924 4564 14976 4616
rect 15384 4564 15436 4616
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 17132 4632 17184 4684
rect 19340 4743 19392 4752
rect 19340 4709 19349 4743
rect 19349 4709 19383 4743
rect 19383 4709 19392 4743
rect 19340 4700 19392 4709
rect 19892 4700 19944 4752
rect 20444 4768 20496 4820
rect 12256 4496 12308 4548
rect 12716 4539 12768 4548
rect 12716 4505 12725 4539
rect 12725 4505 12759 4539
rect 12759 4505 12768 4539
rect 12716 4496 12768 4505
rect 13268 4539 13320 4548
rect 13268 4505 13277 4539
rect 13277 4505 13311 4539
rect 13311 4505 13320 4539
rect 13268 4496 13320 4505
rect 13360 4496 13412 4548
rect 16672 4539 16724 4548
rect 16672 4505 16681 4539
rect 16681 4505 16715 4539
rect 16715 4505 16724 4539
rect 16672 4496 16724 4505
rect 17224 4539 17276 4548
rect 17224 4505 17233 4539
rect 17233 4505 17267 4539
rect 17267 4505 17276 4539
rect 17224 4496 17276 4505
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 18328 4564 18380 4616
rect 20260 4632 20312 4684
rect 22100 4768 22152 4820
rect 22652 4768 22704 4820
rect 21456 4700 21508 4752
rect 18604 4539 18656 4548
rect 18604 4505 18613 4539
rect 18613 4505 18647 4539
rect 18647 4505 18656 4539
rect 18604 4496 18656 4505
rect 18788 4496 18840 4548
rect 19616 4564 19668 4616
rect 19524 4428 19576 4480
rect 19892 4471 19944 4480
rect 19892 4437 19901 4471
rect 19901 4437 19935 4471
rect 19935 4437 19944 4471
rect 19892 4428 19944 4437
rect 20076 4607 20128 4616
rect 20076 4573 20077 4607
rect 20077 4573 20111 4607
rect 20111 4573 20128 4607
rect 20076 4564 20128 4573
rect 20352 4607 20404 4616
rect 20352 4573 20361 4607
rect 20361 4573 20395 4607
rect 20395 4573 20404 4607
rect 20352 4564 20404 4573
rect 20536 4564 20588 4616
rect 20628 4607 20680 4616
rect 20628 4573 20637 4607
rect 20637 4573 20671 4607
rect 20671 4573 20680 4607
rect 20628 4564 20680 4573
rect 20812 4496 20864 4548
rect 21364 4564 21416 4616
rect 21824 4632 21876 4684
rect 22376 4564 22428 4616
rect 22928 4768 22980 4820
rect 23204 4768 23256 4820
rect 23480 4768 23532 4820
rect 23756 4768 23808 4820
rect 23572 4564 23624 4616
rect 24032 4768 24084 4820
rect 24400 4768 24452 4820
rect 24676 4768 24728 4820
rect 24860 4768 24912 4820
rect 25964 4768 26016 4820
rect 27620 4811 27672 4820
rect 27620 4777 27629 4811
rect 27629 4777 27663 4811
rect 27663 4777 27672 4811
rect 27620 4768 27672 4777
rect 24492 4564 24544 4616
rect 24952 4700 25004 4752
rect 25228 4700 25280 4752
rect 25504 4700 25556 4752
rect 26332 4743 26384 4752
rect 26332 4709 26341 4743
rect 26341 4709 26375 4743
rect 26375 4709 26384 4743
rect 26332 4700 26384 4709
rect 26240 4632 26292 4684
rect 20076 4428 20128 4480
rect 20260 4428 20312 4480
rect 20904 4428 20956 4480
rect 21088 4428 21140 4480
rect 22284 4471 22336 4480
rect 22284 4437 22293 4471
rect 22293 4437 22327 4471
rect 22327 4437 22336 4471
rect 22284 4428 22336 4437
rect 22468 4428 22520 4480
rect 22652 4471 22704 4480
rect 22652 4437 22661 4471
rect 22661 4437 22695 4471
rect 22695 4437 22704 4471
rect 22652 4428 22704 4437
rect 22744 4428 22796 4480
rect 24124 4496 24176 4548
rect 23848 4471 23900 4480
rect 23848 4437 23857 4471
rect 23857 4437 23891 4471
rect 23891 4437 23900 4471
rect 23848 4428 23900 4437
rect 25044 4496 25096 4548
rect 28172 4768 28224 4820
rect 28448 4811 28500 4820
rect 28448 4777 28457 4811
rect 28457 4777 28491 4811
rect 28491 4777 28500 4811
rect 28448 4768 28500 4777
rect 28724 4768 28776 4820
rect 28908 4768 28960 4820
rect 29000 4811 29052 4820
rect 29000 4777 29009 4811
rect 29009 4777 29043 4811
rect 29043 4777 29052 4811
rect 29000 4768 29052 4777
rect 30564 4768 30616 4820
rect 30840 4768 30892 4820
rect 31116 4768 31168 4820
rect 33508 4768 33560 4820
rect 34428 4811 34480 4820
rect 34428 4777 34437 4811
rect 34437 4777 34471 4811
rect 34471 4777 34480 4811
rect 34428 4768 34480 4777
rect 34796 4811 34848 4820
rect 34796 4777 34805 4811
rect 34805 4777 34839 4811
rect 34839 4777 34848 4811
rect 34796 4768 34848 4777
rect 35256 4811 35308 4820
rect 35256 4777 35265 4811
rect 35265 4777 35299 4811
rect 35299 4777 35308 4811
rect 35256 4768 35308 4777
rect 35348 4768 35400 4820
rect 35808 4768 35860 4820
rect 36636 4768 36688 4820
rect 37740 4768 37792 4820
rect 38384 4768 38436 4820
rect 28908 4564 28960 4616
rect 29184 4607 29236 4616
rect 29184 4573 29193 4607
rect 29193 4573 29227 4607
rect 29227 4573 29236 4607
rect 29184 4564 29236 4573
rect 29920 4607 29972 4616
rect 29920 4573 29929 4607
rect 29929 4573 29963 4607
rect 29963 4573 29972 4607
rect 29920 4564 29972 4573
rect 31760 4700 31812 4752
rect 31852 4700 31904 4752
rect 32036 4743 32088 4752
rect 32036 4709 32045 4743
rect 32045 4709 32079 4743
rect 32079 4709 32088 4743
rect 32036 4700 32088 4709
rect 36176 4700 36228 4752
rect 37280 4700 37332 4752
rect 38568 4700 38620 4752
rect 39672 4768 39724 4820
rect 40224 4768 40276 4820
rect 39948 4700 40000 4752
rect 24952 4471 25004 4480
rect 24952 4437 24961 4471
rect 24961 4437 24995 4471
rect 24995 4437 25004 4471
rect 24952 4428 25004 4437
rect 25136 4428 25188 4480
rect 25504 4471 25556 4480
rect 25504 4437 25513 4471
rect 25513 4437 25547 4471
rect 25547 4437 25556 4471
rect 25504 4428 25556 4437
rect 27988 4496 28040 4548
rect 28080 4428 28132 4480
rect 29736 4471 29788 4480
rect 29736 4437 29745 4471
rect 29745 4437 29779 4471
rect 29779 4437 29788 4471
rect 29736 4428 29788 4437
rect 31024 4471 31076 4480
rect 31024 4437 31033 4471
rect 31033 4437 31067 4471
rect 31067 4437 31076 4471
rect 31024 4428 31076 4437
rect 31392 4471 31444 4480
rect 31392 4437 31401 4471
rect 31401 4437 31435 4471
rect 31435 4437 31444 4471
rect 31392 4428 31444 4437
rect 33232 4564 33284 4616
rect 34428 4564 34480 4616
rect 35072 4607 35124 4616
rect 35072 4573 35081 4607
rect 35081 4573 35115 4607
rect 35115 4573 35124 4607
rect 35072 4564 35124 4573
rect 35164 4564 35216 4616
rect 35624 4607 35676 4616
rect 35624 4573 35633 4607
rect 35633 4573 35667 4607
rect 35667 4573 35676 4607
rect 35624 4564 35676 4573
rect 40132 4632 40184 4684
rect 40316 4564 40368 4616
rect 41512 4607 41564 4616
rect 41512 4573 41521 4607
rect 41521 4573 41555 4607
rect 41555 4573 41564 4607
rect 41512 4564 41564 4573
rect 32956 4428 33008 4480
rect 37096 4539 37148 4548
rect 37096 4505 37105 4539
rect 37105 4505 37139 4539
rect 37139 4505 37148 4539
rect 37096 4496 37148 4505
rect 37648 4539 37700 4548
rect 37648 4505 37657 4539
rect 37657 4505 37691 4539
rect 37691 4505 37700 4539
rect 37648 4496 37700 4505
rect 37740 4496 37792 4548
rect 39304 4539 39356 4548
rect 39304 4505 39313 4539
rect 39313 4505 39347 4539
rect 39347 4505 39356 4539
rect 39304 4496 39356 4505
rect 39948 4539 40000 4548
rect 39948 4505 39957 4539
rect 39957 4505 39991 4539
rect 39991 4505 40000 4539
rect 39948 4496 40000 4505
rect 38660 4428 38712 4480
rect 41696 4471 41748 4480
rect 41696 4437 41705 4471
rect 41705 4437 41739 4471
rect 41739 4437 41748 4471
rect 41696 4428 41748 4437
rect 42708 4428 42760 4480
rect 11896 4326 11948 4378
rect 11960 4326 12012 4378
rect 12024 4326 12076 4378
rect 12088 4326 12140 4378
rect 12152 4326 12204 4378
rect 22843 4326 22895 4378
rect 22907 4326 22959 4378
rect 22971 4326 23023 4378
rect 23035 4326 23087 4378
rect 23099 4326 23151 4378
rect 33790 4326 33842 4378
rect 33854 4326 33906 4378
rect 33918 4326 33970 4378
rect 33982 4326 34034 4378
rect 34046 4326 34098 4378
rect 44737 4326 44789 4378
rect 44801 4326 44853 4378
rect 44865 4326 44917 4378
rect 44929 4326 44981 4378
rect 44993 4326 45045 4378
rect 10784 4224 10836 4276
rect 11152 4267 11204 4276
rect 11152 4233 11161 4267
rect 11161 4233 11195 4267
rect 11195 4233 11204 4267
rect 11152 4224 11204 4233
rect 11336 4224 11388 4276
rect 12624 4267 12676 4276
rect 12624 4233 12633 4267
rect 12633 4233 12667 4267
rect 12667 4233 12676 4267
rect 12624 4224 12676 4233
rect 13084 4224 13136 4276
rect 15384 4224 15436 4276
rect 16580 4224 16632 4276
rect 17224 4224 17276 4276
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 18052 4267 18104 4276
rect 18052 4233 18061 4267
rect 18061 4233 18095 4267
rect 18095 4233 18104 4267
rect 18052 4224 18104 4233
rect 18604 4267 18656 4276
rect 18604 4233 18613 4267
rect 18613 4233 18647 4267
rect 18647 4233 18656 4267
rect 18604 4224 18656 4233
rect 18880 4267 18932 4276
rect 18880 4233 18889 4267
rect 18889 4233 18923 4267
rect 18923 4233 18932 4267
rect 18880 4224 18932 4233
rect 18972 4224 19024 4276
rect 19708 4224 19760 4276
rect 11244 4156 11296 4208
rect 11796 4199 11848 4208
rect 11796 4165 11805 4199
rect 11805 4165 11839 4199
rect 11839 4165 11848 4199
rect 11796 4156 11848 4165
rect 12532 4199 12584 4208
rect 12532 4165 12541 4199
rect 12541 4165 12575 4199
rect 12575 4165 12584 4199
rect 12532 4156 12584 4165
rect 13268 4199 13320 4208
rect 13268 4165 13277 4199
rect 13277 4165 13311 4199
rect 13311 4165 13320 4199
rect 13268 4156 13320 4165
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9588 4088 9640 4140
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 12624 4020 12676 4072
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 11980 3995 12032 4004
rect 11980 3961 11989 3995
rect 11989 3961 12023 3995
rect 12023 3961 12032 3995
rect 11980 3952 12032 3961
rect 12256 3952 12308 4004
rect 13452 3995 13504 4004
rect 13452 3961 13461 3995
rect 13461 3961 13495 3995
rect 13495 3961 13504 3995
rect 13452 3952 13504 3961
rect 13636 3952 13688 4004
rect 14004 4199 14056 4208
rect 14004 4165 14013 4199
rect 14013 4165 14047 4199
rect 14047 4165 14056 4199
rect 14004 4156 14056 4165
rect 14372 4199 14424 4208
rect 14372 4165 14381 4199
rect 14381 4165 14415 4199
rect 14415 4165 14424 4199
rect 14372 4156 14424 4165
rect 15016 4199 15068 4208
rect 15016 4165 15025 4199
rect 15025 4165 15059 4199
rect 15059 4165 15068 4199
rect 15016 4156 15068 4165
rect 15476 4199 15528 4208
rect 15476 4165 15485 4199
rect 15485 4165 15519 4199
rect 15519 4165 15528 4199
rect 15476 4156 15528 4165
rect 14648 4131 14700 4140
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 15384 4088 15436 4140
rect 15752 4088 15804 4140
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 16580 4020 16632 4072
rect 14188 3995 14240 4004
rect 14188 3961 14197 3995
rect 14197 3961 14231 3995
rect 14231 3961 14240 3995
rect 14188 3952 14240 3961
rect 14556 3995 14608 4004
rect 14556 3961 14565 3995
rect 14565 3961 14599 3995
rect 14599 3961 14608 3995
rect 14556 3952 14608 3961
rect 16764 3952 16816 4004
rect 15568 3884 15620 3936
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 17868 4020 17920 4072
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 19340 4131 19392 4140
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 19432 4020 19484 4072
rect 19524 3952 19576 4004
rect 19800 4088 19852 4140
rect 20812 4156 20864 4208
rect 20904 4156 20956 4208
rect 21272 4156 21324 4208
rect 25044 4224 25096 4276
rect 25504 4224 25556 4276
rect 21916 4156 21968 4208
rect 23940 4088 23992 4140
rect 25872 4224 25924 4276
rect 26240 4224 26292 4276
rect 31024 4224 31076 4276
rect 31392 4224 31444 4276
rect 34520 4224 34572 4276
rect 34336 4156 34388 4208
rect 37096 4224 37148 4276
rect 36728 4156 36780 4208
rect 30472 4088 30524 4140
rect 35716 4131 35768 4140
rect 35716 4097 35725 4131
rect 35725 4097 35759 4131
rect 35759 4097 35768 4131
rect 35716 4088 35768 4097
rect 35992 4131 36044 4140
rect 35992 4097 36001 4131
rect 36001 4097 36035 4131
rect 36035 4097 36044 4131
rect 35992 4088 36044 4097
rect 36268 4131 36320 4140
rect 36268 4097 36277 4131
rect 36277 4097 36311 4131
rect 36311 4097 36320 4131
rect 36268 4088 36320 4097
rect 36544 4131 36596 4140
rect 36544 4097 36553 4131
rect 36553 4097 36587 4131
rect 36587 4097 36596 4131
rect 36544 4088 36596 4097
rect 39120 4131 39172 4140
rect 39120 4097 39129 4131
rect 39129 4097 39163 4131
rect 39163 4097 39172 4131
rect 39120 4088 39172 4097
rect 24400 4020 24452 4072
rect 26700 4020 26752 4072
rect 27344 4020 27396 4072
rect 33692 4020 33744 4072
rect 26240 3952 26292 4004
rect 26516 3952 26568 4004
rect 36084 3952 36136 4004
rect 37188 3952 37240 4004
rect 38200 3952 38252 4004
rect 19892 3884 19944 3936
rect 19984 3884 20036 3936
rect 20812 3927 20864 3936
rect 20812 3893 20821 3927
rect 20821 3893 20855 3927
rect 20855 3893 20864 3927
rect 20812 3884 20864 3893
rect 33140 3884 33192 3936
rect 37280 3884 37332 3936
rect 39672 3884 39724 3936
rect 40408 3884 40460 3936
rect 41420 3884 41472 3936
rect 6423 3782 6475 3834
rect 6487 3782 6539 3834
rect 6551 3782 6603 3834
rect 6615 3782 6667 3834
rect 6679 3782 6731 3834
rect 17370 3782 17422 3834
rect 17434 3782 17486 3834
rect 17498 3782 17550 3834
rect 17562 3782 17614 3834
rect 17626 3782 17678 3834
rect 28317 3782 28369 3834
rect 28381 3782 28433 3834
rect 28445 3782 28497 3834
rect 28509 3782 28561 3834
rect 28573 3782 28625 3834
rect 39264 3782 39316 3834
rect 39328 3782 39380 3834
rect 39392 3782 39444 3834
rect 39456 3782 39508 3834
rect 39520 3782 39572 3834
rect 11336 3680 11388 3732
rect 14740 3680 14792 3732
rect 18788 3680 18840 3732
rect 27252 3680 27304 3732
rect 27344 3680 27396 3732
rect 12992 3612 13044 3664
rect 17224 3612 17276 3664
rect 19340 3612 19392 3664
rect 19432 3612 19484 3664
rect 12624 3476 12676 3528
rect 15752 3408 15804 3460
rect 17132 3476 17184 3528
rect 24400 3476 24452 3528
rect 20720 3408 20772 3460
rect 26240 3544 26292 3596
rect 34612 3680 34664 3732
rect 36544 3680 36596 3732
rect 38200 3680 38252 3732
rect 39120 3680 39172 3732
rect 33416 3544 33468 3596
rect 26976 3408 27028 3460
rect 32496 3476 32548 3528
rect 33600 3519 33652 3528
rect 33600 3485 33609 3519
rect 33609 3485 33643 3519
rect 33643 3485 33652 3519
rect 33600 3476 33652 3485
rect 34152 3476 34204 3528
rect 34244 3408 34296 3460
rect 17960 3340 18012 3392
rect 27896 3340 27948 3392
rect 31484 3383 31536 3392
rect 31484 3349 31493 3383
rect 31493 3349 31527 3383
rect 31527 3349 31536 3383
rect 31484 3340 31536 3349
rect 11896 3238 11948 3290
rect 11960 3238 12012 3290
rect 12024 3238 12076 3290
rect 12088 3238 12140 3290
rect 12152 3238 12204 3290
rect 22843 3238 22895 3290
rect 22907 3238 22959 3290
rect 22971 3238 23023 3290
rect 23035 3238 23087 3290
rect 23099 3238 23151 3290
rect 33790 3238 33842 3290
rect 33854 3238 33906 3290
rect 33918 3238 33970 3290
rect 33982 3238 34034 3290
rect 34046 3238 34098 3290
rect 44737 3238 44789 3290
rect 44801 3238 44853 3290
rect 44865 3238 44917 3290
rect 44929 3238 44981 3290
rect 44993 3238 45045 3290
rect 2688 3136 2740 3188
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 15292 3136 15344 3188
rect 15660 3136 15712 3188
rect 16488 3136 16540 3188
rect 16672 3136 16724 3188
rect 16948 3136 17000 3188
rect 18512 3136 18564 3188
rect 848 3000 900 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11244 3043 11296 3052
rect 11244 3009 11253 3043
rect 11253 3009 11287 3043
rect 11287 3009 11296 3043
rect 11244 3000 11296 3009
rect 17776 3068 17828 3120
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 1676 2907 1728 2916
rect 1676 2873 1685 2907
rect 1685 2873 1719 2907
rect 1719 2873 1728 2907
rect 1676 2864 1728 2873
rect 5632 2907 5684 2916
rect 5632 2873 5641 2907
rect 5641 2873 5675 2907
rect 5675 2873 5684 2907
rect 5632 2864 5684 2873
rect 10508 2907 10560 2916
rect 10508 2873 10517 2907
rect 10517 2873 10551 2907
rect 10551 2873 10560 2907
rect 10508 2864 10560 2873
rect 13176 2864 13228 2916
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 16764 2932 16816 2984
rect 20168 3000 20220 3052
rect 23388 3136 23440 3188
rect 24216 3179 24268 3188
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 25412 3136 25464 3188
rect 31944 3136 31996 3188
rect 32312 3136 32364 3188
rect 23940 3000 23992 3052
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 25504 3043 25556 3052
rect 25504 3009 25513 3043
rect 25513 3009 25547 3043
rect 25547 3009 25556 3043
rect 25504 3000 25556 3009
rect 26240 3043 26292 3052
rect 26240 3009 26249 3043
rect 26249 3009 26283 3043
rect 26283 3009 26292 3043
rect 26240 3000 26292 3009
rect 27160 3043 27212 3052
rect 27160 3009 27169 3043
rect 27169 3009 27203 3043
rect 27203 3009 27212 3043
rect 27160 3000 27212 3009
rect 27712 3043 27764 3052
rect 27712 3009 27721 3043
rect 27721 3009 27755 3043
rect 27755 3009 27764 3043
rect 27712 3000 27764 3009
rect 19708 2932 19760 2984
rect 16856 2864 16908 2916
rect 26056 2839 26108 2848
rect 26056 2805 26065 2839
rect 26065 2805 26099 2839
rect 26099 2805 26108 2839
rect 26056 2796 26108 2805
rect 32496 2839 32548 2848
rect 32496 2805 32505 2839
rect 32505 2805 32539 2839
rect 32539 2805 32548 2839
rect 32496 2796 32548 2805
rect 33048 3136 33100 3188
rect 43168 3136 43220 3188
rect 34796 3043 34848 3052
rect 34796 3009 34805 3043
rect 34805 3009 34839 3043
rect 34839 3009 34848 3043
rect 34796 3000 34848 3009
rect 33324 2796 33376 2848
rect 35532 2796 35584 2848
rect 44640 2864 44692 2916
rect 44272 2839 44324 2848
rect 44272 2805 44281 2839
rect 44281 2805 44315 2839
rect 44315 2805 44324 2839
rect 44272 2796 44324 2805
rect 6423 2694 6475 2746
rect 6487 2694 6539 2746
rect 6551 2694 6603 2746
rect 6615 2694 6667 2746
rect 6679 2694 6731 2746
rect 17370 2694 17422 2746
rect 17434 2694 17486 2746
rect 17498 2694 17550 2746
rect 17562 2694 17614 2746
rect 17626 2694 17678 2746
rect 28317 2694 28369 2746
rect 28381 2694 28433 2746
rect 28445 2694 28497 2746
rect 28509 2694 28561 2746
rect 28573 2694 28625 2746
rect 39264 2694 39316 2746
rect 39328 2694 39380 2746
rect 39392 2694 39444 2746
rect 39456 2694 39508 2746
rect 39520 2694 39572 2746
rect 1952 2592 2004 2644
rect 10324 2592 10376 2644
rect 11060 2592 11112 2644
rect 11796 2592 11848 2644
rect 12532 2592 12584 2644
rect 13268 2592 13320 2644
rect 14004 2592 14056 2644
rect 14372 2635 14424 2644
rect 14372 2601 14381 2635
rect 14381 2601 14415 2635
rect 14415 2601 14424 2635
rect 14372 2592 14424 2601
rect 15476 2592 15528 2644
rect 16212 2592 16264 2644
rect 16580 2592 16632 2644
rect 17132 2635 17184 2644
rect 17132 2601 17141 2635
rect 17141 2601 17175 2635
rect 17175 2601 17184 2635
rect 17132 2592 17184 2601
rect 17224 2592 17276 2644
rect 17776 2592 17828 2644
rect 19708 2592 19760 2644
rect 20168 2592 20220 2644
rect 25504 2592 25556 2644
rect 26240 2592 26292 2644
rect 27160 2592 27212 2644
rect 27712 2592 27764 2644
rect 28908 2635 28960 2644
rect 28908 2601 28917 2635
rect 28917 2601 28951 2635
rect 28951 2601 28960 2635
rect 28908 2592 28960 2601
rect 29184 2592 29236 2644
rect 29920 2592 29972 2644
rect 33140 2592 33192 2644
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 4712 2456 4764 2465
rect 16396 2456 16448 2508
rect 26332 2456 26384 2508
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 5908 2431 5960 2440
rect 5908 2397 5917 2431
rect 5917 2397 5951 2431
rect 5951 2397 5960 2431
rect 5908 2388 5960 2397
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 10508 2431 10560 2440
rect 10508 2397 10517 2431
rect 10517 2397 10551 2431
rect 10551 2397 10560 2431
rect 10508 2388 10560 2397
rect 11520 2431 11572 2440
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 13452 2431 13504 2440
rect 13452 2397 13461 2431
rect 13461 2397 13495 2431
rect 13495 2397 13504 2431
rect 13452 2388 13504 2397
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 16580 2388 16632 2440
rect 17040 2388 17092 2440
rect 17776 2388 17828 2440
rect 18512 2388 18564 2440
rect 19248 2388 19300 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 20996 2431 21048 2440
rect 20996 2397 21005 2431
rect 21005 2397 21039 2431
rect 21039 2397 21048 2431
rect 20996 2388 21048 2397
rect 21456 2388 21508 2440
rect 22192 2388 22244 2440
rect 23204 2431 23256 2440
rect 23204 2397 23213 2431
rect 23213 2397 23247 2431
rect 23247 2397 23256 2431
rect 23204 2388 23256 2397
rect 23664 2388 23716 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 25136 2388 25188 2440
rect 26148 2431 26200 2440
rect 26148 2397 26157 2431
rect 26157 2397 26191 2431
rect 26191 2397 26200 2431
rect 26148 2388 26200 2397
rect 26608 2388 26660 2440
rect 27620 2431 27672 2440
rect 27620 2397 27629 2431
rect 27629 2397 27663 2431
rect 27663 2397 27672 2431
rect 27620 2388 27672 2397
rect 28080 2388 28132 2440
rect 28816 2388 28868 2440
rect 29828 2431 29880 2440
rect 29828 2397 29837 2431
rect 29837 2397 29871 2431
rect 29871 2397 29880 2431
rect 29828 2388 29880 2397
rect 30288 2388 30340 2440
rect 31484 2431 31536 2440
rect 31484 2397 31493 2431
rect 31493 2397 31527 2431
rect 31527 2397 31536 2431
rect 31484 2388 31536 2397
rect 32036 2388 32088 2440
rect 1768 2363 1820 2372
rect 1768 2329 1777 2363
rect 1777 2329 1811 2363
rect 1811 2329 1820 2363
rect 1768 2320 1820 2329
rect 3424 2363 3476 2372
rect 3424 2329 3433 2363
rect 3433 2329 3467 2363
rect 3467 2329 3476 2363
rect 3424 2320 3476 2329
rect 3608 2363 3660 2372
rect 3608 2329 3617 2363
rect 3617 2329 3651 2363
rect 3651 2329 3660 2363
rect 3608 2320 3660 2329
rect 16764 2320 16816 2372
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 16948 2252 17000 2304
rect 20076 2295 20128 2304
rect 20076 2261 20085 2295
rect 20085 2261 20119 2295
rect 20119 2261 20128 2295
rect 20076 2252 20128 2261
rect 20812 2295 20864 2304
rect 20812 2261 20821 2295
rect 20821 2261 20855 2295
rect 20855 2261 20864 2295
rect 20812 2252 20864 2261
rect 21824 2295 21876 2304
rect 21824 2261 21833 2295
rect 21833 2261 21867 2295
rect 21867 2261 21876 2295
rect 21824 2252 21876 2261
rect 31116 2363 31168 2372
rect 31116 2329 31125 2363
rect 31125 2329 31159 2363
rect 31159 2329 31168 2363
rect 31116 2320 31168 2329
rect 32128 2363 32180 2372
rect 32128 2329 32137 2363
rect 32137 2329 32171 2363
rect 32171 2329 32180 2363
rect 32128 2320 32180 2329
rect 32496 2431 32548 2440
rect 32496 2397 32505 2431
rect 32505 2397 32539 2431
rect 32539 2397 32548 2431
rect 32496 2388 32548 2397
rect 32956 2388 33008 2440
rect 33508 2388 33560 2440
rect 34244 2388 34296 2440
rect 34336 2388 34388 2440
rect 34520 2388 34572 2440
rect 36084 2388 36136 2440
rect 37280 2388 37332 2440
rect 39672 2388 39724 2440
rect 40408 2388 40460 2440
rect 41420 2388 41472 2440
rect 41696 2388 41748 2440
rect 42708 2388 42760 2440
rect 43168 2388 43220 2440
rect 24492 2295 24544 2304
rect 24492 2261 24501 2295
rect 24501 2261 24535 2295
rect 24535 2261 24544 2295
rect 24492 2252 24544 2261
rect 32496 2252 32548 2304
rect 33508 2295 33560 2304
rect 33508 2261 33517 2295
rect 33517 2261 33551 2295
rect 33551 2261 33560 2295
rect 33508 2252 33560 2261
rect 34244 2295 34296 2304
rect 34244 2261 34253 2295
rect 34253 2261 34287 2295
rect 34287 2261 34296 2295
rect 34244 2252 34296 2261
rect 34980 2295 35032 2304
rect 34980 2261 34989 2295
rect 34989 2261 35023 2295
rect 35023 2261 35032 2295
rect 34980 2252 35032 2261
rect 35900 2295 35952 2304
rect 35900 2261 35909 2295
rect 35909 2261 35943 2295
rect 35943 2261 35952 2295
rect 35900 2252 35952 2261
rect 36452 2295 36504 2304
rect 36452 2261 36461 2295
rect 36461 2261 36495 2295
rect 36495 2261 36504 2295
rect 36452 2252 36504 2261
rect 37188 2252 37240 2304
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 38384 2252 38436 2304
rect 39396 2295 39448 2304
rect 39396 2261 39405 2295
rect 39405 2261 39439 2295
rect 39439 2261 39448 2295
rect 39396 2252 39448 2261
rect 39856 2252 39908 2304
rect 40868 2295 40920 2304
rect 40868 2261 40877 2295
rect 40877 2261 40911 2295
rect 40911 2261 40920 2295
rect 40868 2252 40920 2261
rect 41328 2252 41380 2304
rect 42432 2252 42484 2304
rect 43168 2295 43220 2304
rect 43168 2261 43177 2295
rect 43177 2261 43211 2295
rect 43211 2261 43220 2295
rect 43168 2252 43220 2261
rect 43812 2295 43864 2304
rect 43812 2261 43821 2295
rect 43821 2261 43855 2295
rect 43855 2261 43864 2295
rect 43812 2252 43864 2261
rect 11896 2150 11948 2202
rect 11960 2150 12012 2202
rect 12024 2150 12076 2202
rect 12088 2150 12140 2202
rect 12152 2150 12204 2202
rect 22843 2150 22895 2202
rect 22907 2150 22959 2202
rect 22971 2150 23023 2202
rect 23035 2150 23087 2202
rect 23099 2150 23151 2202
rect 33790 2150 33842 2202
rect 33854 2150 33906 2202
rect 33918 2150 33970 2202
rect 33982 2150 34034 2202
rect 34046 2150 34098 2202
rect 44737 2150 44789 2202
rect 44801 2150 44853 2202
rect 44865 2150 44917 2202
rect 44929 2150 44981 2202
rect 44993 2150 45045 2202
rect 7932 2048 7984 2100
rect 15384 2048 15436 2100
rect 20076 2048 20128 2100
rect 24032 1980 24084 2032
rect 15752 1912 15804 1964
rect 21824 1912 21876 1964
rect 12808 1844 12860 1896
rect 20812 1844 20864 1896
rect 16856 1776 16908 1828
rect 24492 1776 24544 1828
rect 1676 1300 1728 1352
rect 33600 1300 33652 1352
rect 3608 1232 3660 1284
rect 34796 1232 34848 1284
rect 5632 1164 5684 1216
rect 35716 1164 35768 1216
<< metal2 >>
rect 5722 7840 5778 8000
rect 5998 7840 6054 8000
rect 6274 7840 6330 8000
rect 6550 7840 6606 8000
rect 6826 7840 6882 8000
rect 7102 7970 7158 8000
rect 7102 7942 7328 7970
rect 7102 7840 7158 7942
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 848 3052 900 3058
rect 848 2994 900 3000
rect 860 160 888 2994
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1688 1358 1716 2858
rect 1964 2650 1992 6190
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 3194 2728 6122
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 4172 3058 4200 6258
rect 5736 4758 5764 7840
rect 5908 6520 5960 6526
rect 5908 6462 5960 6468
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5920 4622 5948 6462
rect 6012 5370 6040 7840
rect 6182 5808 6238 5817
rect 6182 5743 6238 5752
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6104 4826 6132 5170
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6196 4622 6224 5743
rect 6288 4758 6316 7840
rect 6564 5166 6592 7840
rect 6734 5672 6790 5681
rect 6734 5607 6790 5616
rect 6748 5234 6776 5607
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6423 4924 6731 4933
rect 6423 4922 6429 4924
rect 6485 4922 6509 4924
rect 6565 4922 6589 4924
rect 6645 4922 6669 4924
rect 6725 4922 6731 4924
rect 6485 4870 6487 4922
rect 6667 4870 6669 4922
rect 6423 4868 6429 4870
rect 6485 4868 6509 4870
rect 6565 4868 6589 4870
rect 6645 4868 6669 4870
rect 6725 4868 6731 4870
rect 6423 4859 6731 4868
rect 6840 4758 6868 7840
rect 7010 5264 7066 5273
rect 7010 5199 7012 5208
rect 7064 5199 7066 5208
rect 7012 5170 7064 5176
rect 7300 4826 7328 7942
rect 7378 7840 7434 8000
rect 7654 7970 7710 8000
rect 7654 7942 7880 7970
rect 7654 7840 7710 7942
rect 7392 5370 7420 7840
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 7668 4554 7696 6326
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7760 5302 7788 5578
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 7852 4826 7880 7942
rect 7930 7840 7986 8000
rect 8206 7840 8262 8000
rect 8482 7840 8538 8000
rect 8758 7970 8814 8000
rect 8758 7942 8892 7970
rect 8758 7840 8814 7942
rect 7944 5370 7972 7840
rect 8116 6044 8168 6050
rect 8116 5986 8168 5992
rect 8024 5976 8076 5982
rect 8024 5918 8076 5924
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 8036 4622 8064 5918
rect 8128 4622 8156 5986
rect 8220 4808 8248 7840
rect 8496 5370 8524 7840
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8392 4820 8444 4826
rect 8220 4780 8392 4808
rect 8392 4762 8444 4768
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 8864 4146 8892 7942
rect 9034 7840 9090 8000
rect 9310 7840 9366 8000
rect 9586 7840 9642 8000
rect 9862 7840 9918 8000
rect 10138 7840 10194 8000
rect 10414 7840 10470 8000
rect 10690 7970 10746 8000
rect 10520 7942 10746 7970
rect 9048 5370 9076 7840
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9324 4826 9352 7840
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9416 5302 9444 5646
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9508 4622 9536 6394
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9416 4457 9444 4490
rect 9402 4448 9458 4457
rect 9402 4383 9458 4392
rect 9600 4146 9628 7840
rect 9876 4826 9904 7840
rect 10152 5370 10180 7840
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10428 4826 10456 7840
rect 10520 5234 10548 7942
rect 10690 7840 10746 7942
rect 10966 7840 11022 8000
rect 11242 7840 11298 8000
rect 11518 7970 11574 8000
rect 11440 7942 11574 7970
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 10416 4820 10468 4826
rect 10980 4808 11008 7840
rect 11256 5370 11284 7840
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11060 4820 11112 4826
rect 10980 4780 11060 4808
rect 10416 4762 10468 4768
rect 11060 4762 11112 4768
rect 10784 4548 10836 4554
rect 10784 4490 10836 4496
rect 10796 4282 10824 4490
rect 11164 4282 11192 5170
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11256 4729 11284 4966
rect 11242 4720 11298 4729
rect 11242 4655 11298 4664
rect 11348 4282 11376 5170
rect 11440 4826 11468 7942
rect 11518 7840 11574 7942
rect 11794 7840 11850 8000
rect 12070 7970 12126 8000
rect 12070 7942 12296 7970
rect 12070 7840 12126 7942
rect 11808 5250 11836 7840
rect 11896 5468 12204 5477
rect 11896 5466 11902 5468
rect 11958 5466 11982 5468
rect 12038 5466 12062 5468
rect 12118 5466 12142 5468
rect 12198 5466 12204 5468
rect 11958 5414 11960 5466
rect 12140 5414 12142 5466
rect 11896 5412 11902 5414
rect 11958 5412 11982 5414
rect 12038 5412 12062 5414
rect 12118 5412 12142 5414
rect 12198 5412 12204 5414
rect 11896 5403 12204 5412
rect 11624 5234 11836 5250
rect 11612 5228 11836 5234
rect 11664 5222 11836 5228
rect 11612 5170 11664 5176
rect 11520 5024 11572 5030
rect 11888 5024 11940 5030
rect 11520 4966 11572 4972
rect 11886 4992 11888 5001
rect 11940 4992 11942 5001
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11532 4706 11560 4966
rect 11886 4927 11942 4936
rect 11702 4856 11758 4865
rect 11702 4791 11758 4800
rect 12072 4820 12124 4826
rect 11716 4758 11744 4791
rect 12268 4808 12296 7942
rect 12346 7840 12402 8000
rect 12622 7970 12678 8000
rect 12544 7942 12678 7970
rect 12360 5522 12388 7840
rect 12360 5494 12480 5522
rect 12452 4826 12480 5494
rect 12544 5370 12572 7942
rect 12622 7840 12678 7942
rect 12898 7840 12954 8000
rect 13174 7840 13230 8000
rect 13450 7970 13506 8000
rect 13450 7942 13584 7970
rect 13450 7840 13506 7942
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 12124 4780 12296 4808
rect 12440 4820 12492 4826
rect 12072 4762 12124 4768
rect 12440 4762 12492 4768
rect 11440 4678 11560 4706
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 12346 4720 12402 4729
rect 11440 4622 11468 4678
rect 12402 4678 12480 4706
rect 12346 4655 12402 4664
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 12256 4548 12308 4554
rect 12256 4490 12308 4496
rect 11896 4380 12204 4389
rect 11896 4378 11902 4380
rect 11958 4378 11982 4380
rect 12038 4378 12062 4380
rect 12118 4378 12142 4380
rect 12198 4378 12204 4380
rect 11958 4326 11960 4378
rect 12140 4326 12142 4378
rect 11896 4324 11902 4326
rect 11958 4324 11982 4326
rect 12038 4324 12062 4326
rect 12118 4324 12142 4326
rect 12198 4324 12204 4326
rect 11896 4315 12204 4324
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11244 4208 11296 4214
rect 11242 4176 11244 4185
rect 11796 4208 11848 4214
rect 11296 4176 11298 4185
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 9588 4140 9640 4146
rect 11796 4150 11848 4156
rect 11242 4111 11298 4120
rect 11336 4140 11388 4146
rect 9588 4082 9640 4088
rect 11336 4082 11388 4088
rect 6423 3836 6731 3845
rect 6423 3834 6429 3836
rect 6485 3834 6509 3836
rect 6565 3834 6589 3836
rect 6645 3834 6669 3836
rect 6725 3834 6731 3836
rect 6485 3782 6487 3834
rect 6667 3782 6669 3834
rect 6423 3780 6429 3782
rect 6485 3780 6509 3782
rect 6565 3780 6589 3782
rect 6645 3780 6669 3782
rect 6725 3780 6731 3782
rect 6423 3771 6731 3780
rect 11348 3738 11376 4082
rect 11336 3732 11388 3738
rect 11336 3674 11388 3680
rect 11242 3088 11298 3097
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 11060 3052 11112 3058
rect 11242 3023 11244 3032
rect 11060 2994 11112 3000
rect 11296 3023 11298 3032
rect 11244 2994 11296 3000
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 1676 1352 1728 1358
rect 1676 1294 1728 1300
rect 846 0 902 160
rect 1582 82 1638 160
rect 1780 82 1808 2314
rect 1582 54 1808 82
rect 2318 82 2374 160
rect 2516 82 2544 2994
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 3424 2372 3476 2378
rect 3424 2314 3476 2320
rect 3608 2372 3660 2378
rect 3608 2314 3660 2320
rect 2318 54 2544 82
rect 3054 82 3110 160
rect 3436 82 3464 2314
rect 3620 1290 3648 2314
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 3054 54 3464 82
rect 3790 82 3846 160
rect 3896 82 3924 2926
rect 4710 2544 4766 2553
rect 4710 2479 4712 2488
rect 4764 2479 4766 2488
rect 4712 2450 4764 2456
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 3790 54 3924 82
rect 4448 82 4476 2382
rect 4526 82 4582 160
rect 4448 54 4582 82
rect 1582 0 1638 54
rect 2318 0 2374 54
rect 3054 0 3110 54
rect 3790 0 3846 54
rect 4526 0 4582 54
rect 5262 82 5318 160
rect 5460 82 5488 2994
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5644 1222 5672 2858
rect 6423 2748 6731 2757
rect 6423 2746 6429 2748
rect 6485 2746 6509 2748
rect 6565 2746 6589 2748
rect 6645 2746 6669 2748
rect 6725 2746 6731 2748
rect 6485 2694 6487 2746
rect 6667 2694 6669 2746
rect 6423 2692 6429 2694
rect 6485 2692 6509 2694
rect 6565 2692 6589 2694
rect 6645 2692 6669 2694
rect 6725 2692 6731 2694
rect 6423 2683 6731 2692
rect 10336 2650 10364 2994
rect 10506 2952 10562 2961
rect 10506 2887 10508 2896
rect 10560 2887 10562 2896
rect 10508 2858 10560 2864
rect 11072 2650 11100 2994
rect 11808 2650 11836 4150
rect 12268 4010 12296 4490
rect 12452 4321 12480 4678
rect 12438 4312 12494 4321
rect 12636 4282 12664 5714
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12438 4247 12494 4256
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 11980 4004 12032 4010
rect 11980 3946 12032 3952
rect 12256 4004 12308 4010
rect 12256 3946 12308 3952
rect 11992 3641 12020 3946
rect 11978 3632 12034 3641
rect 11978 3567 12034 3576
rect 11896 3292 12204 3301
rect 11896 3290 11902 3292
rect 11958 3290 11982 3292
rect 12038 3290 12062 3292
rect 12118 3290 12142 3292
rect 12198 3290 12204 3292
rect 11958 3238 11960 3290
rect 12140 3238 12142 3290
rect 11896 3236 11902 3238
rect 11958 3236 11982 3238
rect 12038 3236 12062 3238
rect 12118 3236 12142 3238
rect 12198 3236 12204 3238
rect 11896 3227 12204 3236
rect 12544 2650 12572 4150
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 12636 3534 12664 4014
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12728 3194 12756 4490
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 5908 2440 5960 2446
rect 5906 2408 5908 2417
rect 6184 2440 6236 2446
rect 5960 2408 5962 2417
rect 6184 2382 6236 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7748 2440 7800 2446
rect 8300 2440 8352 2446
rect 7748 2382 7800 2388
rect 8220 2400 8300 2428
rect 5906 2343 5962 2352
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 5262 54 5488 82
rect 5998 82 6054 160
rect 6196 82 6224 2382
rect 5998 54 6224 82
rect 6734 82 6790 160
rect 6840 82 6868 2382
rect 7116 1737 7144 2382
rect 7102 1728 7158 1737
rect 7102 1663 7158 1672
rect 6734 54 6868 82
rect 7470 82 7526 160
rect 7760 82 7788 2382
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 2106 7972 2246
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8220 160 8248 2400
rect 8300 2382 8352 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 11520 2440 11572 2446
rect 11980 2440 12032 2446
rect 11520 2382 11572 2388
rect 11808 2400 11980 2428
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 2009 8524 2246
rect 8482 2000 8538 2009
rect 8482 1935 8538 1944
rect 7470 54 7788 82
rect 5262 0 5318 54
rect 5998 0 6054 54
rect 6734 0 6790 54
rect 7470 0 7526 54
rect 8206 0 8262 160
rect 8942 82 8998 160
rect 9048 82 9076 2382
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1873 9260 2246
rect 9218 1864 9274 1873
rect 9218 1799 9274 1808
rect 8942 54 9076 82
rect 9678 82 9734 160
rect 9784 82 9812 2382
rect 9678 54 9812 82
rect 10414 82 10470 160
rect 10520 82 10548 2382
rect 10414 54 10548 82
rect 11150 82 11206 160
rect 11532 82 11560 2382
rect 11150 54 11560 82
rect 11808 82 11836 2400
rect 11980 2382 12032 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 11896 2204 12204 2213
rect 11896 2202 11902 2204
rect 11958 2202 11982 2204
rect 12038 2202 12062 2204
rect 12118 2202 12142 2204
rect 12198 2202 12204 2204
rect 11958 2150 11960 2202
rect 12140 2150 12142 2202
rect 11896 2148 11902 2150
rect 11958 2148 11982 2150
rect 12038 2148 12062 2150
rect 12118 2148 12142 2150
rect 12198 2148 12204 2150
rect 11896 2139 12204 2148
rect 11886 82 11942 160
rect 11808 54 11942 82
rect 8942 0 8998 54
rect 9678 0 9734 54
rect 10414 0 10470 54
rect 11150 0 11206 54
rect 11886 0 11942 54
rect 12622 82 12678 160
rect 12728 82 12756 2382
rect 12820 1902 12848 4966
rect 12912 4808 12940 7840
rect 13188 5370 13216 7840
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12992 4820 13044 4826
rect 12912 4780 12992 4808
rect 12992 4762 13044 4768
rect 13096 4282 13124 5170
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 13004 3670 13032 4082
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 13188 2922 13216 5170
rect 13268 5092 13320 5098
rect 13320 5052 13400 5080
rect 13268 5034 13320 5040
rect 13266 4584 13322 4593
rect 13372 4554 13400 5052
rect 13556 4826 13584 7942
rect 13726 7840 13782 8000
rect 14002 7840 14058 8000
rect 14278 7840 14334 8000
rect 14554 7970 14610 8000
rect 14554 7942 14688 7970
rect 14554 7840 14610 7942
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5302 13676 6054
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13740 5030 13768 7840
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13266 4519 13268 4528
rect 13320 4519 13322 4528
rect 13360 4548 13412 4554
rect 13268 4490 13320 4496
rect 13360 4490 13412 4496
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 13280 2650 13308 4150
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13636 4004 13688 4010
rect 13832 3992 13860 4966
rect 14016 4808 14044 7840
rect 14292 5370 14320 7840
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14188 4820 14240 4826
rect 14016 4780 14188 4808
rect 14188 4762 14240 4768
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 14372 4208 14424 4214
rect 14372 4150 14424 4156
rect 13688 3964 13860 3992
rect 13636 3946 13688 3952
rect 13464 3641 13492 3946
rect 13450 3632 13506 3641
rect 13450 3567 13506 3576
rect 14016 2650 14044 4150
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 14200 3913 14228 3946
rect 14186 3904 14242 3913
rect 14186 3839 14242 3848
rect 14384 2650 14412 4150
rect 14660 4146 14688 7942
rect 14830 7840 14886 8000
rect 15106 7840 15162 8000
rect 15382 7840 15438 8000
rect 15658 7840 15714 8000
rect 15934 7840 15990 8000
rect 16210 7840 16266 8000
rect 16486 7840 16542 8000
rect 16762 7840 16818 8000
rect 17038 7840 17094 8000
rect 17314 7840 17370 8000
rect 17590 7840 17646 8000
rect 17866 7840 17922 8000
rect 18142 7840 18198 8000
rect 18418 7840 18474 8000
rect 18694 7840 18750 8000
rect 18970 7970 19026 8000
rect 18892 7942 19026 7970
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14568 3505 14596 3946
rect 14752 3738 14780 5170
rect 14844 4758 14872 7840
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14832 4752 14884 4758
rect 14832 4694 14884 4700
rect 14936 4622 14964 5510
rect 15120 5370 15148 7840
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15106 5128 15162 5137
rect 15028 5086 15106 5114
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15028 4214 15056 5086
rect 15106 5063 15162 5072
rect 15106 4720 15162 4729
rect 15106 4655 15108 4664
rect 15160 4655 15162 4664
rect 15108 4626 15160 4632
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14554 3496 14610 3505
rect 14554 3431 14610 3440
rect 15212 3233 15240 5170
rect 15198 3224 15254 3233
rect 15304 3194 15332 5170
rect 15396 4758 15424 7840
rect 15672 5370 15700 7840
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15384 4752 15436 4758
rect 15384 4694 15436 4700
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15396 4282 15424 4558
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15198 3159 15254 3168
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 12808 1896 12860 1902
rect 12808 1838 12860 1844
rect 12622 54 12756 82
rect 13358 82 13414 160
rect 13464 82 13492 2382
rect 13358 54 13492 82
rect 14094 82 14150 160
rect 14200 82 14228 2382
rect 14094 54 14228 82
rect 14830 82 14886 160
rect 14936 82 14964 2382
rect 15396 2106 15424 4082
rect 15488 2650 15516 4150
rect 15580 3942 15608 4558
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15672 3194 15700 4626
rect 15764 4146 15792 5782
rect 15948 4826 15976 7840
rect 16224 5370 16252 7840
rect 16396 5908 16448 5914
rect 16396 5850 16448 5856
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 16026 4992 16082 5001
rect 16026 4927 16082 4936
rect 16040 4826 16068 4927
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 16212 4140 16264 4146
rect 16212 4082 16264 4088
rect 16224 3482 16252 4082
rect 16408 3618 16436 5850
rect 16500 4758 16528 7840
rect 16776 5370 16804 7840
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16948 5296 17000 5302
rect 16948 5238 17000 5244
rect 16578 4856 16634 4865
rect 16578 4791 16634 4800
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16592 4282 16620 4791
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16408 3590 16528 3618
rect 15752 3460 15804 3466
rect 16224 3454 16436 3482
rect 15752 3402 15804 3408
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15660 2440 15712 2446
rect 15580 2400 15660 2428
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15580 160 15608 2400
rect 15660 2382 15712 2388
rect 15764 1970 15792 3402
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16224 2650 16252 2994
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16408 2514 16436 3454
rect 16500 3194 16528 3590
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16592 2650 16620 4014
rect 16684 3194 16712 4490
rect 16764 4004 16816 4010
rect 16816 3964 16896 3992
rect 16764 3946 16816 3952
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16868 3074 16896 3964
rect 16960 3194 16988 5238
rect 17052 4758 17080 7840
rect 17328 6202 17356 7840
rect 17236 6174 17356 6202
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 17144 4690 17172 5238
rect 17236 4808 17264 6174
rect 17604 5370 17632 7840
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17370 4924 17678 4933
rect 17370 4922 17376 4924
rect 17432 4922 17456 4924
rect 17512 4922 17536 4924
rect 17592 4922 17616 4924
rect 17672 4922 17678 4924
rect 17432 4870 17434 4922
rect 17614 4870 17616 4922
rect 17370 4868 17376 4870
rect 17432 4868 17456 4870
rect 17512 4868 17536 4870
rect 17592 4868 17616 4870
rect 17672 4868 17678 4870
rect 17370 4859 17678 4868
rect 17316 4820 17368 4826
rect 17236 4780 17316 4808
rect 17316 4762 17368 4768
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 17224 4548 17276 4554
rect 17224 4490 17276 4496
rect 17236 4282 17264 4490
rect 17788 4282 17816 5170
rect 17880 4826 17908 7840
rect 18156 5370 18184 7840
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17972 4706 18000 5170
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 17880 4678 18000 4706
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17880 4078 17908 4678
rect 18340 4622 18368 5102
rect 18432 4826 18460 7840
rect 18708 5370 18736 7840
rect 18892 5370 18920 7942
rect 18970 7840 19026 7942
rect 19246 7840 19302 8000
rect 19522 7840 19578 8000
rect 19798 7840 19854 8000
rect 20074 7840 20130 8000
rect 20350 7840 20406 8000
rect 20626 7840 20682 8000
rect 20902 7840 20958 8000
rect 21178 7840 21234 8000
rect 21454 7970 21510 8000
rect 21454 7942 21680 7970
rect 21454 7840 21510 7942
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 19260 5302 19288 7840
rect 19338 5808 19394 5817
rect 19338 5743 19394 5752
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18064 4282 18092 4558
rect 18800 4554 18828 4762
rect 18604 4548 18656 4554
rect 18604 4490 18656 4496
rect 18788 4548 18840 4554
rect 18788 4490 18840 4496
rect 18616 4282 18644 4490
rect 18892 4282 18920 5170
rect 18984 4282 19012 5170
rect 19352 4758 19380 5743
rect 19536 5370 19564 7840
rect 19812 6474 19840 7840
rect 19984 6520 20036 6526
rect 19812 6446 19932 6474
rect 19984 6462 20036 6468
rect 19614 5672 19670 5681
rect 19614 5607 19670 5616
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19522 4992 19578 5001
rect 19444 4950 19522 4978
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 19444 4162 19472 4950
rect 19522 4927 19578 4936
rect 19628 4622 19656 5607
rect 19798 5400 19854 5409
rect 19798 5335 19854 5344
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19524 4480 19576 4486
rect 19576 4440 19656 4468
rect 19524 4422 19576 4428
rect 19628 4162 19656 4440
rect 19720 4282 19748 5170
rect 19812 4826 19840 5335
rect 19904 5302 19932 6446
rect 19892 5296 19944 5302
rect 19892 5238 19944 5244
rect 19890 4856 19946 4865
rect 19800 4820 19852 4826
rect 19890 4791 19946 4800
rect 19800 4762 19852 4768
rect 19904 4758 19932 4791
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19708 4276 19760 4282
rect 19708 4218 19760 4224
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 19340 4140 19392 4146
rect 19444 4134 19564 4162
rect 19628 4146 19840 4162
rect 19628 4140 19852 4146
rect 19628 4134 19800 4140
rect 19340 4082 19392 4088
rect 17868 4072 17920 4078
rect 17868 4014 17920 4020
rect 17370 3836 17678 3845
rect 17370 3834 17376 3836
rect 17432 3834 17456 3836
rect 17512 3834 17536 3836
rect 17592 3834 17616 3836
rect 17672 3834 17678 3836
rect 17432 3782 17434 3834
rect 17614 3782 17616 3834
rect 17370 3780 17376 3782
rect 17432 3780 17456 3782
rect 17512 3780 17536 3782
rect 17592 3780 17616 3782
rect 17672 3780 17678 3782
rect 17370 3771 17678 3780
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16868 3046 16988 3074
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 16592 1442 16620 2382
rect 16776 2378 16804 2926
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 16868 1834 16896 2858
rect 16960 2310 16988 3046
rect 17144 2650 17172 3470
rect 17236 2650 17264 3606
rect 17972 3398 18000 4082
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 17960 3392 18012 3398
rect 18248 3369 18276 3975
rect 17960 3334 18012 3340
rect 18234 3360 18290 3369
rect 18234 3295 18290 3304
rect 18524 3194 18552 4082
rect 18800 3738 18828 4082
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 19352 3670 19380 4082
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19444 3670 19472 4014
rect 19536 4010 19564 4134
rect 19800 4082 19852 4088
rect 19524 4004 19576 4010
rect 19524 3946 19576 3952
rect 19904 3942 19932 4422
rect 19996 3942 20024 6462
rect 20088 4622 20116 7840
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20180 4672 20208 5170
rect 20260 4684 20312 4690
rect 20180 4644 20260 4672
rect 20260 4626 20312 4632
rect 20364 4622 20392 7840
rect 20442 5400 20498 5409
rect 20442 5335 20498 5344
rect 20456 4826 20484 5335
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20548 4622 20576 4966
rect 20640 4622 20668 7840
rect 20916 5114 20944 7840
rect 21192 5216 21220 7840
rect 21652 5234 21680 7942
rect 21730 7840 21786 8000
rect 22006 7840 22062 8000
rect 22282 7840 22338 8000
rect 22558 7840 22614 8000
rect 22834 7840 22890 8000
rect 23110 7840 23166 8000
rect 23386 7840 23442 8000
rect 23662 7840 23718 8000
rect 23938 7840 23994 8000
rect 24214 7840 24270 8000
rect 24490 7970 24546 8000
rect 24490 7942 24716 7970
rect 24490 7840 24546 7942
rect 21744 5234 21772 7840
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21364 5228 21416 5234
rect 21192 5188 21364 5216
rect 21364 5170 21416 5176
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 20916 5086 21404 5114
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20076 4480 20128 4486
rect 20260 4480 20312 4486
rect 20128 4440 20260 4468
rect 20076 4422 20128 4428
rect 20260 4422 20312 4428
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 20732 3466 20760 4966
rect 20824 4554 21128 4570
rect 20812 4548 21128 4554
rect 20864 4542 21128 4548
rect 20812 4490 20864 4496
rect 21100 4486 21128 4542
rect 20904 4480 20956 4486
rect 20904 4422 20956 4428
rect 21088 4480 21140 4486
rect 21088 4422 21140 4428
rect 20916 4214 20944 4422
rect 21284 4214 21312 4966
rect 21376 4622 21404 5086
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21454 4856 21510 4865
rect 21454 4791 21510 4800
rect 21468 4758 21496 4791
rect 21456 4752 21508 4758
rect 21456 4694 21508 4700
rect 21836 4690 21864 4966
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21928 4214 21956 5306
rect 22020 5216 22048 7840
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22100 5228 22152 5234
rect 22020 5188 22100 5216
rect 22100 5170 22152 5176
rect 22204 5114 22232 5646
rect 22296 5216 22324 7840
rect 22572 6610 22600 7840
rect 22848 6610 22876 7840
rect 22572 6582 22692 6610
rect 22560 5228 22612 5234
rect 22296 5188 22560 5216
rect 22664 5216 22692 6582
rect 22756 6582 22876 6610
rect 23124 6610 23152 7840
rect 23124 6582 23244 6610
rect 22756 5352 22784 6582
rect 22843 5468 23151 5477
rect 22843 5466 22849 5468
rect 22905 5466 22929 5468
rect 22985 5466 23009 5468
rect 23065 5466 23089 5468
rect 23145 5466 23151 5468
rect 22905 5414 22907 5466
rect 23087 5414 23089 5466
rect 22843 5412 22849 5414
rect 22905 5412 22929 5414
rect 22985 5412 23009 5414
rect 23065 5412 23089 5414
rect 23145 5412 23151 5414
rect 22843 5403 23151 5412
rect 22756 5324 23152 5352
rect 23124 5234 23152 5324
rect 22836 5228 22888 5234
rect 22664 5188 22836 5216
rect 22560 5170 22612 5176
rect 22836 5170 22888 5176
rect 23112 5228 23164 5234
rect 23216 5216 23244 6582
rect 23400 5522 23428 7840
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23400 5494 23520 5522
rect 23492 5234 23520 5494
rect 23388 5228 23440 5234
rect 23216 5188 23388 5216
rect 23112 5170 23164 5176
rect 23388 5170 23440 5176
rect 23480 5228 23532 5234
rect 23480 5170 23532 5176
rect 23020 5160 23072 5166
rect 22008 5092 22060 5098
rect 22204 5086 22508 5114
rect 23020 5102 23072 5108
rect 23386 5128 23442 5137
rect 22008 5034 22060 5040
rect 22020 4865 22048 5034
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22006 4856 22062 4865
rect 22112 4826 22140 4966
rect 22204 4865 22232 4966
rect 22190 4856 22246 4865
rect 22006 4791 22062 4800
rect 22100 4820 22152 4826
rect 22190 4791 22246 4800
rect 22100 4762 22152 4768
rect 22388 4622 22416 4966
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22480 4486 22508 5086
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22664 4826 22692 4966
rect 22940 4826 22968 4966
rect 23032 4865 23060 5102
rect 23386 5063 23442 5072
rect 23204 5024 23256 5030
rect 23204 4966 23256 4972
rect 23018 4856 23074 4865
rect 22652 4820 22704 4826
rect 22652 4762 22704 4768
rect 22928 4820 22980 4826
rect 23216 4826 23244 4966
rect 23018 4791 23074 4800
rect 23204 4820 23256 4826
rect 22928 4762 22980 4768
rect 23204 4762 23256 4768
rect 22284 4480 22336 4486
rect 22282 4448 22284 4457
rect 22468 4480 22520 4486
rect 22336 4448 22338 4457
rect 22468 4422 22520 4428
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 22282 4383 22338 4392
rect 22664 4321 22692 4422
rect 22650 4312 22706 4321
rect 22650 4247 22706 4256
rect 20812 4208 20864 4214
rect 20812 4150 20864 4156
rect 20904 4208 20956 4214
rect 20904 4150 20956 4156
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21916 4208 21968 4214
rect 22756 4185 22784 4422
rect 22843 4380 23151 4389
rect 22843 4378 22849 4380
rect 22905 4378 22929 4380
rect 22985 4378 23009 4380
rect 23065 4378 23089 4380
rect 23145 4378 23151 4380
rect 22905 4326 22907 4378
rect 23087 4326 23089 4378
rect 22843 4324 22849 4326
rect 22905 4324 22929 4326
rect 22985 4324 23009 4326
rect 23065 4324 23089 4326
rect 23145 4324 23151 4326
rect 22843 4315 23151 4324
rect 21916 4150 21968 4156
rect 22742 4176 22798 4185
rect 20824 3942 20852 4150
rect 22742 4111 22798 4120
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 22843 3292 23151 3301
rect 22843 3290 22849 3292
rect 22905 3290 22929 3292
rect 22985 3290 23009 3292
rect 23065 3290 23089 3292
rect 23145 3290 23151 3292
rect 22905 3238 22907 3290
rect 23087 3238 23089 3290
rect 22843 3236 22849 3238
rect 22905 3236 22929 3238
rect 22985 3236 23009 3238
rect 23065 3236 23089 3238
rect 23145 3236 23151 3238
rect 22650 3224 22706 3233
rect 22843 3227 23151 3236
rect 18512 3188 18564 3194
rect 23400 3194 23428 5063
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 4826 23520 4966
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 23584 4622 23612 6394
rect 23676 5658 23704 7840
rect 23676 5630 23796 5658
rect 23768 5234 23796 5630
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23768 4826 23796 4966
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23860 4486 23888 5578
rect 23952 5216 23980 7840
rect 24228 6610 24256 7840
rect 24228 6582 24348 6610
rect 24124 6044 24176 6050
rect 24124 5986 24176 5992
rect 24032 5228 24084 5234
rect 23952 5188 24032 5216
rect 24032 5170 24084 5176
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24044 4826 24072 4966
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24136 4554 24164 5986
rect 24320 5234 24348 6582
rect 24398 5264 24454 5273
rect 24308 5228 24360 5234
rect 24454 5222 24532 5250
rect 24398 5199 24454 5208
rect 24308 5170 24360 5176
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24412 4826 24440 4966
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24504 4622 24532 5222
rect 24688 5216 24716 7942
rect 24766 7840 24822 8000
rect 25042 7840 25098 8000
rect 25318 7840 25374 8000
rect 25594 7970 25650 8000
rect 25870 7970 25926 8000
rect 25594 7942 25820 7970
rect 25594 7840 25650 7942
rect 24780 5370 24808 7840
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 24860 5228 24912 5234
rect 24688 5188 24860 5216
rect 24860 5170 24912 5176
rect 24964 5114 24992 5238
rect 25056 5166 25084 7840
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 25136 5976 25188 5982
rect 25136 5918 25188 5924
rect 24872 5086 24992 5114
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4826 24716 4966
rect 24872 4826 24900 5086
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24860 4820 24912 4826
rect 24860 4762 24912 4768
rect 24964 4758 24992 4966
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 24492 4616 24544 4622
rect 24492 4558 24544 4564
rect 24124 4548 24176 4554
rect 24124 4490 24176 4496
rect 25044 4548 25096 4554
rect 25044 4490 25096 4496
rect 23848 4480 23900 4486
rect 23848 4422 23900 4428
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24214 4176 24270 4185
rect 23940 4140 23992 4146
rect 24964 4162 24992 4422
rect 25056 4282 25084 4490
rect 25148 4486 25176 5918
rect 25240 5114 25268 6326
rect 25332 5302 25360 7840
rect 25412 5568 25464 5574
rect 25412 5510 25464 5516
rect 25320 5296 25372 5302
rect 25320 5238 25372 5244
rect 25240 5086 25360 5114
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25240 4758 25268 4966
rect 25228 4752 25280 4758
rect 25228 4694 25280 4700
rect 25136 4480 25188 4486
rect 25136 4422 25188 4428
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 25332 4162 25360 5086
rect 24964 4134 25360 4162
rect 24214 4111 24270 4120
rect 23940 4082 23992 4088
rect 22650 3159 22706 3168
rect 23388 3188 23440 3194
rect 18512 3130 18564 3136
rect 17776 3120 17828 3126
rect 17776 3062 17828 3068
rect 17370 2748 17678 2757
rect 17370 2746 17376 2748
rect 17432 2746 17456 2748
rect 17512 2746 17536 2748
rect 17592 2746 17616 2748
rect 17672 2746 17678 2748
rect 17432 2694 17434 2746
rect 17614 2694 17616 2746
rect 17370 2692 17376 2694
rect 17432 2692 17456 2694
rect 17512 2692 17536 2694
rect 17592 2692 17616 2694
rect 17672 2692 17678 2694
rect 17370 2683 17678 2692
rect 17788 2650 17816 3062
rect 20168 3052 20220 3058
rect 20168 2994 20220 3000
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19720 2650 19748 2926
rect 20180 2650 20208 2994
rect 22664 2825 22692 3159
rect 23388 3130 23440 3136
rect 23952 3058 23980 4082
rect 24228 3194 24256 4111
rect 24400 4072 24452 4078
rect 24400 4014 24452 4020
rect 24412 3534 24440 4014
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 25424 3194 25452 5510
rect 25792 5234 25820 7942
rect 25870 7942 26096 7970
rect 25870 7840 25926 7942
rect 25872 5296 25924 5302
rect 25872 5238 25924 5244
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25504 5024 25556 5030
rect 25504 4966 25556 4972
rect 25516 4758 25544 4966
rect 25504 4752 25556 4758
rect 25504 4694 25556 4700
rect 25504 4480 25556 4486
rect 25504 4422 25556 4428
rect 25516 4282 25544 4422
rect 25884 4282 25912 5238
rect 26068 5234 26096 7942
rect 26146 7840 26202 8000
rect 26422 7840 26478 8000
rect 26698 7840 26754 8000
rect 26974 7840 27030 8000
rect 27250 7970 27306 8000
rect 27250 7942 27476 7970
rect 27250 7840 27306 7942
rect 26056 5228 26108 5234
rect 26160 5216 26188 7840
rect 26332 5228 26384 5234
rect 26160 5188 26332 5216
rect 26056 5170 26108 5176
rect 26436 5216 26464 7840
rect 26712 5234 26740 7840
rect 26988 5302 27016 7840
rect 26976 5296 27028 5302
rect 26976 5238 27028 5244
rect 26608 5228 26660 5234
rect 26436 5188 26608 5216
rect 26332 5170 26384 5176
rect 26608 5170 26660 5176
rect 26700 5228 26752 5234
rect 27448 5216 27476 7942
rect 27526 7840 27582 8000
rect 27802 7840 27858 8000
rect 28078 7840 28134 8000
rect 28354 7840 28410 8000
rect 28630 7840 28686 8000
rect 28906 7840 28962 8000
rect 29182 7840 29238 8000
rect 29458 7840 29514 8000
rect 29734 7840 29790 8000
rect 30010 7970 30066 8000
rect 30010 7942 30144 7970
rect 30010 7840 30066 7942
rect 27540 5352 27568 7840
rect 27620 5364 27672 5370
rect 27540 5324 27620 5352
rect 27620 5306 27672 5312
rect 27712 5228 27764 5234
rect 27448 5188 27712 5216
rect 26700 5170 26752 5176
rect 27712 5170 27764 5176
rect 27816 5166 27844 7840
rect 28092 6594 28120 7840
rect 28080 6588 28132 6594
rect 28080 6530 28132 6536
rect 28368 5302 28396 7840
rect 28644 6610 28672 7840
rect 28540 6588 28592 6594
rect 28644 6582 28764 6610
rect 28540 6530 28592 6536
rect 28356 5296 28408 5302
rect 28356 5238 28408 5244
rect 28552 5234 28580 6530
rect 28736 5302 28764 6582
rect 29000 6112 29052 6118
rect 29000 6054 29052 6060
rect 28724 5296 28776 5302
rect 28724 5238 28776 5244
rect 28540 5228 28592 5234
rect 28540 5170 28592 5176
rect 27804 5160 27856 5166
rect 27804 5102 27856 5108
rect 27988 5092 28040 5098
rect 27988 5034 28040 5040
rect 25964 5024 26016 5030
rect 25964 4966 26016 4972
rect 26240 5024 26292 5030
rect 26240 4966 26292 4972
rect 26516 5024 26568 5030
rect 26516 4966 26568 4972
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 26976 5024 27028 5030
rect 26976 4966 27028 4972
rect 27252 5024 27304 5030
rect 27804 5024 27856 5030
rect 27252 4966 27304 4972
rect 27802 4992 27804 5001
rect 27896 5024 27948 5030
rect 27856 4992 27858 5001
rect 25976 4826 26004 4966
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 26252 4690 26280 4966
rect 26332 4752 26384 4758
rect 26332 4694 26384 4700
rect 26240 4684 26292 4690
rect 26240 4626 26292 4632
rect 26252 4282 26280 4626
rect 25504 4276 25556 4282
rect 25504 4218 25556 4224
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 26240 4276 26292 4282
rect 26240 4218 26292 4224
rect 26240 4004 26292 4010
rect 26240 3946 26292 3952
rect 26252 3602 26280 3946
rect 26240 3596 26292 3602
rect 26240 3538 26292 3544
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 25504 3052 25556 3058
rect 25504 2994 25556 3000
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 22650 2816 22706 2825
rect 22650 2751 22706 2760
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 23204 2440 23256 2446
rect 23204 2382 23256 2388
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 16316 1414 16620 1442
rect 16316 160 16344 1414
rect 17052 160 17080 2382
rect 17788 160 17816 2382
rect 18524 160 18552 2382
rect 19260 160 19288 2382
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 20088 2106 20116 2246
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 14830 54 14964 82
rect 12622 0 12678 54
rect 13358 0 13414 54
rect 14094 0 14150 54
rect 14830 0 14886 54
rect 15566 0 15622 160
rect 16302 0 16358 160
rect 17038 0 17094 160
rect 17774 0 17830 160
rect 18510 0 18566 160
rect 19246 0 19302 160
rect 19982 82 20038 160
rect 20272 82 20300 2382
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20824 1902 20852 2246
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 19982 54 20300 82
rect 20718 82 20774 160
rect 21008 82 21036 2382
rect 21468 160 21496 2382
rect 21824 2304 21876 2310
rect 21824 2246 21876 2252
rect 21836 1970 21864 2246
rect 21824 1964 21876 1970
rect 21824 1906 21876 1912
rect 22204 160 22232 2382
rect 22843 2204 23151 2213
rect 22843 2202 22849 2204
rect 22905 2202 22929 2204
rect 22985 2202 23009 2204
rect 23065 2202 23089 2204
rect 23145 2202 23151 2204
rect 22905 2150 22907 2202
rect 23087 2150 23089 2202
rect 22843 2148 22849 2150
rect 22905 2148 22929 2150
rect 22985 2148 23009 2150
rect 23065 2148 23089 2150
rect 23145 2148 23151 2150
rect 22843 2139 23151 2148
rect 20718 54 21036 82
rect 19982 0 20038 54
rect 20718 0 20774 54
rect 21454 0 21510 160
rect 22190 0 22246 160
rect 22926 82 22982 160
rect 23216 82 23244 2382
rect 23676 160 23704 2382
rect 24044 2038 24072 2994
rect 25516 2650 25544 2994
rect 26056 2848 26108 2854
rect 26054 2816 26056 2825
rect 26108 2816 26110 2825
rect 26054 2751 26110 2760
rect 26252 2650 26280 2994
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26344 2514 26372 4694
rect 26528 4010 26556 4966
rect 26712 4078 26740 4966
rect 26700 4072 26752 4078
rect 26700 4014 26752 4020
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26988 3466 27016 4966
rect 27264 3738 27292 4966
rect 27896 4966 27948 4972
rect 27802 4927 27858 4936
rect 27618 4856 27674 4865
rect 27618 4791 27620 4800
rect 27672 4791 27674 4800
rect 27620 4762 27672 4768
rect 27344 4072 27396 4078
rect 27344 4014 27396 4020
rect 27356 3738 27384 4014
rect 27252 3732 27304 3738
rect 27252 3674 27304 3680
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 27908 3398 27936 4966
rect 28000 4672 28028 5034
rect 28264 5024 28316 5030
rect 28184 4984 28264 5012
rect 28184 4826 28212 4984
rect 28264 4966 28316 4972
rect 28724 5024 28776 5030
rect 28724 4966 28776 4972
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 28317 4924 28625 4933
rect 28317 4922 28323 4924
rect 28379 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28625 4924
rect 28379 4870 28381 4922
rect 28561 4870 28563 4922
rect 28317 4868 28323 4870
rect 28379 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28625 4870
rect 28317 4859 28625 4868
rect 28736 4826 28764 4966
rect 28920 4826 28948 4966
rect 29012 4826 29040 6054
rect 30116 5234 30144 7942
rect 30286 7840 30342 8000
rect 30562 7970 30618 8000
rect 30562 7942 30696 7970
rect 30562 7840 30618 7942
rect 30104 5228 30156 5234
rect 30300 5216 30328 7840
rect 30668 5234 30696 7942
rect 30838 7840 30894 8000
rect 31114 7970 31170 8000
rect 31390 7970 31446 8000
rect 31114 7942 31248 7970
rect 31114 7840 31170 7942
rect 30380 5228 30432 5234
rect 30300 5188 30380 5216
rect 30104 5170 30156 5176
rect 30380 5170 30432 5176
rect 30656 5228 30708 5234
rect 30852 5216 30880 7840
rect 31220 5234 31248 7942
rect 31390 7942 31524 7970
rect 31390 7840 31446 7942
rect 31496 5234 31524 7942
rect 31666 7840 31722 8000
rect 31942 7970 31998 8000
rect 31942 7942 32168 7970
rect 31942 7840 31998 7942
rect 30932 5228 30984 5234
rect 30852 5188 30932 5216
rect 30656 5170 30708 5176
rect 30932 5170 30984 5176
rect 31208 5228 31260 5234
rect 31208 5170 31260 5176
rect 31484 5228 31536 5234
rect 31680 5216 31708 7840
rect 32140 5234 32168 7942
rect 32218 7840 32274 8000
rect 32494 7840 32550 8000
rect 32770 7840 32826 8000
rect 33046 7840 33102 8000
rect 33322 7970 33378 8000
rect 33322 7942 33548 7970
rect 33322 7840 33378 7942
rect 31760 5228 31812 5234
rect 31680 5188 31760 5216
rect 31484 5170 31536 5176
rect 31760 5170 31812 5176
rect 32128 5228 32180 5234
rect 32232 5216 32260 7840
rect 32404 5228 32456 5234
rect 32232 5188 32404 5216
rect 32128 5170 32180 5176
rect 32508 5216 32536 7840
rect 32680 5228 32732 5234
rect 32508 5188 32680 5216
rect 32404 5170 32456 5176
rect 32784 5216 32812 7840
rect 33060 5234 33088 7840
rect 33232 6248 33284 6254
rect 33232 6190 33284 6196
rect 32956 5228 33008 5234
rect 32784 5188 32956 5216
rect 32680 5170 32732 5176
rect 32956 5170 33008 5176
rect 33048 5228 33100 5234
rect 33048 5170 33100 5176
rect 33138 5128 33194 5137
rect 31852 5092 31904 5098
rect 31852 5034 31904 5040
rect 32496 5092 32548 5098
rect 32496 5034 32548 5040
rect 33048 5092 33100 5098
rect 33138 5063 33140 5072
rect 33048 5034 33100 5040
rect 33192 5063 33194 5072
rect 33140 5034 33192 5040
rect 30472 5024 30524 5030
rect 30472 4966 30524 4972
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 31116 5024 31168 5030
rect 31116 4966 31168 4972
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 28172 4820 28224 4826
rect 28172 4762 28224 4768
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 28724 4820 28776 4826
rect 28724 4762 28776 4768
rect 28908 4820 28960 4826
rect 28908 4762 28960 4768
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 28460 4729 28488 4762
rect 28446 4720 28502 4729
rect 28000 4644 28120 4672
rect 28446 4655 28502 4664
rect 27988 4548 28040 4554
rect 27988 4490 28040 4496
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27172 2650 27200 2994
rect 27724 2650 27752 2994
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26608 2440 26660 2446
rect 27620 2440 27672 2446
rect 26608 2382 26660 2388
rect 27540 2400 27620 2428
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24032 2032 24084 2038
rect 24032 1974 24084 1980
rect 24504 1834 24532 2246
rect 24492 1828 24544 1834
rect 24492 1770 24544 1776
rect 22926 54 23244 82
rect 22926 0 22982 54
rect 23662 0 23718 160
rect 24398 82 24454 160
rect 24688 82 24716 2382
rect 25148 160 25176 2382
rect 24398 54 24716 82
rect 24398 0 24454 54
rect 25134 0 25190 160
rect 25870 82 25926 160
rect 26160 82 26188 2382
rect 26620 160 26648 2382
rect 25870 54 26188 82
rect 25870 0 25926 54
rect 26606 0 26662 160
rect 27342 82 27398 160
rect 27540 82 27568 2400
rect 27620 2382 27672 2388
rect 28000 1873 28028 4490
rect 28092 4486 28120 4644
rect 28908 4616 28960 4622
rect 28908 4558 28960 4564
rect 29184 4616 29236 4622
rect 29920 4616 29972 4622
rect 29184 4558 29236 4564
rect 29734 4584 29790 4593
rect 28080 4480 28132 4486
rect 28080 4422 28132 4428
rect 28184 3998 28764 4026
rect 28184 3913 28212 3998
rect 28736 3913 28764 3998
rect 28170 3904 28226 3913
rect 28170 3839 28226 3848
rect 28722 3904 28778 3913
rect 28317 3836 28625 3845
rect 28722 3839 28778 3848
rect 28317 3834 28323 3836
rect 28379 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28625 3836
rect 28379 3782 28381 3834
rect 28561 3782 28563 3834
rect 28317 3780 28323 3782
rect 28379 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28625 3782
rect 28317 3771 28625 3780
rect 28317 2748 28625 2757
rect 28317 2746 28323 2748
rect 28379 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28625 2748
rect 28379 2694 28381 2746
rect 28561 2694 28563 2746
rect 28317 2692 28323 2694
rect 28379 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28625 2694
rect 28317 2683 28625 2692
rect 28920 2650 28948 4558
rect 29196 2650 29224 4558
rect 29920 4558 29972 4564
rect 29734 4519 29790 4528
rect 29748 4486 29776 4519
rect 29736 4480 29788 4486
rect 29736 4422 29788 4428
rect 29932 2650 29960 4558
rect 30484 4146 30512 4966
rect 30576 4826 30604 4966
rect 30852 4826 30880 4966
rect 31128 4826 31156 4966
rect 30564 4820 30616 4826
rect 30564 4762 30616 4768
rect 30840 4820 30892 4826
rect 30840 4762 30892 4768
rect 31116 4820 31168 4826
rect 31116 4762 31168 4768
rect 31772 4758 31800 4966
rect 31864 4758 31892 5034
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 32312 5024 32364 5030
rect 32312 4966 32364 4972
rect 31760 4752 31812 4758
rect 31760 4694 31812 4700
rect 31852 4752 31904 4758
rect 31852 4694 31904 4700
rect 31024 4480 31076 4486
rect 31024 4422 31076 4428
rect 31392 4480 31444 4486
rect 31392 4422 31444 4428
rect 31036 4282 31064 4422
rect 31404 4282 31432 4422
rect 31024 4276 31076 4282
rect 31024 4218 31076 4224
rect 31392 4276 31444 4282
rect 31392 4218 31444 4224
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 31484 3392 31536 3398
rect 31484 3334 31536 3340
rect 28908 2644 28960 2650
rect 28908 2586 28960 2592
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29920 2644 29972 2650
rect 29920 2586 29972 2592
rect 31496 2446 31524 3334
rect 31956 3194 31984 4966
rect 32036 4752 32088 4758
rect 32036 4694 32088 4700
rect 31944 3188 31996 3194
rect 31944 3130 31996 3136
rect 32048 2446 32076 4694
rect 32324 3194 32352 4966
rect 32508 3534 32536 5034
rect 32956 4480 33008 4486
rect 32956 4422 33008 4428
rect 32496 3528 32548 3534
rect 32496 3470 32548 3476
rect 32312 3188 32364 3194
rect 32312 3130 32364 3136
rect 32496 2848 32548 2854
rect 32496 2790 32548 2796
rect 32508 2446 32536 2790
rect 32968 2446 32996 4422
rect 33060 3194 33088 5034
rect 33244 4622 33272 6190
rect 33520 5234 33548 7942
rect 33598 7840 33654 8000
rect 33874 7970 33930 8000
rect 34150 7970 34206 8000
rect 33874 7942 34100 7970
rect 33874 7840 33930 7942
rect 33508 5228 33560 5234
rect 33612 5216 33640 7840
rect 34072 7698 34100 7942
rect 34150 7942 34376 7970
rect 34150 7840 34206 7942
rect 34072 7670 34192 7698
rect 33790 5468 34098 5477
rect 33790 5466 33796 5468
rect 33852 5466 33876 5468
rect 33932 5466 33956 5468
rect 34012 5466 34036 5468
rect 34092 5466 34098 5468
rect 33852 5414 33854 5466
rect 34034 5414 34036 5466
rect 33790 5412 33796 5414
rect 33852 5412 33876 5414
rect 33932 5412 33956 5414
rect 34012 5412 34036 5414
rect 34092 5412 34098 5414
rect 33790 5403 34098 5412
rect 33784 5228 33836 5234
rect 33612 5188 33784 5216
rect 33508 5170 33560 5176
rect 34164 5216 34192 7670
rect 34348 5234 34376 7942
rect 34426 7840 34482 8000
rect 34702 7970 34758 8000
rect 34702 7942 34836 7970
rect 34702 7840 34758 7942
rect 34440 5522 34468 7840
rect 34440 5494 34652 5522
rect 34518 5400 34574 5409
rect 34624 5370 34652 5494
rect 34518 5335 34520 5344
rect 34572 5335 34574 5344
rect 34612 5364 34664 5370
rect 34520 5306 34572 5312
rect 34612 5306 34664 5312
rect 34244 5228 34296 5234
rect 34164 5188 34244 5216
rect 33784 5170 33836 5176
rect 34244 5170 34296 5176
rect 34336 5228 34388 5234
rect 34336 5170 34388 5176
rect 34612 5228 34664 5234
rect 34612 5170 34664 5176
rect 33324 5092 33376 5098
rect 33324 5034 33376 5040
rect 34428 5092 34480 5098
rect 34428 5034 34480 5040
rect 33232 4616 33284 4622
rect 33232 4558 33284 4564
rect 33140 3936 33192 3942
rect 33140 3878 33192 3884
rect 33048 3188 33100 3194
rect 33048 3130 33100 3136
rect 33152 2650 33180 3878
rect 33336 2854 33364 5034
rect 33416 5024 33468 5030
rect 33416 4966 33468 4972
rect 33692 5024 33744 5030
rect 33692 4966 33744 4972
rect 34152 5024 34204 5030
rect 34152 4966 34204 4972
rect 33428 3602 33456 4966
rect 33508 4820 33560 4826
rect 33508 4762 33560 4768
rect 33416 3596 33468 3602
rect 33416 3538 33468 3544
rect 33324 2848 33376 2854
rect 33324 2790 33376 2796
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33520 2446 33548 4762
rect 33704 4078 33732 4966
rect 33790 4380 34098 4389
rect 33790 4378 33796 4380
rect 33852 4378 33876 4380
rect 33932 4378 33956 4380
rect 34012 4378 34036 4380
rect 34092 4378 34098 4380
rect 33852 4326 33854 4378
rect 34034 4326 34036 4378
rect 33790 4324 33796 4326
rect 33852 4324 33876 4326
rect 33932 4324 33956 4326
rect 34012 4324 34036 4326
rect 34092 4324 34098 4326
rect 33790 4315 34098 4324
rect 33692 4072 33744 4078
rect 33692 4014 33744 4020
rect 34164 3534 34192 4966
rect 34440 4826 34468 5034
rect 34428 4820 34480 4826
rect 34428 4762 34480 4768
rect 34428 4616 34480 4622
rect 34428 4558 34480 4564
rect 34336 4208 34388 4214
rect 34336 4150 34388 4156
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34152 3528 34204 3534
rect 34152 3470 34204 3476
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 29828 2440 29880 2446
rect 29828 2382 29880 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 31484 2440 31536 2446
rect 31484 2382 31536 2388
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 27986 1864 28042 1873
rect 27986 1799 28042 1808
rect 28092 160 28120 2382
rect 28828 160 28856 2382
rect 27342 54 27568 82
rect 27342 0 27398 54
rect 28078 0 28134 160
rect 28814 0 28870 160
rect 29550 82 29606 160
rect 29840 82 29868 2382
rect 30300 160 30328 2382
rect 31116 2372 31168 2378
rect 31116 2314 31168 2320
rect 32128 2372 32180 2378
rect 32128 2314 32180 2320
rect 29550 54 29868 82
rect 29550 0 29606 54
rect 30286 0 30342 160
rect 31022 82 31078 160
rect 31128 82 31156 2314
rect 31022 54 31156 82
rect 31758 82 31814 160
rect 32140 82 32168 2314
rect 32496 2304 32548 2310
rect 32496 2246 32548 2252
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 32508 160 32536 2246
rect 31758 54 32168 82
rect 31022 0 31078 54
rect 31758 0 31814 54
rect 32494 0 32550 160
rect 33230 82 33286 160
rect 33520 82 33548 2246
rect 33612 1358 33640 3470
rect 34244 3460 34296 3466
rect 34244 3402 34296 3408
rect 33790 3292 34098 3301
rect 33790 3290 33796 3292
rect 33852 3290 33876 3292
rect 33932 3290 33956 3292
rect 34012 3290 34036 3292
rect 34092 3290 34098 3292
rect 33852 3238 33854 3290
rect 34034 3238 34036 3290
rect 33790 3236 33796 3238
rect 33852 3236 33876 3238
rect 33932 3236 33956 3238
rect 34012 3236 34036 3238
rect 34092 3236 34098 3238
rect 33790 3227 34098 3236
rect 34256 2446 34284 3402
rect 34348 2446 34376 4150
rect 34244 2440 34296 2446
rect 34244 2382 34296 2388
rect 34336 2440 34388 2446
rect 34336 2382 34388 2388
rect 34244 2304 34296 2310
rect 34244 2246 34296 2252
rect 33790 2204 34098 2213
rect 33790 2202 33796 2204
rect 33852 2202 33876 2204
rect 33932 2202 33956 2204
rect 34012 2202 34036 2204
rect 34092 2202 34098 2204
rect 33852 2150 33854 2202
rect 34034 2150 34036 2202
rect 33790 2148 33796 2150
rect 33852 2148 33876 2150
rect 33932 2148 33956 2150
rect 34012 2148 34036 2150
rect 34092 2148 34098 2150
rect 33790 2139 34098 2148
rect 33600 1352 33652 1358
rect 33600 1294 33652 1300
rect 33230 54 33548 82
rect 33966 82 34022 160
rect 34256 82 34284 2246
rect 34440 2009 34468 4558
rect 34520 4276 34572 4282
rect 34520 4218 34572 4224
rect 34532 2446 34560 4218
rect 34624 3738 34652 5170
rect 34808 4826 34836 7942
rect 34978 7840 35034 8000
rect 35254 7970 35310 8000
rect 35530 7970 35586 8000
rect 35254 7942 35480 7970
rect 35254 7840 35310 7942
rect 34992 5370 35020 7840
rect 35452 7698 35480 7942
rect 35530 7942 35756 7970
rect 35530 7840 35586 7942
rect 35452 7670 35572 7698
rect 35164 6316 35216 6322
rect 35164 6258 35216 6264
rect 35072 6180 35124 6186
rect 35072 6122 35124 6128
rect 34980 5364 35032 5370
rect 34980 5306 35032 5312
rect 34796 4820 34848 4826
rect 34796 4762 34848 4768
rect 35084 4622 35112 6122
rect 35176 4622 35204 6258
rect 35544 5370 35572 7670
rect 35532 5364 35584 5370
rect 35532 5306 35584 5312
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 35256 5160 35308 5166
rect 35256 5102 35308 5108
rect 35268 4826 35296 5102
rect 35360 4826 35388 5170
rect 35532 5160 35584 5166
rect 35532 5102 35584 5108
rect 35256 4820 35308 4826
rect 35256 4762 35308 4768
rect 35348 4820 35400 4826
rect 35348 4762 35400 4768
rect 35072 4616 35124 4622
rect 35072 4558 35124 4564
rect 35164 4616 35216 4622
rect 35164 4558 35216 4564
rect 34612 3732 34664 3738
rect 34612 3674 34664 3680
rect 34796 3052 34848 3058
rect 34796 2994 34848 3000
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 34426 2000 34482 2009
rect 34426 1935 34482 1944
rect 34808 1290 34836 2994
rect 35544 2854 35572 5102
rect 35728 5030 35756 7942
rect 35806 7840 35862 8000
rect 36082 7840 36138 8000
rect 36358 7970 36414 8000
rect 36358 7942 36584 7970
rect 36358 7840 36414 7942
rect 35716 5024 35768 5030
rect 35716 4966 35768 4972
rect 35820 4826 35848 7840
rect 36096 6202 36124 7840
rect 36096 6174 36216 6202
rect 35808 4820 35860 4826
rect 35808 4762 35860 4768
rect 36188 4758 36216 6174
rect 36556 5370 36584 7942
rect 36634 7840 36690 8000
rect 36910 7840 36966 8000
rect 37186 7840 37242 8000
rect 37462 7970 37518 8000
rect 37462 7942 37688 7970
rect 37462 7840 37518 7942
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36648 4826 36676 7840
rect 36728 5228 36780 5234
rect 36728 5170 36780 5176
rect 36636 4820 36688 4826
rect 36636 4762 36688 4768
rect 36176 4752 36228 4758
rect 36176 4694 36228 4700
rect 35624 4616 35676 4622
rect 35624 4558 35676 4564
rect 35532 2848 35584 2854
rect 35532 2790 35584 2796
rect 35636 2689 35664 4558
rect 36740 4214 36768 5170
rect 36924 5030 36952 7840
rect 37200 5522 37228 7840
rect 37200 5494 37320 5522
rect 37188 5160 37240 5166
rect 37188 5102 37240 5108
rect 36912 5024 36964 5030
rect 36912 4966 36964 4972
rect 37096 4548 37148 4554
rect 37096 4490 37148 4496
rect 37108 4282 37136 4490
rect 37096 4276 37148 4282
rect 37096 4218 37148 4224
rect 36728 4208 36780 4214
rect 36728 4150 36780 4156
rect 35716 4140 35768 4146
rect 35716 4082 35768 4088
rect 35992 4140 36044 4146
rect 35992 4082 36044 4088
rect 36268 4140 36320 4146
rect 36268 4082 36320 4088
rect 36544 4140 36596 4146
rect 36544 4082 36596 4088
rect 35622 2680 35678 2689
rect 35622 2615 35678 2624
rect 34980 2304 35032 2310
rect 34980 2246 35032 2252
rect 34796 1284 34848 1290
rect 34796 1226 34848 1232
rect 33966 54 34284 82
rect 34702 82 34758 160
rect 34992 82 35020 2246
rect 35728 1222 35756 4082
rect 36004 2417 36032 4082
rect 36084 4004 36136 4010
rect 36084 3946 36136 3952
rect 36096 2446 36124 3946
rect 36084 2440 36136 2446
rect 35990 2408 36046 2417
rect 36084 2382 36136 2388
rect 35990 2343 36046 2352
rect 35900 2304 35952 2310
rect 35900 2246 35952 2252
rect 35912 1442 35940 2246
rect 36280 1737 36308 4082
rect 36556 3738 36584 4082
rect 37200 4010 37228 5102
rect 37292 4758 37320 5494
rect 37660 5098 37688 7942
rect 37738 7840 37794 8000
rect 38014 7970 38070 8000
rect 38014 7942 38240 7970
rect 38014 7840 38070 7942
rect 37648 5092 37700 5098
rect 37648 5034 37700 5040
rect 37752 4826 37780 7840
rect 38212 5370 38240 7942
rect 38290 7840 38346 8000
rect 38566 7840 38622 8000
rect 38842 7970 38898 8000
rect 38842 7942 39068 7970
rect 38842 7840 38898 7942
rect 38200 5364 38252 5370
rect 38200 5306 38252 5312
rect 38016 5160 38068 5166
rect 38016 5102 38068 5108
rect 37740 4820 37792 4826
rect 37740 4762 37792 4768
rect 37280 4752 37332 4758
rect 37280 4694 37332 4700
rect 37648 4548 37700 4554
rect 37648 4490 37700 4496
rect 37740 4548 37792 4554
rect 37740 4490 37792 4496
rect 37660 4185 37688 4490
rect 37646 4176 37702 4185
rect 37646 4111 37702 4120
rect 37188 4004 37240 4010
rect 37188 3946 37240 3952
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 37292 2446 37320 3878
rect 37752 3097 37780 4490
rect 37738 3088 37794 3097
rect 37738 3023 37794 3032
rect 38028 2961 38056 5102
rect 38304 4808 38332 7840
rect 38384 4820 38436 4826
rect 38304 4780 38384 4808
rect 38384 4762 38436 4768
rect 38580 4758 38608 7840
rect 38660 5772 38712 5778
rect 38660 5714 38712 5720
rect 38672 5302 38700 5714
rect 38660 5296 38712 5302
rect 38660 5238 38712 5244
rect 39040 5012 39068 7942
rect 39118 7840 39174 8000
rect 39394 7970 39450 8000
rect 39670 7970 39726 8000
rect 39394 7942 39620 7970
rect 39394 7840 39450 7942
rect 39132 5250 39160 7840
rect 39592 7698 39620 7942
rect 39670 7942 39896 7970
rect 39670 7840 39726 7942
rect 39592 7670 39712 7698
rect 39684 5370 39712 7670
rect 39672 5364 39724 5370
rect 39672 5306 39724 5312
rect 39132 5222 39712 5250
rect 39304 5024 39356 5030
rect 39040 4984 39304 5012
rect 39304 4966 39356 4972
rect 39264 4924 39572 4933
rect 39264 4922 39270 4924
rect 39326 4922 39350 4924
rect 39406 4922 39430 4924
rect 39486 4922 39510 4924
rect 39566 4922 39572 4924
rect 39326 4870 39328 4922
rect 39508 4870 39510 4922
rect 39264 4868 39270 4870
rect 39326 4868 39350 4870
rect 39406 4868 39430 4870
rect 39486 4868 39510 4870
rect 39566 4868 39572 4870
rect 39264 4859 39572 4868
rect 39684 4826 39712 5222
rect 39672 4820 39724 4826
rect 39672 4762 39724 4768
rect 38568 4752 38620 4758
rect 38568 4694 38620 4700
rect 39868 4706 39896 7942
rect 39946 7840 40002 8000
rect 40222 7840 40278 8000
rect 39960 5522 39988 7840
rect 39960 5494 40080 5522
rect 40052 5302 40080 5494
rect 40130 5400 40186 5409
rect 40130 5335 40186 5344
rect 40040 5296 40092 5302
rect 40040 5238 40092 5244
rect 39948 4752 40000 4758
rect 39868 4700 39948 4706
rect 39868 4694 40000 4700
rect 39868 4678 39988 4694
rect 40144 4690 40172 5335
rect 40236 4826 40264 7840
rect 40316 5908 40368 5914
rect 40316 5850 40368 5856
rect 40224 4820 40276 4826
rect 40224 4762 40276 4768
rect 40132 4684 40184 4690
rect 40132 4626 40184 4632
rect 40328 4622 40356 5850
rect 40592 5840 40644 5846
rect 40592 5782 40644 5788
rect 40604 5234 40632 5782
rect 44737 5468 45045 5477
rect 44737 5466 44743 5468
rect 44799 5466 44823 5468
rect 44879 5466 44903 5468
rect 44959 5466 44983 5468
rect 45039 5466 45045 5468
rect 44799 5414 44801 5466
rect 44981 5414 44983 5466
rect 44737 5412 44743 5414
rect 44799 5412 44823 5414
rect 44879 5412 44903 5414
rect 44959 5412 44983 5414
rect 45039 5412 45045 5414
rect 44737 5403 45045 5412
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40592 5228 40644 5234
rect 40592 5170 40644 5176
rect 40316 4616 40368 4622
rect 40316 4558 40368 4564
rect 39304 4548 39356 4554
rect 39304 4490 39356 4496
rect 39948 4548 40000 4554
rect 39948 4490 40000 4496
rect 38660 4480 38712 4486
rect 38660 4422 38712 4428
rect 38200 4004 38252 4010
rect 38200 3946 38252 3952
rect 38212 3738 38240 3946
rect 38200 3732 38252 3738
rect 38200 3674 38252 3680
rect 38672 3505 38700 4422
rect 39120 4140 39172 4146
rect 39120 4082 39172 4088
rect 39132 3738 39160 4082
rect 39316 4049 39344 4490
rect 39302 4040 39358 4049
rect 39302 3975 39358 3984
rect 39672 3936 39724 3942
rect 39672 3878 39724 3884
rect 39264 3836 39572 3845
rect 39264 3834 39270 3836
rect 39326 3834 39350 3836
rect 39406 3834 39430 3836
rect 39486 3834 39510 3836
rect 39566 3834 39572 3836
rect 39326 3782 39328 3834
rect 39508 3782 39510 3834
rect 39264 3780 39270 3782
rect 39326 3780 39350 3782
rect 39406 3780 39430 3782
rect 39486 3780 39510 3782
rect 39566 3780 39572 3782
rect 39264 3771 39572 3780
rect 39120 3732 39172 3738
rect 39120 3674 39172 3680
rect 38658 3496 38714 3505
rect 38658 3431 38714 3440
rect 38014 2952 38070 2961
rect 38014 2887 38070 2896
rect 39264 2748 39572 2757
rect 39264 2746 39270 2748
rect 39326 2746 39350 2748
rect 39406 2746 39430 2748
rect 39486 2746 39510 2748
rect 39566 2746 39572 2748
rect 39326 2694 39328 2746
rect 39508 2694 39510 2746
rect 39264 2692 39270 2694
rect 39326 2692 39350 2694
rect 39406 2692 39430 2694
rect 39486 2692 39510 2694
rect 39566 2692 39572 2694
rect 39264 2683 39572 2692
rect 39684 2446 39712 3878
rect 39960 3641 39988 4490
rect 40512 4321 40540 5170
rect 41510 5128 41566 5137
rect 41510 5063 41566 5072
rect 41524 4622 41552 5063
rect 41512 4616 41564 4622
rect 41512 4558 41564 4564
rect 41696 4480 41748 4486
rect 41696 4422 41748 4428
rect 42708 4480 42760 4486
rect 42708 4422 42760 4428
rect 40498 4312 40554 4321
rect 40498 4247 40554 4256
rect 40408 3936 40460 3942
rect 40408 3878 40460 3884
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 39946 3632 40002 3641
rect 39946 3567 40002 3576
rect 40420 2446 40448 3878
rect 41432 2446 41460 3878
rect 41708 2446 41736 4422
rect 42720 2446 42748 4422
rect 44737 4380 45045 4389
rect 44737 4378 44743 4380
rect 44799 4378 44823 4380
rect 44879 4378 44903 4380
rect 44959 4378 44983 4380
rect 45039 4378 45045 4380
rect 44799 4326 44801 4378
rect 44981 4326 44983 4378
rect 44737 4324 44743 4326
rect 44799 4324 44823 4326
rect 44879 4324 44903 4326
rect 44959 4324 44983 4326
rect 45039 4324 45045 4326
rect 44737 4315 45045 4324
rect 44737 3292 45045 3301
rect 44737 3290 44743 3292
rect 44799 3290 44823 3292
rect 44879 3290 44903 3292
rect 44959 3290 44983 3292
rect 45039 3290 45045 3292
rect 44799 3238 44801 3290
rect 44981 3238 44983 3290
rect 44737 3236 44743 3238
rect 44799 3236 44823 3238
rect 44879 3236 44903 3238
rect 44959 3236 44983 3238
rect 45039 3236 45045 3238
rect 44737 3227 45045 3236
rect 43168 3188 43220 3194
rect 43168 3130 43220 3136
rect 43180 2446 43208 3130
rect 44640 2916 44692 2922
rect 44640 2858 44692 2864
rect 44272 2848 44324 2854
rect 44272 2790 44324 2796
rect 37280 2440 37332 2446
rect 37280 2382 37332 2388
rect 39672 2440 39724 2446
rect 39672 2382 39724 2388
rect 40408 2440 40460 2446
rect 40408 2382 40460 2388
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 41696 2440 41748 2446
rect 41696 2382 41748 2388
rect 42708 2440 42760 2446
rect 42708 2382 42760 2388
rect 43168 2440 43220 2446
rect 43168 2382 43220 2388
rect 36452 2304 36504 2310
rect 36452 2246 36504 2252
rect 37188 2304 37240 2310
rect 37188 2246 37240 2252
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38384 2304 38436 2310
rect 38384 2246 38436 2252
rect 39396 2304 39448 2310
rect 39396 2246 39448 2252
rect 39856 2304 39908 2310
rect 39856 2246 39908 2252
rect 40868 2304 40920 2310
rect 40868 2246 40920 2252
rect 41328 2304 41380 2310
rect 41328 2246 41380 2252
rect 42432 2304 42484 2310
rect 42432 2246 42484 2252
rect 43168 2304 43220 2310
rect 43168 2246 43220 2252
rect 43812 2304 43864 2310
rect 43812 2246 43864 2252
rect 36266 1728 36322 1737
rect 36266 1663 36322 1672
rect 35820 1414 35940 1442
rect 35716 1216 35768 1222
rect 35716 1158 35768 1164
rect 34702 54 35020 82
rect 35438 82 35494 160
rect 35820 82 35848 1414
rect 35438 54 35848 82
rect 36174 82 36230 160
rect 36464 82 36492 2246
rect 36174 54 36492 82
rect 36910 82 36966 160
rect 37200 82 37228 2246
rect 36910 54 37228 82
rect 37646 82 37702 160
rect 38028 82 38056 2246
rect 38396 160 38424 2246
rect 37646 54 38056 82
rect 33230 0 33286 54
rect 33966 0 34022 54
rect 34702 0 34758 54
rect 35438 0 35494 54
rect 36174 0 36230 54
rect 36910 0 36966 54
rect 37646 0 37702 54
rect 38382 0 38438 160
rect 39118 82 39174 160
rect 39408 82 39436 2246
rect 39868 160 39896 2246
rect 39118 54 39436 82
rect 39118 0 39174 54
rect 39854 0 39910 160
rect 40590 82 40646 160
rect 40880 82 40908 2246
rect 41340 160 41368 2246
rect 42076 190 42196 218
rect 42076 160 42104 190
rect 40590 54 40908 82
rect 40590 0 40646 54
rect 41326 0 41382 160
rect 42062 0 42118 160
rect 42168 82 42196 190
rect 42444 82 42472 2246
rect 42168 54 42472 82
rect 42798 82 42854 160
rect 43180 82 43208 2246
rect 42798 54 43208 82
rect 43534 82 43590 160
rect 43824 82 43852 2246
rect 44284 160 44312 2790
rect 43534 54 43852 82
rect 42798 0 42854 54
rect 43534 0 43590 54
rect 44270 0 44326 160
rect 44652 82 44680 2858
rect 44737 2204 45045 2213
rect 44737 2202 44743 2204
rect 44799 2202 44823 2204
rect 44879 2202 44903 2204
rect 44959 2202 44983 2204
rect 45039 2202 45045 2204
rect 44799 2150 44801 2202
rect 44981 2150 44983 2202
rect 44737 2148 44743 2150
rect 44799 2148 44823 2150
rect 44879 2148 44903 2150
rect 44959 2148 44983 2150
rect 45039 2148 45045 2150
rect 44737 2139 45045 2148
rect 45006 82 45062 160
rect 44652 54 45062 82
rect 45006 0 45062 54
<< via2 >>
rect 6182 5752 6238 5808
rect 6734 5616 6790 5672
rect 6429 4922 6485 4924
rect 6509 4922 6565 4924
rect 6589 4922 6645 4924
rect 6669 4922 6725 4924
rect 6429 4870 6475 4922
rect 6475 4870 6485 4922
rect 6509 4870 6539 4922
rect 6539 4870 6551 4922
rect 6551 4870 6565 4922
rect 6589 4870 6603 4922
rect 6603 4870 6615 4922
rect 6615 4870 6645 4922
rect 6669 4870 6679 4922
rect 6679 4870 6725 4922
rect 6429 4868 6485 4870
rect 6509 4868 6565 4870
rect 6589 4868 6645 4870
rect 6669 4868 6725 4870
rect 7010 5228 7066 5264
rect 7010 5208 7012 5228
rect 7012 5208 7064 5228
rect 7064 5208 7066 5228
rect 9402 4392 9458 4448
rect 11242 4664 11298 4720
rect 11902 5466 11958 5468
rect 11982 5466 12038 5468
rect 12062 5466 12118 5468
rect 12142 5466 12198 5468
rect 11902 5414 11948 5466
rect 11948 5414 11958 5466
rect 11982 5414 12012 5466
rect 12012 5414 12024 5466
rect 12024 5414 12038 5466
rect 12062 5414 12076 5466
rect 12076 5414 12088 5466
rect 12088 5414 12118 5466
rect 12142 5414 12152 5466
rect 12152 5414 12198 5466
rect 11902 5412 11958 5414
rect 11982 5412 12038 5414
rect 12062 5412 12118 5414
rect 12142 5412 12198 5414
rect 11886 4972 11888 4992
rect 11888 4972 11940 4992
rect 11940 4972 11942 4992
rect 11886 4936 11942 4972
rect 11702 4800 11758 4856
rect 12346 4664 12402 4720
rect 11902 4378 11958 4380
rect 11982 4378 12038 4380
rect 12062 4378 12118 4380
rect 12142 4378 12198 4380
rect 11902 4326 11948 4378
rect 11948 4326 11958 4378
rect 11982 4326 12012 4378
rect 12012 4326 12024 4378
rect 12024 4326 12038 4378
rect 12062 4326 12076 4378
rect 12076 4326 12088 4378
rect 12088 4326 12118 4378
rect 12142 4326 12152 4378
rect 12152 4326 12198 4378
rect 11902 4324 11958 4326
rect 11982 4324 12038 4326
rect 12062 4324 12118 4326
rect 12142 4324 12198 4326
rect 11242 4156 11244 4176
rect 11244 4156 11296 4176
rect 11296 4156 11298 4176
rect 11242 4120 11298 4156
rect 6429 3834 6485 3836
rect 6509 3834 6565 3836
rect 6589 3834 6645 3836
rect 6669 3834 6725 3836
rect 6429 3782 6475 3834
rect 6475 3782 6485 3834
rect 6509 3782 6539 3834
rect 6539 3782 6551 3834
rect 6551 3782 6565 3834
rect 6589 3782 6603 3834
rect 6603 3782 6615 3834
rect 6615 3782 6645 3834
rect 6669 3782 6679 3834
rect 6679 3782 6725 3834
rect 6429 3780 6485 3782
rect 6509 3780 6565 3782
rect 6589 3780 6645 3782
rect 6669 3780 6725 3782
rect 11242 3052 11298 3088
rect 11242 3032 11244 3052
rect 11244 3032 11296 3052
rect 11296 3032 11298 3052
rect 4710 2508 4766 2544
rect 4710 2488 4712 2508
rect 4712 2488 4764 2508
rect 4764 2488 4766 2508
rect 6429 2746 6485 2748
rect 6509 2746 6565 2748
rect 6589 2746 6645 2748
rect 6669 2746 6725 2748
rect 6429 2694 6475 2746
rect 6475 2694 6485 2746
rect 6509 2694 6539 2746
rect 6539 2694 6551 2746
rect 6551 2694 6565 2746
rect 6589 2694 6603 2746
rect 6603 2694 6615 2746
rect 6615 2694 6645 2746
rect 6669 2694 6679 2746
rect 6679 2694 6725 2746
rect 6429 2692 6485 2694
rect 6509 2692 6565 2694
rect 6589 2692 6645 2694
rect 6669 2692 6725 2694
rect 10506 2916 10562 2952
rect 10506 2896 10508 2916
rect 10508 2896 10560 2916
rect 10560 2896 10562 2916
rect 12438 4256 12494 4312
rect 11978 3576 12034 3632
rect 11902 3290 11958 3292
rect 11982 3290 12038 3292
rect 12062 3290 12118 3292
rect 12142 3290 12198 3292
rect 11902 3238 11948 3290
rect 11948 3238 11958 3290
rect 11982 3238 12012 3290
rect 12012 3238 12024 3290
rect 12024 3238 12038 3290
rect 12062 3238 12076 3290
rect 12076 3238 12088 3290
rect 12088 3238 12118 3290
rect 12142 3238 12152 3290
rect 12152 3238 12198 3290
rect 11902 3236 11958 3238
rect 11982 3236 12038 3238
rect 12062 3236 12118 3238
rect 12142 3236 12198 3238
rect 5906 2388 5908 2408
rect 5908 2388 5960 2408
rect 5960 2388 5962 2408
rect 5906 2352 5962 2388
rect 7102 1672 7158 1728
rect 8482 1944 8538 2000
rect 9218 1808 9274 1864
rect 11902 2202 11958 2204
rect 11982 2202 12038 2204
rect 12062 2202 12118 2204
rect 12142 2202 12198 2204
rect 11902 2150 11948 2202
rect 11948 2150 11958 2202
rect 11982 2150 12012 2202
rect 12012 2150 12024 2202
rect 12024 2150 12038 2202
rect 12062 2150 12076 2202
rect 12076 2150 12088 2202
rect 12088 2150 12118 2202
rect 12142 2150 12152 2202
rect 12152 2150 12198 2202
rect 11902 2148 11958 2150
rect 11982 2148 12038 2150
rect 12062 2148 12118 2150
rect 12142 2148 12198 2150
rect 13266 4548 13322 4584
rect 13266 4528 13268 4548
rect 13268 4528 13320 4548
rect 13320 4528 13322 4548
rect 13450 3576 13506 3632
rect 14186 3848 14242 3904
rect 15106 5072 15162 5128
rect 15106 4684 15162 4720
rect 15106 4664 15108 4684
rect 15108 4664 15160 4684
rect 15160 4664 15162 4684
rect 14554 3440 14610 3496
rect 15198 3168 15254 3224
rect 16026 4936 16082 4992
rect 16578 4800 16634 4856
rect 17376 4922 17432 4924
rect 17456 4922 17512 4924
rect 17536 4922 17592 4924
rect 17616 4922 17672 4924
rect 17376 4870 17422 4922
rect 17422 4870 17432 4922
rect 17456 4870 17486 4922
rect 17486 4870 17498 4922
rect 17498 4870 17512 4922
rect 17536 4870 17550 4922
rect 17550 4870 17562 4922
rect 17562 4870 17592 4922
rect 17616 4870 17626 4922
rect 17626 4870 17672 4922
rect 17376 4868 17432 4870
rect 17456 4868 17512 4870
rect 17536 4868 17592 4870
rect 17616 4868 17672 4870
rect 19338 5752 19394 5808
rect 19614 5616 19670 5672
rect 19522 4936 19578 4992
rect 19798 5344 19854 5400
rect 19890 4800 19946 4856
rect 17376 3834 17432 3836
rect 17456 3834 17512 3836
rect 17536 3834 17592 3836
rect 17616 3834 17672 3836
rect 17376 3782 17422 3834
rect 17422 3782 17432 3834
rect 17456 3782 17486 3834
rect 17486 3782 17498 3834
rect 17498 3782 17512 3834
rect 17536 3782 17550 3834
rect 17550 3782 17562 3834
rect 17562 3782 17592 3834
rect 17616 3782 17626 3834
rect 17626 3782 17672 3834
rect 17376 3780 17432 3782
rect 17456 3780 17512 3782
rect 17536 3780 17592 3782
rect 17616 3780 17672 3782
rect 18234 3984 18290 4040
rect 18234 3304 18290 3360
rect 20442 5344 20498 5400
rect 21454 4800 21510 4856
rect 22849 5466 22905 5468
rect 22929 5466 22985 5468
rect 23009 5466 23065 5468
rect 23089 5466 23145 5468
rect 22849 5414 22895 5466
rect 22895 5414 22905 5466
rect 22929 5414 22959 5466
rect 22959 5414 22971 5466
rect 22971 5414 22985 5466
rect 23009 5414 23023 5466
rect 23023 5414 23035 5466
rect 23035 5414 23065 5466
rect 23089 5414 23099 5466
rect 23099 5414 23145 5466
rect 22849 5412 22905 5414
rect 22929 5412 22985 5414
rect 23009 5412 23065 5414
rect 23089 5412 23145 5414
rect 22006 4800 22062 4856
rect 22190 4800 22246 4856
rect 23386 5072 23442 5128
rect 23018 4800 23074 4856
rect 22282 4428 22284 4448
rect 22284 4428 22336 4448
rect 22336 4428 22338 4448
rect 22282 4392 22338 4428
rect 22650 4256 22706 4312
rect 22849 4378 22905 4380
rect 22929 4378 22985 4380
rect 23009 4378 23065 4380
rect 23089 4378 23145 4380
rect 22849 4326 22895 4378
rect 22895 4326 22905 4378
rect 22929 4326 22959 4378
rect 22959 4326 22971 4378
rect 22971 4326 22985 4378
rect 23009 4326 23023 4378
rect 23023 4326 23035 4378
rect 23035 4326 23065 4378
rect 23089 4326 23099 4378
rect 23099 4326 23145 4378
rect 22849 4324 22905 4326
rect 22929 4324 22985 4326
rect 23009 4324 23065 4326
rect 23089 4324 23145 4326
rect 22742 4120 22798 4176
rect 22849 3290 22905 3292
rect 22929 3290 22985 3292
rect 23009 3290 23065 3292
rect 23089 3290 23145 3292
rect 22849 3238 22895 3290
rect 22895 3238 22905 3290
rect 22929 3238 22959 3290
rect 22959 3238 22971 3290
rect 22971 3238 22985 3290
rect 23009 3238 23023 3290
rect 23023 3238 23035 3290
rect 23035 3238 23065 3290
rect 23089 3238 23099 3290
rect 23099 3238 23145 3290
rect 22849 3236 22905 3238
rect 22929 3236 22985 3238
rect 23009 3236 23065 3238
rect 23089 3236 23145 3238
rect 22650 3168 22706 3224
rect 24398 5208 24454 5264
rect 24214 4120 24270 4176
rect 17376 2746 17432 2748
rect 17456 2746 17512 2748
rect 17536 2746 17592 2748
rect 17616 2746 17672 2748
rect 17376 2694 17422 2746
rect 17422 2694 17432 2746
rect 17456 2694 17486 2746
rect 17486 2694 17498 2746
rect 17498 2694 17512 2746
rect 17536 2694 17550 2746
rect 17550 2694 17562 2746
rect 17562 2694 17592 2746
rect 17616 2694 17626 2746
rect 17626 2694 17672 2746
rect 17376 2692 17432 2694
rect 17456 2692 17512 2694
rect 17536 2692 17592 2694
rect 17616 2692 17672 2694
rect 27802 4972 27804 4992
rect 27804 4972 27856 4992
rect 27856 4972 27858 4992
rect 22650 2760 22706 2816
rect 22849 2202 22905 2204
rect 22929 2202 22985 2204
rect 23009 2202 23065 2204
rect 23089 2202 23145 2204
rect 22849 2150 22895 2202
rect 22895 2150 22905 2202
rect 22929 2150 22959 2202
rect 22959 2150 22971 2202
rect 22971 2150 22985 2202
rect 23009 2150 23023 2202
rect 23023 2150 23035 2202
rect 23035 2150 23065 2202
rect 23089 2150 23099 2202
rect 23099 2150 23145 2202
rect 22849 2148 22905 2150
rect 22929 2148 22985 2150
rect 23009 2148 23065 2150
rect 23089 2148 23145 2150
rect 26054 2796 26056 2816
rect 26056 2796 26108 2816
rect 26108 2796 26110 2816
rect 26054 2760 26110 2796
rect 27802 4936 27858 4972
rect 27618 4820 27674 4856
rect 27618 4800 27620 4820
rect 27620 4800 27672 4820
rect 27672 4800 27674 4820
rect 28323 4922 28379 4924
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28323 4870 28369 4922
rect 28369 4870 28379 4922
rect 28403 4870 28433 4922
rect 28433 4870 28445 4922
rect 28445 4870 28459 4922
rect 28483 4870 28497 4922
rect 28497 4870 28509 4922
rect 28509 4870 28539 4922
rect 28563 4870 28573 4922
rect 28573 4870 28619 4922
rect 28323 4868 28379 4870
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 33138 5092 33194 5128
rect 33138 5072 33140 5092
rect 33140 5072 33192 5092
rect 33192 5072 33194 5092
rect 28446 4664 28502 4720
rect 28170 3848 28226 3904
rect 28722 3848 28778 3904
rect 28323 3834 28379 3836
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28323 3782 28369 3834
rect 28369 3782 28379 3834
rect 28403 3782 28433 3834
rect 28433 3782 28445 3834
rect 28445 3782 28459 3834
rect 28483 3782 28497 3834
rect 28497 3782 28509 3834
rect 28509 3782 28539 3834
rect 28563 3782 28573 3834
rect 28573 3782 28619 3834
rect 28323 3780 28379 3782
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28323 2746 28379 2748
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28323 2694 28369 2746
rect 28369 2694 28379 2746
rect 28403 2694 28433 2746
rect 28433 2694 28445 2746
rect 28445 2694 28459 2746
rect 28483 2694 28497 2746
rect 28497 2694 28509 2746
rect 28509 2694 28539 2746
rect 28563 2694 28573 2746
rect 28573 2694 28619 2746
rect 28323 2692 28379 2694
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 29734 4528 29790 4584
rect 33796 5466 33852 5468
rect 33876 5466 33932 5468
rect 33956 5466 34012 5468
rect 34036 5466 34092 5468
rect 33796 5414 33842 5466
rect 33842 5414 33852 5466
rect 33876 5414 33906 5466
rect 33906 5414 33918 5466
rect 33918 5414 33932 5466
rect 33956 5414 33970 5466
rect 33970 5414 33982 5466
rect 33982 5414 34012 5466
rect 34036 5414 34046 5466
rect 34046 5414 34092 5466
rect 33796 5412 33852 5414
rect 33876 5412 33932 5414
rect 33956 5412 34012 5414
rect 34036 5412 34092 5414
rect 34518 5364 34574 5400
rect 34518 5344 34520 5364
rect 34520 5344 34572 5364
rect 34572 5344 34574 5364
rect 33796 4378 33852 4380
rect 33876 4378 33932 4380
rect 33956 4378 34012 4380
rect 34036 4378 34092 4380
rect 33796 4326 33842 4378
rect 33842 4326 33852 4378
rect 33876 4326 33906 4378
rect 33906 4326 33918 4378
rect 33918 4326 33932 4378
rect 33956 4326 33970 4378
rect 33970 4326 33982 4378
rect 33982 4326 34012 4378
rect 34036 4326 34046 4378
rect 34046 4326 34092 4378
rect 33796 4324 33852 4326
rect 33876 4324 33932 4326
rect 33956 4324 34012 4326
rect 34036 4324 34092 4326
rect 27986 1808 28042 1864
rect 33796 3290 33852 3292
rect 33876 3290 33932 3292
rect 33956 3290 34012 3292
rect 34036 3290 34092 3292
rect 33796 3238 33842 3290
rect 33842 3238 33852 3290
rect 33876 3238 33906 3290
rect 33906 3238 33918 3290
rect 33918 3238 33932 3290
rect 33956 3238 33970 3290
rect 33970 3238 33982 3290
rect 33982 3238 34012 3290
rect 34036 3238 34046 3290
rect 34046 3238 34092 3290
rect 33796 3236 33852 3238
rect 33876 3236 33932 3238
rect 33956 3236 34012 3238
rect 34036 3236 34092 3238
rect 33796 2202 33852 2204
rect 33876 2202 33932 2204
rect 33956 2202 34012 2204
rect 34036 2202 34092 2204
rect 33796 2150 33842 2202
rect 33842 2150 33852 2202
rect 33876 2150 33906 2202
rect 33906 2150 33918 2202
rect 33918 2150 33932 2202
rect 33956 2150 33970 2202
rect 33970 2150 33982 2202
rect 33982 2150 34012 2202
rect 34036 2150 34046 2202
rect 34046 2150 34092 2202
rect 33796 2148 33852 2150
rect 33876 2148 33932 2150
rect 33956 2148 34012 2150
rect 34036 2148 34092 2150
rect 34426 1944 34482 2000
rect 35622 2624 35678 2680
rect 35990 2352 36046 2408
rect 37646 4120 37702 4176
rect 37738 3032 37794 3088
rect 39270 4922 39326 4924
rect 39350 4922 39406 4924
rect 39430 4922 39486 4924
rect 39510 4922 39566 4924
rect 39270 4870 39316 4922
rect 39316 4870 39326 4922
rect 39350 4870 39380 4922
rect 39380 4870 39392 4922
rect 39392 4870 39406 4922
rect 39430 4870 39444 4922
rect 39444 4870 39456 4922
rect 39456 4870 39486 4922
rect 39510 4870 39520 4922
rect 39520 4870 39566 4922
rect 39270 4868 39326 4870
rect 39350 4868 39406 4870
rect 39430 4868 39486 4870
rect 39510 4868 39566 4870
rect 40130 5344 40186 5400
rect 44743 5466 44799 5468
rect 44823 5466 44879 5468
rect 44903 5466 44959 5468
rect 44983 5466 45039 5468
rect 44743 5414 44789 5466
rect 44789 5414 44799 5466
rect 44823 5414 44853 5466
rect 44853 5414 44865 5466
rect 44865 5414 44879 5466
rect 44903 5414 44917 5466
rect 44917 5414 44929 5466
rect 44929 5414 44959 5466
rect 44983 5414 44993 5466
rect 44993 5414 45039 5466
rect 44743 5412 44799 5414
rect 44823 5412 44879 5414
rect 44903 5412 44959 5414
rect 44983 5412 45039 5414
rect 39302 3984 39358 4040
rect 39270 3834 39326 3836
rect 39350 3834 39406 3836
rect 39430 3834 39486 3836
rect 39510 3834 39566 3836
rect 39270 3782 39316 3834
rect 39316 3782 39326 3834
rect 39350 3782 39380 3834
rect 39380 3782 39392 3834
rect 39392 3782 39406 3834
rect 39430 3782 39444 3834
rect 39444 3782 39456 3834
rect 39456 3782 39486 3834
rect 39510 3782 39520 3834
rect 39520 3782 39566 3834
rect 39270 3780 39326 3782
rect 39350 3780 39406 3782
rect 39430 3780 39486 3782
rect 39510 3780 39566 3782
rect 38658 3440 38714 3496
rect 38014 2896 38070 2952
rect 39270 2746 39326 2748
rect 39350 2746 39406 2748
rect 39430 2746 39486 2748
rect 39510 2746 39566 2748
rect 39270 2694 39316 2746
rect 39316 2694 39326 2746
rect 39350 2694 39380 2746
rect 39380 2694 39392 2746
rect 39392 2694 39406 2746
rect 39430 2694 39444 2746
rect 39444 2694 39456 2746
rect 39456 2694 39486 2746
rect 39510 2694 39520 2746
rect 39520 2694 39566 2746
rect 39270 2692 39326 2694
rect 39350 2692 39406 2694
rect 39430 2692 39486 2694
rect 39510 2692 39566 2694
rect 41510 5072 41566 5128
rect 40498 4256 40554 4312
rect 39946 3576 40002 3632
rect 44743 4378 44799 4380
rect 44823 4378 44879 4380
rect 44903 4378 44959 4380
rect 44983 4378 45039 4380
rect 44743 4326 44789 4378
rect 44789 4326 44799 4378
rect 44823 4326 44853 4378
rect 44853 4326 44865 4378
rect 44865 4326 44879 4378
rect 44903 4326 44917 4378
rect 44917 4326 44929 4378
rect 44929 4326 44959 4378
rect 44983 4326 44993 4378
rect 44993 4326 45039 4378
rect 44743 4324 44799 4326
rect 44823 4324 44879 4326
rect 44903 4324 44959 4326
rect 44983 4324 45039 4326
rect 44743 3290 44799 3292
rect 44823 3290 44879 3292
rect 44903 3290 44959 3292
rect 44983 3290 45039 3292
rect 44743 3238 44789 3290
rect 44789 3238 44799 3290
rect 44823 3238 44853 3290
rect 44853 3238 44865 3290
rect 44865 3238 44879 3290
rect 44903 3238 44917 3290
rect 44917 3238 44929 3290
rect 44929 3238 44959 3290
rect 44983 3238 44993 3290
rect 44993 3238 45039 3290
rect 44743 3236 44799 3238
rect 44823 3236 44879 3238
rect 44903 3236 44959 3238
rect 44983 3236 45039 3238
rect 36266 1672 36322 1728
rect 44743 2202 44799 2204
rect 44823 2202 44879 2204
rect 44903 2202 44959 2204
rect 44983 2202 45039 2204
rect 44743 2150 44789 2202
rect 44789 2150 44799 2202
rect 44823 2150 44853 2202
rect 44853 2150 44865 2202
rect 44865 2150 44879 2202
rect 44903 2150 44917 2202
rect 44917 2150 44929 2202
rect 44929 2150 44959 2202
rect 44983 2150 44993 2202
rect 44993 2150 45039 2202
rect 44743 2148 44799 2150
rect 44823 2148 44879 2150
rect 44903 2148 44959 2150
rect 44983 2148 45039 2150
<< metal3 >>
rect 6177 5810 6243 5813
rect 19333 5810 19399 5813
rect 6177 5808 19399 5810
rect 6177 5752 6182 5808
rect 6238 5752 19338 5808
rect 19394 5752 19399 5808
rect 6177 5750 19399 5752
rect 6177 5747 6243 5750
rect 19333 5747 19399 5750
rect 6729 5674 6795 5677
rect 19609 5674 19675 5677
rect 6729 5672 19675 5674
rect 6729 5616 6734 5672
rect 6790 5616 19614 5672
rect 19670 5616 19675 5672
rect 6729 5614 19675 5616
rect 6729 5611 6795 5614
rect 19609 5611 19675 5614
rect 11892 5472 12208 5473
rect 11892 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12208 5472
rect 11892 5407 12208 5408
rect 22839 5472 23155 5473
rect 22839 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23155 5472
rect 22839 5407 23155 5408
rect 33786 5472 34102 5473
rect 33786 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34102 5472
rect 33786 5407 34102 5408
rect 44733 5472 45049 5473
rect 44733 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45049 5472
rect 44733 5407 45049 5408
rect 19793 5402 19859 5405
rect 20437 5402 20503 5405
rect 19793 5400 20503 5402
rect 19793 5344 19798 5400
rect 19854 5344 20442 5400
rect 20498 5344 20503 5400
rect 19793 5342 20503 5344
rect 19793 5339 19859 5342
rect 20437 5339 20503 5342
rect 34513 5402 34579 5405
rect 40125 5402 40191 5405
rect 34513 5400 40191 5402
rect 34513 5344 34518 5400
rect 34574 5344 40130 5400
rect 40186 5344 40191 5400
rect 34513 5342 40191 5344
rect 34513 5339 34579 5342
rect 40125 5339 40191 5342
rect 7005 5266 7071 5269
rect 24393 5266 24459 5269
rect 7005 5264 24459 5266
rect 7005 5208 7010 5264
rect 7066 5208 24398 5264
rect 24454 5208 24459 5264
rect 7005 5206 24459 5208
rect 7005 5203 7071 5206
rect 24393 5203 24459 5206
rect 15101 5130 15167 5133
rect 23381 5130 23447 5133
rect 15101 5128 23447 5130
rect 15101 5072 15106 5128
rect 15162 5072 23386 5128
rect 23442 5072 23447 5128
rect 15101 5070 23447 5072
rect 15101 5067 15167 5070
rect 23381 5067 23447 5070
rect 33133 5130 33199 5133
rect 41505 5130 41571 5133
rect 33133 5128 41571 5130
rect 33133 5072 33138 5128
rect 33194 5072 41510 5128
rect 41566 5072 41571 5128
rect 33133 5070 41571 5072
rect 33133 5067 33199 5070
rect 41505 5067 41571 5070
rect 11881 4994 11947 4997
rect 16021 4994 16087 4997
rect 11881 4992 16087 4994
rect 11881 4936 11886 4992
rect 11942 4936 16026 4992
rect 16082 4936 16087 4992
rect 11881 4934 16087 4936
rect 11881 4931 11947 4934
rect 16021 4931 16087 4934
rect 19517 4994 19583 4997
rect 27797 4994 27863 4997
rect 19517 4992 27863 4994
rect 19517 4936 19522 4992
rect 19578 4936 27802 4992
rect 27858 4936 27863 4992
rect 19517 4934 27863 4936
rect 19517 4931 19583 4934
rect 27797 4931 27863 4934
rect 6419 4928 6735 4929
rect 6419 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6735 4928
rect 6419 4863 6735 4864
rect 17366 4928 17682 4929
rect 17366 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17682 4928
rect 17366 4863 17682 4864
rect 28313 4928 28629 4929
rect 28313 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28629 4928
rect 28313 4863 28629 4864
rect 39260 4928 39576 4929
rect 39260 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39576 4928
rect 39260 4863 39576 4864
rect 11697 4858 11763 4861
rect 16573 4858 16639 4861
rect 11697 4856 16639 4858
rect 11697 4800 11702 4856
rect 11758 4800 16578 4856
rect 16634 4800 16639 4856
rect 11697 4798 16639 4800
rect 11697 4795 11763 4798
rect 16573 4795 16639 4798
rect 19885 4858 19951 4861
rect 21449 4858 21515 4861
rect 19885 4856 21515 4858
rect 19885 4800 19890 4856
rect 19946 4800 21454 4856
rect 21510 4800 21515 4856
rect 19885 4798 21515 4800
rect 19885 4795 19951 4798
rect 21449 4795 21515 4798
rect 22001 4858 22067 4861
rect 22185 4858 22251 4861
rect 22001 4856 22251 4858
rect 22001 4800 22006 4856
rect 22062 4800 22190 4856
rect 22246 4800 22251 4856
rect 22001 4798 22251 4800
rect 22001 4795 22067 4798
rect 22185 4795 22251 4798
rect 23013 4858 23079 4861
rect 27613 4858 27679 4861
rect 23013 4856 27679 4858
rect 23013 4800 23018 4856
rect 23074 4800 27618 4856
rect 27674 4800 27679 4856
rect 23013 4798 27679 4800
rect 23013 4795 23079 4798
rect 27613 4795 27679 4798
rect 11237 4722 11303 4725
rect 12341 4722 12407 4725
rect 11237 4720 12407 4722
rect 11237 4664 11242 4720
rect 11298 4664 12346 4720
rect 12402 4664 12407 4720
rect 11237 4662 12407 4664
rect 11237 4659 11303 4662
rect 12341 4659 12407 4662
rect 15101 4722 15167 4725
rect 28441 4722 28507 4725
rect 15101 4720 28507 4722
rect 15101 4664 15106 4720
rect 15162 4664 28446 4720
rect 28502 4664 28507 4720
rect 15101 4662 28507 4664
rect 15101 4659 15167 4662
rect 28441 4659 28507 4662
rect 13261 4586 13327 4589
rect 29729 4586 29795 4589
rect 10918 4526 12450 4586
rect 9397 4450 9463 4453
rect 10918 4450 10978 4526
rect 9397 4448 10978 4450
rect 9397 4392 9402 4448
rect 9458 4392 10978 4448
rect 9397 4390 10978 4392
rect 12390 4450 12450 4526
rect 13261 4584 29795 4586
rect 13261 4528 13266 4584
rect 13322 4528 29734 4584
rect 29790 4528 29795 4584
rect 13261 4526 29795 4528
rect 13261 4523 13327 4526
rect 29729 4523 29795 4526
rect 22277 4450 22343 4453
rect 12390 4448 22343 4450
rect 12390 4392 22282 4448
rect 22338 4392 22343 4448
rect 12390 4390 22343 4392
rect 9397 4387 9463 4390
rect 22277 4387 22343 4390
rect 11892 4384 12208 4385
rect 11892 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12208 4384
rect 11892 4319 12208 4320
rect 22839 4384 23155 4385
rect 22839 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23155 4384
rect 22839 4319 23155 4320
rect 33786 4384 34102 4385
rect 33786 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34102 4384
rect 33786 4319 34102 4320
rect 44733 4384 45049 4385
rect 44733 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45049 4384
rect 44733 4319 45049 4320
rect 12433 4314 12499 4317
rect 22645 4314 22711 4317
rect 12433 4312 22711 4314
rect 12433 4256 12438 4312
rect 12494 4256 22650 4312
rect 22706 4256 22711 4312
rect 12433 4254 22711 4256
rect 12433 4251 12499 4254
rect 22645 4251 22711 4254
rect 37222 4252 37228 4316
rect 37292 4314 37298 4316
rect 40493 4314 40559 4317
rect 37292 4312 40559 4314
rect 37292 4256 40498 4312
rect 40554 4256 40559 4312
rect 37292 4254 40559 4256
rect 37292 4252 37298 4254
rect 40493 4251 40559 4254
rect 11237 4178 11303 4181
rect 22737 4178 22803 4181
rect 11237 4176 22803 4178
rect 11237 4120 11242 4176
rect 11298 4120 22742 4176
rect 22798 4120 22803 4176
rect 11237 4118 22803 4120
rect 11237 4115 11303 4118
rect 22737 4115 22803 4118
rect 24209 4178 24275 4181
rect 37641 4178 37707 4181
rect 24209 4176 37707 4178
rect 24209 4120 24214 4176
rect 24270 4120 37646 4176
rect 37702 4120 37707 4176
rect 24209 4118 37707 4120
rect 24209 4115 24275 4118
rect 37641 4115 37707 4118
rect 18229 4042 18295 4045
rect 39297 4042 39363 4045
rect 17174 3982 18154 4042
rect 14181 3906 14247 3909
rect 17174 3906 17234 3982
rect 14181 3904 17234 3906
rect 14181 3848 14186 3904
rect 14242 3848 17234 3904
rect 14181 3846 17234 3848
rect 18094 3906 18154 3982
rect 18229 4040 39363 4042
rect 18229 3984 18234 4040
rect 18290 3984 39302 4040
rect 39358 3984 39363 4040
rect 18229 3982 39363 3984
rect 18229 3979 18295 3982
rect 39297 3979 39363 3982
rect 28165 3906 28231 3909
rect 18094 3904 28231 3906
rect 18094 3848 28170 3904
rect 28226 3848 28231 3904
rect 18094 3846 28231 3848
rect 14181 3843 14247 3846
rect 28165 3843 28231 3846
rect 28717 3906 28783 3909
rect 37222 3906 37228 3908
rect 28717 3904 37228 3906
rect 28717 3848 28722 3904
rect 28778 3848 37228 3904
rect 28717 3846 37228 3848
rect 28717 3843 28783 3846
rect 37222 3844 37228 3846
rect 37292 3844 37298 3908
rect 6419 3840 6735 3841
rect 6419 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6735 3840
rect 6419 3775 6735 3776
rect 17366 3840 17682 3841
rect 17366 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17682 3840
rect 17366 3775 17682 3776
rect 28313 3840 28629 3841
rect 28313 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28629 3840
rect 28313 3775 28629 3776
rect 39260 3840 39576 3841
rect 39260 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39576 3840
rect 39260 3775 39576 3776
rect 11973 3634 12039 3637
rect 13445 3634 13511 3637
rect 39941 3634 40007 3637
rect 11973 3632 12450 3634
rect 11973 3576 11978 3632
rect 12034 3576 12450 3632
rect 11973 3574 12450 3576
rect 11973 3571 12039 3574
rect 12390 3362 12450 3574
rect 13445 3632 40007 3634
rect 13445 3576 13450 3632
rect 13506 3576 39946 3632
rect 40002 3576 40007 3632
rect 13445 3574 40007 3576
rect 13445 3571 13511 3574
rect 39941 3571 40007 3574
rect 14549 3498 14615 3501
rect 38653 3498 38719 3501
rect 14549 3496 38719 3498
rect 14549 3440 14554 3496
rect 14610 3440 38658 3496
rect 38714 3440 38719 3496
rect 14549 3438 38719 3440
rect 14549 3435 14615 3438
rect 38653 3435 38719 3438
rect 18229 3362 18295 3365
rect 12390 3360 18295 3362
rect 12390 3304 18234 3360
rect 18290 3304 18295 3360
rect 12390 3302 18295 3304
rect 18229 3299 18295 3302
rect 11892 3296 12208 3297
rect 11892 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12208 3296
rect 11892 3231 12208 3232
rect 22839 3296 23155 3297
rect 22839 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23155 3296
rect 22839 3231 23155 3232
rect 33786 3296 34102 3297
rect 33786 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34102 3296
rect 33786 3231 34102 3232
rect 44733 3296 45049 3297
rect 44733 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45049 3296
rect 44733 3231 45049 3232
rect 15193 3226 15259 3229
rect 22645 3226 22711 3229
rect 15193 3224 22711 3226
rect 15193 3168 15198 3224
rect 15254 3168 22650 3224
rect 22706 3168 22711 3224
rect 15193 3166 22711 3168
rect 15193 3163 15259 3166
rect 22645 3163 22711 3166
rect 11237 3090 11303 3093
rect 37733 3090 37799 3093
rect 11237 3088 37799 3090
rect 11237 3032 11242 3088
rect 11298 3032 37738 3088
rect 37794 3032 37799 3088
rect 11237 3030 37799 3032
rect 11237 3027 11303 3030
rect 37733 3027 37799 3030
rect 10501 2954 10567 2957
rect 38009 2954 38075 2957
rect 10501 2952 38075 2954
rect 10501 2896 10506 2952
rect 10562 2896 38014 2952
rect 38070 2896 38075 2952
rect 10501 2894 38075 2896
rect 10501 2891 10567 2894
rect 38009 2891 38075 2894
rect 22645 2818 22711 2821
rect 26049 2818 26115 2821
rect 22645 2816 26115 2818
rect 22645 2760 22650 2816
rect 22706 2760 26054 2816
rect 26110 2760 26115 2816
rect 22645 2758 26115 2760
rect 22645 2755 22711 2758
rect 26049 2755 26115 2758
rect 6419 2752 6735 2753
rect 6419 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6735 2752
rect 6419 2687 6735 2688
rect 17366 2752 17682 2753
rect 17366 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17682 2752
rect 17366 2687 17682 2688
rect 28313 2752 28629 2753
rect 28313 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28629 2752
rect 28313 2687 28629 2688
rect 39260 2752 39576 2753
rect 39260 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39576 2752
rect 39260 2687 39576 2688
rect 35617 2682 35683 2685
rect 30974 2680 35683 2682
rect 30974 2624 35622 2680
rect 35678 2624 35683 2680
rect 30974 2622 35683 2624
rect 4705 2546 4771 2549
rect 30974 2546 31034 2622
rect 35617 2619 35683 2622
rect 4705 2544 31034 2546
rect 4705 2488 4710 2544
rect 4766 2488 31034 2544
rect 4705 2486 31034 2488
rect 4705 2483 4771 2486
rect 5901 2410 5967 2413
rect 35985 2410 36051 2413
rect 5901 2408 36051 2410
rect 5901 2352 5906 2408
rect 5962 2352 35990 2408
rect 36046 2352 36051 2408
rect 5901 2350 36051 2352
rect 5901 2347 5967 2350
rect 35985 2347 36051 2350
rect 11892 2208 12208 2209
rect 11892 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12208 2208
rect 11892 2143 12208 2144
rect 22839 2208 23155 2209
rect 22839 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23155 2208
rect 22839 2143 23155 2144
rect 33786 2208 34102 2209
rect 33786 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34102 2208
rect 33786 2143 34102 2144
rect 44733 2208 45049 2209
rect 44733 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45049 2208
rect 44733 2143 45049 2144
rect 8477 2002 8543 2005
rect 34421 2002 34487 2005
rect 8477 2000 34487 2002
rect 8477 1944 8482 2000
rect 8538 1944 34426 2000
rect 34482 1944 34487 2000
rect 8477 1942 34487 1944
rect 8477 1939 8543 1942
rect 34421 1939 34487 1942
rect 9213 1866 9279 1869
rect 27981 1866 28047 1869
rect 9213 1864 28047 1866
rect 9213 1808 9218 1864
rect 9274 1808 27986 1864
rect 28042 1808 28047 1864
rect 9213 1806 28047 1808
rect 9213 1803 9279 1806
rect 27981 1803 28047 1806
rect 7097 1730 7163 1733
rect 36261 1730 36327 1733
rect 7097 1728 36327 1730
rect 7097 1672 7102 1728
rect 7158 1672 36266 1728
rect 36322 1672 36327 1728
rect 7097 1670 36327 1672
rect 7097 1667 7163 1670
rect 36261 1667 36327 1670
<< via3 >>
rect 11898 5468 11962 5472
rect 11898 5412 11902 5468
rect 11902 5412 11958 5468
rect 11958 5412 11962 5468
rect 11898 5408 11962 5412
rect 11978 5468 12042 5472
rect 11978 5412 11982 5468
rect 11982 5412 12038 5468
rect 12038 5412 12042 5468
rect 11978 5408 12042 5412
rect 12058 5468 12122 5472
rect 12058 5412 12062 5468
rect 12062 5412 12118 5468
rect 12118 5412 12122 5468
rect 12058 5408 12122 5412
rect 12138 5468 12202 5472
rect 12138 5412 12142 5468
rect 12142 5412 12198 5468
rect 12198 5412 12202 5468
rect 12138 5408 12202 5412
rect 22845 5468 22909 5472
rect 22845 5412 22849 5468
rect 22849 5412 22905 5468
rect 22905 5412 22909 5468
rect 22845 5408 22909 5412
rect 22925 5468 22989 5472
rect 22925 5412 22929 5468
rect 22929 5412 22985 5468
rect 22985 5412 22989 5468
rect 22925 5408 22989 5412
rect 23005 5468 23069 5472
rect 23005 5412 23009 5468
rect 23009 5412 23065 5468
rect 23065 5412 23069 5468
rect 23005 5408 23069 5412
rect 23085 5468 23149 5472
rect 23085 5412 23089 5468
rect 23089 5412 23145 5468
rect 23145 5412 23149 5468
rect 23085 5408 23149 5412
rect 33792 5468 33856 5472
rect 33792 5412 33796 5468
rect 33796 5412 33852 5468
rect 33852 5412 33856 5468
rect 33792 5408 33856 5412
rect 33872 5468 33936 5472
rect 33872 5412 33876 5468
rect 33876 5412 33932 5468
rect 33932 5412 33936 5468
rect 33872 5408 33936 5412
rect 33952 5468 34016 5472
rect 33952 5412 33956 5468
rect 33956 5412 34012 5468
rect 34012 5412 34016 5468
rect 33952 5408 34016 5412
rect 34032 5468 34096 5472
rect 34032 5412 34036 5468
rect 34036 5412 34092 5468
rect 34092 5412 34096 5468
rect 34032 5408 34096 5412
rect 44739 5468 44803 5472
rect 44739 5412 44743 5468
rect 44743 5412 44799 5468
rect 44799 5412 44803 5468
rect 44739 5408 44803 5412
rect 44819 5468 44883 5472
rect 44819 5412 44823 5468
rect 44823 5412 44879 5468
rect 44879 5412 44883 5468
rect 44819 5408 44883 5412
rect 44899 5468 44963 5472
rect 44899 5412 44903 5468
rect 44903 5412 44959 5468
rect 44959 5412 44963 5468
rect 44899 5408 44963 5412
rect 44979 5468 45043 5472
rect 44979 5412 44983 5468
rect 44983 5412 45039 5468
rect 45039 5412 45043 5468
rect 44979 5408 45043 5412
rect 6425 4924 6489 4928
rect 6425 4868 6429 4924
rect 6429 4868 6485 4924
rect 6485 4868 6489 4924
rect 6425 4864 6489 4868
rect 6505 4924 6569 4928
rect 6505 4868 6509 4924
rect 6509 4868 6565 4924
rect 6565 4868 6569 4924
rect 6505 4864 6569 4868
rect 6585 4924 6649 4928
rect 6585 4868 6589 4924
rect 6589 4868 6645 4924
rect 6645 4868 6649 4924
rect 6585 4864 6649 4868
rect 6665 4924 6729 4928
rect 6665 4868 6669 4924
rect 6669 4868 6725 4924
rect 6725 4868 6729 4924
rect 6665 4864 6729 4868
rect 17372 4924 17436 4928
rect 17372 4868 17376 4924
rect 17376 4868 17432 4924
rect 17432 4868 17436 4924
rect 17372 4864 17436 4868
rect 17452 4924 17516 4928
rect 17452 4868 17456 4924
rect 17456 4868 17512 4924
rect 17512 4868 17516 4924
rect 17452 4864 17516 4868
rect 17532 4924 17596 4928
rect 17532 4868 17536 4924
rect 17536 4868 17592 4924
rect 17592 4868 17596 4924
rect 17532 4864 17596 4868
rect 17612 4924 17676 4928
rect 17612 4868 17616 4924
rect 17616 4868 17672 4924
rect 17672 4868 17676 4924
rect 17612 4864 17676 4868
rect 28319 4924 28383 4928
rect 28319 4868 28323 4924
rect 28323 4868 28379 4924
rect 28379 4868 28383 4924
rect 28319 4864 28383 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 39266 4924 39330 4928
rect 39266 4868 39270 4924
rect 39270 4868 39326 4924
rect 39326 4868 39330 4924
rect 39266 4864 39330 4868
rect 39346 4924 39410 4928
rect 39346 4868 39350 4924
rect 39350 4868 39406 4924
rect 39406 4868 39410 4924
rect 39346 4864 39410 4868
rect 39426 4924 39490 4928
rect 39426 4868 39430 4924
rect 39430 4868 39486 4924
rect 39486 4868 39490 4924
rect 39426 4864 39490 4868
rect 39506 4924 39570 4928
rect 39506 4868 39510 4924
rect 39510 4868 39566 4924
rect 39566 4868 39570 4924
rect 39506 4864 39570 4868
rect 11898 4380 11962 4384
rect 11898 4324 11902 4380
rect 11902 4324 11958 4380
rect 11958 4324 11962 4380
rect 11898 4320 11962 4324
rect 11978 4380 12042 4384
rect 11978 4324 11982 4380
rect 11982 4324 12038 4380
rect 12038 4324 12042 4380
rect 11978 4320 12042 4324
rect 12058 4380 12122 4384
rect 12058 4324 12062 4380
rect 12062 4324 12118 4380
rect 12118 4324 12122 4380
rect 12058 4320 12122 4324
rect 12138 4380 12202 4384
rect 12138 4324 12142 4380
rect 12142 4324 12198 4380
rect 12198 4324 12202 4380
rect 12138 4320 12202 4324
rect 22845 4380 22909 4384
rect 22845 4324 22849 4380
rect 22849 4324 22905 4380
rect 22905 4324 22909 4380
rect 22845 4320 22909 4324
rect 22925 4380 22989 4384
rect 22925 4324 22929 4380
rect 22929 4324 22985 4380
rect 22985 4324 22989 4380
rect 22925 4320 22989 4324
rect 23005 4380 23069 4384
rect 23005 4324 23009 4380
rect 23009 4324 23065 4380
rect 23065 4324 23069 4380
rect 23005 4320 23069 4324
rect 23085 4380 23149 4384
rect 23085 4324 23089 4380
rect 23089 4324 23145 4380
rect 23145 4324 23149 4380
rect 23085 4320 23149 4324
rect 33792 4380 33856 4384
rect 33792 4324 33796 4380
rect 33796 4324 33852 4380
rect 33852 4324 33856 4380
rect 33792 4320 33856 4324
rect 33872 4380 33936 4384
rect 33872 4324 33876 4380
rect 33876 4324 33932 4380
rect 33932 4324 33936 4380
rect 33872 4320 33936 4324
rect 33952 4380 34016 4384
rect 33952 4324 33956 4380
rect 33956 4324 34012 4380
rect 34012 4324 34016 4380
rect 33952 4320 34016 4324
rect 34032 4380 34096 4384
rect 34032 4324 34036 4380
rect 34036 4324 34092 4380
rect 34092 4324 34096 4380
rect 34032 4320 34096 4324
rect 44739 4380 44803 4384
rect 44739 4324 44743 4380
rect 44743 4324 44799 4380
rect 44799 4324 44803 4380
rect 44739 4320 44803 4324
rect 44819 4380 44883 4384
rect 44819 4324 44823 4380
rect 44823 4324 44879 4380
rect 44879 4324 44883 4380
rect 44819 4320 44883 4324
rect 44899 4380 44963 4384
rect 44899 4324 44903 4380
rect 44903 4324 44959 4380
rect 44959 4324 44963 4380
rect 44899 4320 44963 4324
rect 44979 4380 45043 4384
rect 44979 4324 44983 4380
rect 44983 4324 45039 4380
rect 45039 4324 45043 4380
rect 44979 4320 45043 4324
rect 37228 4252 37292 4316
rect 37228 3844 37292 3908
rect 6425 3836 6489 3840
rect 6425 3780 6429 3836
rect 6429 3780 6485 3836
rect 6485 3780 6489 3836
rect 6425 3776 6489 3780
rect 6505 3836 6569 3840
rect 6505 3780 6509 3836
rect 6509 3780 6565 3836
rect 6565 3780 6569 3836
rect 6505 3776 6569 3780
rect 6585 3836 6649 3840
rect 6585 3780 6589 3836
rect 6589 3780 6645 3836
rect 6645 3780 6649 3836
rect 6585 3776 6649 3780
rect 6665 3836 6729 3840
rect 6665 3780 6669 3836
rect 6669 3780 6725 3836
rect 6725 3780 6729 3836
rect 6665 3776 6729 3780
rect 17372 3836 17436 3840
rect 17372 3780 17376 3836
rect 17376 3780 17432 3836
rect 17432 3780 17436 3836
rect 17372 3776 17436 3780
rect 17452 3836 17516 3840
rect 17452 3780 17456 3836
rect 17456 3780 17512 3836
rect 17512 3780 17516 3836
rect 17452 3776 17516 3780
rect 17532 3836 17596 3840
rect 17532 3780 17536 3836
rect 17536 3780 17592 3836
rect 17592 3780 17596 3836
rect 17532 3776 17596 3780
rect 17612 3836 17676 3840
rect 17612 3780 17616 3836
rect 17616 3780 17672 3836
rect 17672 3780 17676 3836
rect 17612 3776 17676 3780
rect 28319 3836 28383 3840
rect 28319 3780 28323 3836
rect 28323 3780 28379 3836
rect 28379 3780 28383 3836
rect 28319 3776 28383 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 39266 3836 39330 3840
rect 39266 3780 39270 3836
rect 39270 3780 39326 3836
rect 39326 3780 39330 3836
rect 39266 3776 39330 3780
rect 39346 3836 39410 3840
rect 39346 3780 39350 3836
rect 39350 3780 39406 3836
rect 39406 3780 39410 3836
rect 39346 3776 39410 3780
rect 39426 3836 39490 3840
rect 39426 3780 39430 3836
rect 39430 3780 39486 3836
rect 39486 3780 39490 3836
rect 39426 3776 39490 3780
rect 39506 3836 39570 3840
rect 39506 3780 39510 3836
rect 39510 3780 39566 3836
rect 39566 3780 39570 3836
rect 39506 3776 39570 3780
rect 11898 3292 11962 3296
rect 11898 3236 11902 3292
rect 11902 3236 11958 3292
rect 11958 3236 11962 3292
rect 11898 3232 11962 3236
rect 11978 3292 12042 3296
rect 11978 3236 11982 3292
rect 11982 3236 12038 3292
rect 12038 3236 12042 3292
rect 11978 3232 12042 3236
rect 12058 3292 12122 3296
rect 12058 3236 12062 3292
rect 12062 3236 12118 3292
rect 12118 3236 12122 3292
rect 12058 3232 12122 3236
rect 12138 3292 12202 3296
rect 12138 3236 12142 3292
rect 12142 3236 12198 3292
rect 12198 3236 12202 3292
rect 12138 3232 12202 3236
rect 22845 3292 22909 3296
rect 22845 3236 22849 3292
rect 22849 3236 22905 3292
rect 22905 3236 22909 3292
rect 22845 3232 22909 3236
rect 22925 3292 22989 3296
rect 22925 3236 22929 3292
rect 22929 3236 22985 3292
rect 22985 3236 22989 3292
rect 22925 3232 22989 3236
rect 23005 3292 23069 3296
rect 23005 3236 23009 3292
rect 23009 3236 23065 3292
rect 23065 3236 23069 3292
rect 23005 3232 23069 3236
rect 23085 3292 23149 3296
rect 23085 3236 23089 3292
rect 23089 3236 23145 3292
rect 23145 3236 23149 3292
rect 23085 3232 23149 3236
rect 33792 3292 33856 3296
rect 33792 3236 33796 3292
rect 33796 3236 33852 3292
rect 33852 3236 33856 3292
rect 33792 3232 33856 3236
rect 33872 3292 33936 3296
rect 33872 3236 33876 3292
rect 33876 3236 33932 3292
rect 33932 3236 33936 3292
rect 33872 3232 33936 3236
rect 33952 3292 34016 3296
rect 33952 3236 33956 3292
rect 33956 3236 34012 3292
rect 34012 3236 34016 3292
rect 33952 3232 34016 3236
rect 34032 3292 34096 3296
rect 34032 3236 34036 3292
rect 34036 3236 34092 3292
rect 34092 3236 34096 3292
rect 34032 3232 34096 3236
rect 44739 3292 44803 3296
rect 44739 3236 44743 3292
rect 44743 3236 44799 3292
rect 44799 3236 44803 3292
rect 44739 3232 44803 3236
rect 44819 3292 44883 3296
rect 44819 3236 44823 3292
rect 44823 3236 44879 3292
rect 44879 3236 44883 3292
rect 44819 3232 44883 3236
rect 44899 3292 44963 3296
rect 44899 3236 44903 3292
rect 44903 3236 44959 3292
rect 44959 3236 44963 3292
rect 44899 3232 44963 3236
rect 44979 3292 45043 3296
rect 44979 3236 44983 3292
rect 44983 3236 45039 3292
rect 45039 3236 45043 3292
rect 44979 3232 45043 3236
rect 6425 2748 6489 2752
rect 6425 2692 6429 2748
rect 6429 2692 6485 2748
rect 6485 2692 6489 2748
rect 6425 2688 6489 2692
rect 6505 2748 6569 2752
rect 6505 2692 6509 2748
rect 6509 2692 6565 2748
rect 6565 2692 6569 2748
rect 6505 2688 6569 2692
rect 6585 2748 6649 2752
rect 6585 2692 6589 2748
rect 6589 2692 6645 2748
rect 6645 2692 6649 2748
rect 6585 2688 6649 2692
rect 6665 2748 6729 2752
rect 6665 2692 6669 2748
rect 6669 2692 6725 2748
rect 6725 2692 6729 2748
rect 6665 2688 6729 2692
rect 17372 2748 17436 2752
rect 17372 2692 17376 2748
rect 17376 2692 17432 2748
rect 17432 2692 17436 2748
rect 17372 2688 17436 2692
rect 17452 2748 17516 2752
rect 17452 2692 17456 2748
rect 17456 2692 17512 2748
rect 17512 2692 17516 2748
rect 17452 2688 17516 2692
rect 17532 2748 17596 2752
rect 17532 2692 17536 2748
rect 17536 2692 17592 2748
rect 17592 2692 17596 2748
rect 17532 2688 17596 2692
rect 17612 2748 17676 2752
rect 17612 2692 17616 2748
rect 17616 2692 17672 2748
rect 17672 2692 17676 2748
rect 17612 2688 17676 2692
rect 28319 2748 28383 2752
rect 28319 2692 28323 2748
rect 28323 2692 28379 2748
rect 28379 2692 28383 2748
rect 28319 2688 28383 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 39266 2748 39330 2752
rect 39266 2692 39270 2748
rect 39270 2692 39326 2748
rect 39326 2692 39330 2748
rect 39266 2688 39330 2692
rect 39346 2748 39410 2752
rect 39346 2692 39350 2748
rect 39350 2692 39406 2748
rect 39406 2692 39410 2748
rect 39346 2688 39410 2692
rect 39426 2748 39490 2752
rect 39426 2692 39430 2748
rect 39430 2692 39486 2748
rect 39486 2692 39490 2748
rect 39426 2688 39490 2692
rect 39506 2748 39570 2752
rect 39506 2692 39510 2748
rect 39510 2692 39566 2748
rect 39566 2692 39570 2748
rect 39506 2688 39570 2692
rect 11898 2204 11962 2208
rect 11898 2148 11902 2204
rect 11902 2148 11958 2204
rect 11958 2148 11962 2204
rect 11898 2144 11962 2148
rect 11978 2204 12042 2208
rect 11978 2148 11982 2204
rect 11982 2148 12038 2204
rect 12038 2148 12042 2204
rect 11978 2144 12042 2148
rect 12058 2204 12122 2208
rect 12058 2148 12062 2204
rect 12062 2148 12118 2204
rect 12118 2148 12122 2204
rect 12058 2144 12122 2148
rect 12138 2204 12202 2208
rect 12138 2148 12142 2204
rect 12142 2148 12198 2204
rect 12198 2148 12202 2204
rect 12138 2144 12202 2148
rect 22845 2204 22909 2208
rect 22845 2148 22849 2204
rect 22849 2148 22905 2204
rect 22905 2148 22909 2204
rect 22845 2144 22909 2148
rect 22925 2204 22989 2208
rect 22925 2148 22929 2204
rect 22929 2148 22985 2204
rect 22985 2148 22989 2204
rect 22925 2144 22989 2148
rect 23005 2204 23069 2208
rect 23005 2148 23009 2204
rect 23009 2148 23065 2204
rect 23065 2148 23069 2204
rect 23005 2144 23069 2148
rect 23085 2204 23149 2208
rect 23085 2148 23089 2204
rect 23089 2148 23145 2204
rect 23145 2148 23149 2204
rect 23085 2144 23149 2148
rect 33792 2204 33856 2208
rect 33792 2148 33796 2204
rect 33796 2148 33852 2204
rect 33852 2148 33856 2204
rect 33792 2144 33856 2148
rect 33872 2204 33936 2208
rect 33872 2148 33876 2204
rect 33876 2148 33932 2204
rect 33932 2148 33936 2204
rect 33872 2144 33936 2148
rect 33952 2204 34016 2208
rect 33952 2148 33956 2204
rect 33956 2148 34012 2204
rect 34012 2148 34016 2204
rect 33952 2144 34016 2148
rect 34032 2204 34096 2208
rect 34032 2148 34036 2204
rect 34036 2148 34092 2204
rect 34092 2148 34096 2204
rect 34032 2144 34096 2148
rect 44739 2204 44803 2208
rect 44739 2148 44743 2204
rect 44743 2148 44799 2204
rect 44799 2148 44803 2204
rect 44739 2144 44803 2148
rect 44819 2204 44883 2208
rect 44819 2148 44823 2204
rect 44823 2148 44879 2204
rect 44879 2148 44883 2204
rect 44819 2144 44883 2148
rect 44899 2204 44963 2208
rect 44899 2148 44903 2204
rect 44903 2148 44959 2204
rect 44959 2148 44963 2204
rect 44899 2144 44963 2148
rect 44979 2204 45043 2208
rect 44979 2148 44983 2204
rect 44983 2148 45039 2204
rect 45039 2148 45043 2204
rect 44979 2144 45043 2148
<< metal4 >>
rect 6417 4928 6737 5488
rect 6417 4864 6425 4928
rect 6489 4864 6505 4928
rect 6569 4864 6585 4928
rect 6649 4864 6665 4928
rect 6729 4864 6737 4928
rect 6417 3840 6737 4864
rect 6417 3776 6425 3840
rect 6489 3776 6505 3840
rect 6569 3776 6585 3840
rect 6649 3776 6665 3840
rect 6729 3776 6737 3840
rect 6417 2752 6737 3776
rect 6417 2688 6425 2752
rect 6489 2688 6505 2752
rect 6569 2688 6585 2752
rect 6649 2688 6665 2752
rect 6729 2688 6737 2752
rect 6417 2128 6737 2688
rect 11890 5472 12210 5488
rect 11890 5408 11898 5472
rect 11962 5408 11978 5472
rect 12042 5408 12058 5472
rect 12122 5408 12138 5472
rect 12202 5408 12210 5472
rect 11890 4384 12210 5408
rect 11890 4320 11898 4384
rect 11962 4320 11978 4384
rect 12042 4320 12058 4384
rect 12122 4320 12138 4384
rect 12202 4320 12210 4384
rect 11890 3296 12210 4320
rect 11890 3232 11898 3296
rect 11962 3232 11978 3296
rect 12042 3232 12058 3296
rect 12122 3232 12138 3296
rect 12202 3232 12210 3296
rect 11890 2208 12210 3232
rect 11890 2144 11898 2208
rect 11962 2144 11978 2208
rect 12042 2144 12058 2208
rect 12122 2144 12138 2208
rect 12202 2144 12210 2208
rect 11890 2128 12210 2144
rect 17364 4928 17684 5488
rect 17364 4864 17372 4928
rect 17436 4864 17452 4928
rect 17516 4864 17532 4928
rect 17596 4864 17612 4928
rect 17676 4864 17684 4928
rect 17364 3840 17684 4864
rect 17364 3776 17372 3840
rect 17436 3776 17452 3840
rect 17516 3776 17532 3840
rect 17596 3776 17612 3840
rect 17676 3776 17684 3840
rect 17364 2752 17684 3776
rect 17364 2688 17372 2752
rect 17436 2688 17452 2752
rect 17516 2688 17532 2752
rect 17596 2688 17612 2752
rect 17676 2688 17684 2752
rect 17364 2128 17684 2688
rect 22837 5472 23157 5488
rect 22837 5408 22845 5472
rect 22909 5408 22925 5472
rect 22989 5408 23005 5472
rect 23069 5408 23085 5472
rect 23149 5408 23157 5472
rect 22837 4384 23157 5408
rect 22837 4320 22845 4384
rect 22909 4320 22925 4384
rect 22989 4320 23005 4384
rect 23069 4320 23085 4384
rect 23149 4320 23157 4384
rect 22837 3296 23157 4320
rect 22837 3232 22845 3296
rect 22909 3232 22925 3296
rect 22989 3232 23005 3296
rect 23069 3232 23085 3296
rect 23149 3232 23157 3296
rect 22837 2208 23157 3232
rect 22837 2144 22845 2208
rect 22909 2144 22925 2208
rect 22989 2144 23005 2208
rect 23069 2144 23085 2208
rect 23149 2144 23157 2208
rect 22837 2128 23157 2144
rect 28311 4928 28631 5488
rect 28311 4864 28319 4928
rect 28383 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28631 4928
rect 28311 3840 28631 4864
rect 28311 3776 28319 3840
rect 28383 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28631 3840
rect 28311 2752 28631 3776
rect 28311 2688 28319 2752
rect 28383 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28631 2752
rect 28311 2128 28631 2688
rect 33784 5472 34104 5488
rect 33784 5408 33792 5472
rect 33856 5408 33872 5472
rect 33936 5408 33952 5472
rect 34016 5408 34032 5472
rect 34096 5408 34104 5472
rect 33784 4384 34104 5408
rect 33784 4320 33792 4384
rect 33856 4320 33872 4384
rect 33936 4320 33952 4384
rect 34016 4320 34032 4384
rect 34096 4320 34104 4384
rect 33784 3296 34104 4320
rect 39258 4928 39578 5488
rect 39258 4864 39266 4928
rect 39330 4864 39346 4928
rect 39410 4864 39426 4928
rect 39490 4864 39506 4928
rect 39570 4864 39578 4928
rect 37227 4316 37293 4317
rect 37227 4252 37228 4316
rect 37292 4252 37293 4316
rect 37227 4251 37293 4252
rect 37230 3909 37290 4251
rect 37227 3908 37293 3909
rect 37227 3844 37228 3908
rect 37292 3844 37293 3908
rect 37227 3843 37293 3844
rect 33784 3232 33792 3296
rect 33856 3232 33872 3296
rect 33936 3232 33952 3296
rect 34016 3232 34032 3296
rect 34096 3232 34104 3296
rect 33784 2208 34104 3232
rect 33784 2144 33792 2208
rect 33856 2144 33872 2208
rect 33936 2144 33952 2208
rect 34016 2144 34032 2208
rect 34096 2144 34104 2208
rect 33784 2128 34104 2144
rect 39258 3840 39578 4864
rect 39258 3776 39266 3840
rect 39330 3776 39346 3840
rect 39410 3776 39426 3840
rect 39490 3776 39506 3840
rect 39570 3776 39578 3840
rect 39258 2752 39578 3776
rect 39258 2688 39266 2752
rect 39330 2688 39346 2752
rect 39410 2688 39426 2752
rect 39490 2688 39506 2752
rect 39570 2688 39578 2752
rect 39258 2128 39578 2688
rect 44731 5472 45051 5488
rect 44731 5408 44739 5472
rect 44803 5408 44819 5472
rect 44883 5408 44899 5472
rect 44963 5408 44979 5472
rect 45043 5408 45051 5472
rect 44731 4384 45051 5408
rect 44731 4320 44739 4384
rect 44803 4320 44819 4384
rect 44883 4320 44899 4384
rect 44963 4320 44979 4384
rect 45043 4320 45051 4384
rect 44731 3296 45051 4320
rect 44731 3232 44739 3296
rect 44803 3232 44819 3296
rect 44883 3232 44899 3296
rect 44963 3232 44979 3296
rect 45043 3232 45051 3296
rect 44731 2208 45051 3232
rect 44731 2144 44739 2208
rect 44803 2144 44819 2208
rect 44883 2144 44899 2208
rect 44963 2144 44979 2208
rect 45043 2144 45051 2208
rect 44731 2128 45051 2144
use sky130_fd_sc_hd__clkbuf_1  _01_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform -1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform -1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _04_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform -1 0 34500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform -1 0 33120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _07_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _08_
timestamp 1688980957
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _09_
timestamp 1688980957
transform 1 0 11684 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _10_
timestamp 1688980957
transform 1 0 12420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _11_
timestamp 1688980957
transform 1 0 13156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _12_
timestamp 1688980957
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _13_
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _14_
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _15_
timestamp 1688980957
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _16_
timestamp 1688980957
transform -1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_
timestamp 1688980957
transform -1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _18_
timestamp 1688980957
transform -1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _19_
timestamp 1688980957
transform -1 0 17296 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _20_
timestamp 1688980957
transform -1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _21_
timestamp 1688980957
transform -1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _22_
timestamp 1688980957
transform -1 0 24932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _23_
timestamp 1688980957
transform -1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _24_
timestamp 1688980957
transform -1 0 24104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _25_
timestamp 1688980957
transform -1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _26_
timestamp 1688980957
transform -1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _27_
timestamp 1688980957
transform -1 0 23184 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp 1688980957
transform -1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp 1688980957
transform -1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _30_
timestamp 1688980957
transform -1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _31_
timestamp 1688980957
transform -1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _32_
timestamp 1688980957
transform -1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _33_
timestamp 1688980957
transform -1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _34_
timestamp 1688980957
transform -1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 12144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _42_
timestamp 1688980957
transform -1 0 29992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _43_
timestamp 1688980957
transform -1 0 29256 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _44_
timestamp 1688980957
transform -1 0 28704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _45_
timestamp 1688980957
transform -1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _46_
timestamp 1688980957
transform -1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _47_
timestamp 1688980957
transform -1 0 26312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _48_
timestamp 1688980957
transform -1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform 1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 15548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 17112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _56_
timestamp 1688980957
transform -1 0 28428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _57_
timestamp 1688980957
transform -1 0 28152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _58_
timestamp 1688980957
transform -1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1688980957
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1688980957
transform 1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1688980957
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1688980957
transform 1 0 31464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1688980957
transform 1 0 32476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1688980957
transform -1 0 32108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform -1 0 32476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform -1 0 31740 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1688980957
transform -1 0 31464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1688980957
transform -1 0 31096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1688980957
transform -1 0 35696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1688980957
transform -1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _77_
timestamp 1688980957
transform 1 0 26680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _78_
timestamp 1688980957
transform 1 0 26404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _79_
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1688980957
transform -1 0 39376 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1688980957
transform -1 0 40112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1688980957
transform -1 0 40848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1688980957
transform -1 0 41768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1688980957
transform -1 0 42320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _85_
timestamp 1688980957
transform 1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _86_
timestamp 1688980957
transform 1 0 32752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _87_
timestamp 1688980957
transform 1 0 32200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _88_
timestamp 1688980957
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _89_
timestamp 1688980957
transform -1 0 34224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _90_
timestamp 1688980957
transform -1 0 35328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _91_
timestamp 1688980957
transform -1 0 35052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _92_
timestamp 1688980957
transform -1 0 35604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _93_
timestamp 1688980957
transform -1 0 35880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_61
timestamp 1688980957
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_75
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_89
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_116
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_129
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1688980957
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_172
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_185
timestamp 1688980957
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_201
timestamp 1688980957
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_213
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_228
timestamp 1688980957
transform 1 0 22080 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_241
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_257
timestamp 1688980957
transform 1 0 24748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_261
timestamp 1688980957
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_273
timestamp 1688980957
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_284
timestamp 1688980957
transform 1 0 27232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_297
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_301
timestamp 1688980957
transform 1 0 28796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_313
timestamp 1688980957
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_317
timestamp 1688980957
transform 1 0 30268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_325
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_332
timestamp 1688980957
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_356
timestamp 1688980957
transform 1 0 33856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_372
timestamp 1688980957
transform 1 0 35328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_380
timestamp 1688980957
transform 1 0 36064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_388
timestamp 1688980957
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_412
timestamp 1688980957
transform 1 0 39008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_428
timestamp 1688980957
transform 1 0 40480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_436
timestamp 1688980957
transform 1 0 41216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_444
timestamp 1688980957
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_468
timestamp 1688980957
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_472
timestamp 1688980957
transform 1 0 44528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_7
timestamp 1688980957
transform 1 0 1748 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_13
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_18
timestamp 1688980957
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_40
timestamp 1688980957
transform 1 0 4784 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_50
timestamp 1688980957
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_103
timestamp 1688980957
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_129
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_141
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_177
timestamp 1688980957
transform 1 0 17388 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_201
timestamp 1688980957
transform 1 0 19596 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_213 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_221
timestamp 1688980957
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_252
timestamp 1688980957
transform 1 0 24288 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_260
timestamp 1688980957
transform 1 0 25024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_266
timestamp 1688980957
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_270
timestamp 1688980957
transform 1 0 25944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_274
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_284
timestamp 1688980957
transform 1 0 27232 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_290
timestamp 1688980957
transform 1 0 27784 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_302
timestamp 1688980957
transform 1 0 28888 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_314
timestamp 1688980957
transform 1 0 29992 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_326
timestamp 1688980957
transform 1 0 31096 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_334
timestamp 1688980957
transform 1 0 31832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_350
timestamp 1688980957
transform 1 0 33304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_362
timestamp 1688980957
transform 1 0 34408 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_369
timestamp 1688980957
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_381
timestamp 1688980957
transform 1 0 36156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_389
timestamp 1688980957
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_161
timestamp 1688980957
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_166
timestamp 1688980957
transform 1 0 16376 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_178
timestamp 1688980957
transform 1 0 17480 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_190
timestamp 1688980957
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_281
timestamp 1688980957
transform 1 0 26956 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_293
timestamp 1688980957
transform 1 0 28060 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_305
timestamp 1688980957
transform 1 0 29164 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_329
timestamp 1688980957
transform 1 0 31372 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_356
timestamp 1688980957
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_90
timestamp 1688980957
transform 1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_99
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_119
timestamp 1688980957
transform 1 0 12052 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_130
timestamp 1688980957
transform 1 0 13064 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_138
timestamp 1688980957
transform 1 0 13800 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_153
timestamp 1688980957
transform 1 0 15180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_165
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_176
timestamp 1688980957
transform 1 0 17296 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_180
timestamp 1688980957
transform 1 0 17664 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_199
timestamp 1688980957
transform 1 0 19412 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_203
timestamp 1688980957
transform 1 0 19780 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_207
timestamp 1688980957
transform 1 0 20148 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_211
timestamp 1688980957
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_278
timestamp 1688980957
transform 1 0 26680 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_388
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_416
timestamp 1688980957
transform 1 0 39376 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_420
timestamp 1688980957
transform 1 0 39744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_424
timestamp 1688980957
transform 1 0 40112 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_428
timestamp 1688980957
transform 1 0 40480 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_432
timestamp 1688980957
transform 1 0 40848 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_444
timestamp 1688980957
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 1688980957
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_219
timestamp 1688980957
transform 1 0 21252 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_223
timestamp 1688980957
transform 1 0 21620 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_246
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_271
timestamp 1688980957
transform 1 0 26036 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_275
timestamp 1688980957
transform 1 0 26404 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_287
timestamp 1688980957
transform 1 0 27508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_300
timestamp 1688980957
transform 1 0 28704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1688980957
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_314
timestamp 1688980957
transform 1 0 29992 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_322
timestamp 1688980957
transform 1 0 30728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_326
timestamp 1688980957
transform 1 0 31096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_337
timestamp 1688980957
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_341
timestamp 1688980957
transform 1 0 32476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_348
timestamp 1688980957
transform 1 0 33120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_356
timestamp 1688980957
transform 1 0 33856 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_442
timestamp 1688980957
transform 1 0 41768 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_448
timestamp 1688980957
transform 1 0 42320 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_460
timestamp 1688980957
transform 1 0 43424 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_472
timestamp 1688980957
transform 1 0 44528 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_29
timestamp 1688980957
transform 1 0 3772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_41
timestamp 1688980957
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_85
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_197
timestamp 1688980957
transform 1 0 19228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_216
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_309
timestamp 1688980957
transform 1 0 29532 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_389
timestamp 1688980957
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_439
timestamp 1688980957
transform 1 0 41492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1688980957
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1688980957
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1688980957
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 20424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform -1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 23184 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 23736 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 24380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 24656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 24932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 25208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 25484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform -1 0 26036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 28612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform -1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 26312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform -1 0 27232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform -1 0 27508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform -1 0 27784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform -1 0 28060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform -1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 28336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform -1 0 30360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform -1 0 33212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform -1 0 33488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform -1 0 33764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform -1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform 1 0 34040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform -1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform -1 0 30912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform -1 0 31188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform -1 0 31464 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform -1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform -1 0 32016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform -1 0 32384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform -1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform 1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1688980957
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1688980957
transform -1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1688980957
transform -1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1688980957
transform -1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1688980957
transform 1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1688980957
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1688980957
transform 1 0 24472 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1688980957
transform -1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1688980957
transform 1 0 25944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1688980957
transform 1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1688980957
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1688980957
transform 1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1688980957
transform 1 0 29624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output90 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35236 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 38088 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 38916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 38640 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 39192 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 39836 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 40388 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 40388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 40940 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 35788 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 36340 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 35880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 36432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 36984 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 37812 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 37536 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform -1 0 6072 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform -1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform -1 0 6624 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform -1 0 6256 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform -1 0 7176 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform -1 0 7728 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform -1 0 7176 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform -1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform -1 0 7728 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform -1 0 8832 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform -1 0 8280 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform -1 0 9384 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform -1 0 8832 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform -1 0 9568 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform -1 0 10212 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform -1 0 10120 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform -1 0 9752 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform -1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform -1 0 10304 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform -1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform -1 0 14628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform -1 0 13984 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output133
timestamp 1688980957
transform -1 0 15180 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform -1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform -1 0 14904 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform -1 0 15732 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 11224 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform -1 0 11408 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform -1 0 12328 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform -1 0 12880 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform -1 0 12328 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform -1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform -1 0 12880 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform -1 0 13432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform -1 0 15456 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output147
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output148
timestamp 1688980957
transform -1 0 18584 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output149
timestamp 1688980957
transform -1 0 19136 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output150
timestamp 1688980957
transform -1 0 19872 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output151
timestamp 1688980957
transform -1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output152
timestamp 1688980957
transform -1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output153
timestamp 1688980957
transform 1 0 15732 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output154
timestamp 1688980957
transform -1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output155
timestamp 1688980957
transform -1 0 16836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output156
timestamp 1688980957
transform -1 0 16560 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output157
timestamp 1688980957
transform -1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output158
timestamp 1688980957
transform -1 0 17940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output159
timestamp 1688980957
transform -1 0 17480 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output160
timestamp 1688980957
transform 1 0 17940 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output161
timestamp 1688980957
transform -1 0 18032 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output162
timestamp 1688980957
transform -1 0 31648 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output163
timestamp 1688980957
transform -1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output164
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output165
timestamp 1688980957
transform 1 0 33304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output166
timestamp 1688980957
transform 1 0 34040 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output167
timestamp 1688980957
transform 1 0 34776 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output168
timestamp 1688980957
transform 1 0 35512 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output169
timestamp 1688980957
transform 1 0 36248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output170
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output171
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output172
timestamp 1688980957
transform 1 0 38456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output173
timestamp 1688980957
transform 1 0 39192 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output174
timestamp 1688980957
transform 1 0 39928 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output175
timestamp 1688980957
transform 1 0 40664 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output176
timestamp 1688980957
transform 1 0 41400 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output177
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output178
timestamp 1688980957
transform 1 0 42964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output179
timestamp 1688980957
transform 1 0 43608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output180
timestamp 1688980957
transform 1 0 44068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output181
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output182
timestamp 1688980957
transform 1 0 34684 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 44896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 44896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 44896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 44896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 44896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 44896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  S_term_single_183 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 35052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_12 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_13
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_14
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_15
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_16
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_17
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_18
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_19
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 13984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 24288 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 29440 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 34592 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 39744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
<< labels >>
flabel metal2 s 34702 7840 34758 8000 0 FreeSans 224 90 0 0 Co
port 0 nsew signal tristate
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 1 nsew signal input
flabel metal2 s 8942 0 8998 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 2 nsew signal input
flabel metal2 s 9678 0 9734 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 3 nsew signal input
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 4 nsew signal input
flabel metal2 s 11150 0 11206 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 5 nsew signal input
flabel metal2 s 11886 0 11942 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 6 nsew signal input
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 7 nsew signal input
flabel metal2 s 13358 0 13414 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 8 nsew signal input
flabel metal2 s 14094 0 14150 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 9 nsew signal input
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 10 nsew signal input
flabel metal2 s 15566 0 15622 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 11 nsew signal input
flabel metal2 s 2318 0 2374 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 12 nsew signal input
flabel metal2 s 3054 0 3110 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 13 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 14 nsew signal input
flabel metal2 s 4526 0 4582 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 15 nsew signal input
flabel metal2 s 5262 0 5318 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 16 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 17 nsew signal input
flabel metal2 s 6734 0 6790 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 18 nsew signal input
flabel metal2 s 7470 0 7526 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 19 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 20 nsew signal input
flabel metal2 s 34978 7840 35034 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 21 nsew signal tristate
flabel metal2 s 37738 7840 37794 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 22 nsew signal tristate
flabel metal2 s 38014 7840 38070 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 23 nsew signal tristate
flabel metal2 s 38290 7840 38346 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 24 nsew signal tristate
flabel metal2 s 38566 7840 38622 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 25 nsew signal tristate
flabel metal2 s 38842 7840 38898 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 26 nsew signal tristate
flabel metal2 s 39118 7840 39174 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 27 nsew signal tristate
flabel metal2 s 39394 7840 39450 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 28 nsew signal tristate
flabel metal2 s 39670 7840 39726 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 29 nsew signal tristate
flabel metal2 s 39946 7840 40002 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 30 nsew signal tristate
flabel metal2 s 40222 7840 40278 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 31 nsew signal tristate
flabel metal2 s 35254 7840 35310 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 32 nsew signal tristate
flabel metal2 s 35530 7840 35586 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 33 nsew signal tristate
flabel metal2 s 35806 7840 35862 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 34 nsew signal tristate
flabel metal2 s 36082 7840 36138 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 35 nsew signal tristate
flabel metal2 s 36358 7840 36414 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 36 nsew signal tristate
flabel metal2 s 36634 7840 36690 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 37 nsew signal tristate
flabel metal2 s 36910 7840 36966 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 38 nsew signal tristate
flabel metal2 s 37186 7840 37242 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 39 nsew signal tristate
flabel metal2 s 37462 7840 37518 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 40 nsew signal tristate
flabel metal2 s 5722 7840 5778 8000 0 FreeSans 224 90 0 0 N1BEG[0]
port 41 nsew signal tristate
flabel metal2 s 5998 7840 6054 8000 0 FreeSans 224 90 0 0 N1BEG[1]
port 42 nsew signal tristate
flabel metal2 s 6274 7840 6330 8000 0 FreeSans 224 90 0 0 N1BEG[2]
port 43 nsew signal tristate
flabel metal2 s 6550 7840 6606 8000 0 FreeSans 224 90 0 0 N1BEG[3]
port 44 nsew signal tristate
flabel metal2 s 6826 7840 6882 8000 0 FreeSans 224 90 0 0 N2BEG[0]
port 45 nsew signal tristate
flabel metal2 s 7102 7840 7158 8000 0 FreeSans 224 90 0 0 N2BEG[1]
port 46 nsew signal tristate
flabel metal2 s 7378 7840 7434 8000 0 FreeSans 224 90 0 0 N2BEG[2]
port 47 nsew signal tristate
flabel metal2 s 7654 7840 7710 8000 0 FreeSans 224 90 0 0 N2BEG[3]
port 48 nsew signal tristate
flabel metal2 s 7930 7840 7986 8000 0 FreeSans 224 90 0 0 N2BEG[4]
port 49 nsew signal tristate
flabel metal2 s 8206 7840 8262 8000 0 FreeSans 224 90 0 0 N2BEG[5]
port 50 nsew signal tristate
flabel metal2 s 8482 7840 8538 8000 0 FreeSans 224 90 0 0 N2BEG[6]
port 51 nsew signal tristate
flabel metal2 s 8758 7840 8814 8000 0 FreeSans 224 90 0 0 N2BEG[7]
port 52 nsew signal tristate
flabel metal2 s 9034 7840 9090 8000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 53 nsew signal tristate
flabel metal2 s 9310 7840 9366 8000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 54 nsew signal tristate
flabel metal2 s 9586 7840 9642 8000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 55 nsew signal tristate
flabel metal2 s 9862 7840 9918 8000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 56 nsew signal tristate
flabel metal2 s 10138 7840 10194 8000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 57 nsew signal tristate
flabel metal2 s 10414 7840 10470 8000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 58 nsew signal tristate
flabel metal2 s 10690 7840 10746 8000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 59 nsew signal tristate
flabel metal2 s 10966 7840 11022 8000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 60 nsew signal tristate
flabel metal2 s 11242 7840 11298 8000 0 FreeSans 224 90 0 0 N4BEG[0]
port 61 nsew signal tristate
flabel metal2 s 14002 7840 14058 8000 0 FreeSans 224 90 0 0 N4BEG[10]
port 62 nsew signal tristate
flabel metal2 s 14278 7840 14334 8000 0 FreeSans 224 90 0 0 N4BEG[11]
port 63 nsew signal tristate
flabel metal2 s 14554 7840 14610 8000 0 FreeSans 224 90 0 0 N4BEG[12]
port 64 nsew signal tristate
flabel metal2 s 14830 7840 14886 8000 0 FreeSans 224 90 0 0 N4BEG[13]
port 65 nsew signal tristate
flabel metal2 s 15106 7840 15162 8000 0 FreeSans 224 90 0 0 N4BEG[14]
port 66 nsew signal tristate
flabel metal2 s 15382 7840 15438 8000 0 FreeSans 224 90 0 0 N4BEG[15]
port 67 nsew signal tristate
flabel metal2 s 11518 7840 11574 8000 0 FreeSans 224 90 0 0 N4BEG[1]
port 68 nsew signal tristate
flabel metal2 s 11794 7840 11850 8000 0 FreeSans 224 90 0 0 N4BEG[2]
port 69 nsew signal tristate
flabel metal2 s 12070 7840 12126 8000 0 FreeSans 224 90 0 0 N4BEG[3]
port 70 nsew signal tristate
flabel metal2 s 12346 7840 12402 8000 0 FreeSans 224 90 0 0 N4BEG[4]
port 71 nsew signal tristate
flabel metal2 s 12622 7840 12678 8000 0 FreeSans 224 90 0 0 N4BEG[5]
port 72 nsew signal tristate
flabel metal2 s 12898 7840 12954 8000 0 FreeSans 224 90 0 0 N4BEG[6]
port 73 nsew signal tristate
flabel metal2 s 13174 7840 13230 8000 0 FreeSans 224 90 0 0 N4BEG[7]
port 74 nsew signal tristate
flabel metal2 s 13450 7840 13506 8000 0 FreeSans 224 90 0 0 N4BEG[8]
port 75 nsew signal tristate
flabel metal2 s 13726 7840 13782 8000 0 FreeSans 224 90 0 0 N4BEG[9]
port 76 nsew signal tristate
flabel metal2 s 15658 7840 15714 8000 0 FreeSans 224 90 0 0 NN4BEG[0]
port 77 nsew signal tristate
flabel metal2 s 18418 7840 18474 8000 0 FreeSans 224 90 0 0 NN4BEG[10]
port 78 nsew signal tristate
flabel metal2 s 18694 7840 18750 8000 0 FreeSans 224 90 0 0 NN4BEG[11]
port 79 nsew signal tristate
flabel metal2 s 18970 7840 19026 8000 0 FreeSans 224 90 0 0 NN4BEG[12]
port 80 nsew signal tristate
flabel metal2 s 19246 7840 19302 8000 0 FreeSans 224 90 0 0 NN4BEG[13]
port 81 nsew signal tristate
flabel metal2 s 19522 7840 19578 8000 0 FreeSans 224 90 0 0 NN4BEG[14]
port 82 nsew signal tristate
flabel metal2 s 19798 7840 19854 8000 0 FreeSans 224 90 0 0 NN4BEG[15]
port 83 nsew signal tristate
flabel metal2 s 15934 7840 15990 8000 0 FreeSans 224 90 0 0 NN4BEG[1]
port 84 nsew signal tristate
flabel metal2 s 16210 7840 16266 8000 0 FreeSans 224 90 0 0 NN4BEG[2]
port 85 nsew signal tristate
flabel metal2 s 16486 7840 16542 8000 0 FreeSans 224 90 0 0 NN4BEG[3]
port 86 nsew signal tristate
flabel metal2 s 16762 7840 16818 8000 0 FreeSans 224 90 0 0 NN4BEG[4]
port 87 nsew signal tristate
flabel metal2 s 17038 7840 17094 8000 0 FreeSans 224 90 0 0 NN4BEG[5]
port 88 nsew signal tristate
flabel metal2 s 17314 7840 17370 8000 0 FreeSans 224 90 0 0 NN4BEG[6]
port 89 nsew signal tristate
flabel metal2 s 17590 7840 17646 8000 0 FreeSans 224 90 0 0 NN4BEG[7]
port 90 nsew signal tristate
flabel metal2 s 17866 7840 17922 8000 0 FreeSans 224 90 0 0 NN4BEG[8]
port 91 nsew signal tristate
flabel metal2 s 18142 7840 18198 8000 0 FreeSans 224 90 0 0 NN4BEG[9]
port 92 nsew signal tristate
flabel metal2 s 20074 7840 20130 8000 0 FreeSans 224 90 0 0 S1END[0]
port 93 nsew signal input
flabel metal2 s 20350 7840 20406 8000 0 FreeSans 224 90 0 0 S1END[1]
port 94 nsew signal input
flabel metal2 s 20626 7840 20682 8000 0 FreeSans 224 90 0 0 S1END[2]
port 95 nsew signal input
flabel metal2 s 20902 7840 20958 8000 0 FreeSans 224 90 0 0 S1END[3]
port 96 nsew signal input
flabel metal2 s 21178 7840 21234 8000 0 FreeSans 224 90 0 0 S2END[0]
port 97 nsew signal input
flabel metal2 s 21454 7840 21510 8000 0 FreeSans 224 90 0 0 S2END[1]
port 98 nsew signal input
flabel metal2 s 21730 7840 21786 8000 0 FreeSans 224 90 0 0 S2END[2]
port 99 nsew signal input
flabel metal2 s 22006 7840 22062 8000 0 FreeSans 224 90 0 0 S2END[3]
port 100 nsew signal input
flabel metal2 s 22282 7840 22338 8000 0 FreeSans 224 90 0 0 S2END[4]
port 101 nsew signal input
flabel metal2 s 22558 7840 22614 8000 0 FreeSans 224 90 0 0 S2END[5]
port 102 nsew signal input
flabel metal2 s 22834 7840 22890 8000 0 FreeSans 224 90 0 0 S2END[6]
port 103 nsew signal input
flabel metal2 s 23110 7840 23166 8000 0 FreeSans 224 90 0 0 S2END[7]
port 104 nsew signal input
flabel metal2 s 23386 7840 23442 8000 0 FreeSans 224 90 0 0 S2MID[0]
port 105 nsew signal input
flabel metal2 s 23662 7840 23718 8000 0 FreeSans 224 90 0 0 S2MID[1]
port 106 nsew signal input
flabel metal2 s 23938 7840 23994 8000 0 FreeSans 224 90 0 0 S2MID[2]
port 107 nsew signal input
flabel metal2 s 24214 7840 24270 8000 0 FreeSans 224 90 0 0 S2MID[3]
port 108 nsew signal input
flabel metal2 s 24490 7840 24546 8000 0 FreeSans 224 90 0 0 S2MID[4]
port 109 nsew signal input
flabel metal2 s 24766 7840 24822 8000 0 FreeSans 224 90 0 0 S2MID[5]
port 110 nsew signal input
flabel metal2 s 25042 7840 25098 8000 0 FreeSans 224 90 0 0 S2MID[6]
port 111 nsew signal input
flabel metal2 s 25318 7840 25374 8000 0 FreeSans 224 90 0 0 S2MID[7]
port 112 nsew signal input
flabel metal2 s 25594 7840 25650 8000 0 FreeSans 224 90 0 0 S4END[0]
port 113 nsew signal input
flabel metal2 s 28354 7840 28410 8000 0 FreeSans 224 90 0 0 S4END[10]
port 114 nsew signal input
flabel metal2 s 28630 7840 28686 8000 0 FreeSans 224 90 0 0 S4END[11]
port 115 nsew signal input
flabel metal2 s 28906 7840 28962 8000 0 FreeSans 224 90 0 0 S4END[12]
port 116 nsew signal input
flabel metal2 s 29182 7840 29238 8000 0 FreeSans 224 90 0 0 S4END[13]
port 117 nsew signal input
flabel metal2 s 29458 7840 29514 8000 0 FreeSans 224 90 0 0 S4END[14]
port 118 nsew signal input
flabel metal2 s 29734 7840 29790 8000 0 FreeSans 224 90 0 0 S4END[15]
port 119 nsew signal input
flabel metal2 s 25870 7840 25926 8000 0 FreeSans 224 90 0 0 S4END[1]
port 120 nsew signal input
flabel metal2 s 26146 7840 26202 8000 0 FreeSans 224 90 0 0 S4END[2]
port 121 nsew signal input
flabel metal2 s 26422 7840 26478 8000 0 FreeSans 224 90 0 0 S4END[3]
port 122 nsew signal input
flabel metal2 s 26698 7840 26754 8000 0 FreeSans 224 90 0 0 S4END[4]
port 123 nsew signal input
flabel metal2 s 26974 7840 27030 8000 0 FreeSans 224 90 0 0 S4END[5]
port 124 nsew signal input
flabel metal2 s 27250 7840 27306 8000 0 FreeSans 224 90 0 0 S4END[6]
port 125 nsew signal input
flabel metal2 s 27526 7840 27582 8000 0 FreeSans 224 90 0 0 S4END[7]
port 126 nsew signal input
flabel metal2 s 27802 7840 27858 8000 0 FreeSans 224 90 0 0 S4END[8]
port 127 nsew signal input
flabel metal2 s 28078 7840 28134 8000 0 FreeSans 224 90 0 0 S4END[9]
port 128 nsew signal input
flabel metal2 s 30010 7840 30066 8000 0 FreeSans 224 90 0 0 SS4END[0]
port 129 nsew signal input
flabel metal2 s 32770 7840 32826 8000 0 FreeSans 224 90 0 0 SS4END[10]
port 130 nsew signal input
flabel metal2 s 33046 7840 33102 8000 0 FreeSans 224 90 0 0 SS4END[11]
port 131 nsew signal input
flabel metal2 s 33322 7840 33378 8000 0 FreeSans 224 90 0 0 SS4END[12]
port 132 nsew signal input
flabel metal2 s 33598 7840 33654 8000 0 FreeSans 224 90 0 0 SS4END[13]
port 133 nsew signal input
flabel metal2 s 33874 7840 33930 8000 0 FreeSans 224 90 0 0 SS4END[14]
port 134 nsew signal input
flabel metal2 s 34150 7840 34206 8000 0 FreeSans 224 90 0 0 SS4END[15]
port 135 nsew signal input
flabel metal2 s 30286 7840 30342 8000 0 FreeSans 224 90 0 0 SS4END[1]
port 136 nsew signal input
flabel metal2 s 30562 7840 30618 8000 0 FreeSans 224 90 0 0 SS4END[2]
port 137 nsew signal input
flabel metal2 s 30838 7840 30894 8000 0 FreeSans 224 90 0 0 SS4END[3]
port 138 nsew signal input
flabel metal2 s 31114 7840 31170 8000 0 FreeSans 224 90 0 0 SS4END[4]
port 139 nsew signal input
flabel metal2 s 31390 7840 31446 8000 0 FreeSans 224 90 0 0 SS4END[5]
port 140 nsew signal input
flabel metal2 s 31666 7840 31722 8000 0 FreeSans 224 90 0 0 SS4END[6]
port 141 nsew signal input
flabel metal2 s 31942 7840 31998 8000 0 FreeSans 224 90 0 0 SS4END[7]
port 142 nsew signal input
flabel metal2 s 32218 7840 32274 8000 0 FreeSans 224 90 0 0 SS4END[8]
port 143 nsew signal input
flabel metal2 s 32494 7840 32550 8000 0 FreeSans 224 90 0 0 SS4END[9]
port 144 nsew signal input
flabel metal2 s 16302 0 16358 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN0
port 145 nsew signal input
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN1
port 146 nsew signal input
flabel metal2 s 17774 0 17830 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN10
port 147 nsew signal input
flabel metal2 s 18510 0 18566 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN11
port 148 nsew signal input
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN12
port 149 nsew signal input
flabel metal2 s 19982 0 20038 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN13
port 150 nsew signal input
flabel metal2 s 20718 0 20774 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN14
port 151 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN15
port 152 nsew signal input
flabel metal2 s 22190 0 22246 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN16
port 153 nsew signal input
flabel metal2 s 22926 0 22982 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN17
port 154 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN18
port 155 nsew signal input
flabel metal2 s 24398 0 24454 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN19
port 156 nsew signal input
flabel metal2 s 25134 0 25190 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN2
port 157 nsew signal input
flabel metal2 s 25870 0 25926 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN3
port 158 nsew signal input
flabel metal2 s 26606 0 26662 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN4
port 159 nsew signal input
flabel metal2 s 27342 0 27398 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN5
port 160 nsew signal input
flabel metal2 s 28078 0 28134 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN6
port 161 nsew signal input
flabel metal2 s 28814 0 28870 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN7
port 162 nsew signal input
flabel metal2 s 29550 0 29606 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN8
port 163 nsew signal input
flabel metal2 s 30286 0 30342 160 0 FreeSans 224 90 0 0 UIO_BOT_UIN9
port 164 nsew signal input
flabel metal2 s 31022 0 31078 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT0
port 165 nsew signal tristate
flabel metal2 s 31758 0 31814 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT1
port 166 nsew signal tristate
flabel metal2 s 32494 0 32550 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT10
port 167 nsew signal tristate
flabel metal2 s 33230 0 33286 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT11
port 168 nsew signal tristate
flabel metal2 s 33966 0 34022 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT12
port 169 nsew signal tristate
flabel metal2 s 34702 0 34758 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT13
port 170 nsew signal tristate
flabel metal2 s 35438 0 35494 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT14
port 171 nsew signal tristate
flabel metal2 s 36174 0 36230 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT15
port 172 nsew signal tristate
flabel metal2 s 36910 0 36966 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT16
port 173 nsew signal tristate
flabel metal2 s 37646 0 37702 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT17
port 174 nsew signal tristate
flabel metal2 s 38382 0 38438 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT18
port 175 nsew signal tristate
flabel metal2 s 39118 0 39174 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT19
port 176 nsew signal tristate
flabel metal2 s 39854 0 39910 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT2
port 177 nsew signal tristate
flabel metal2 s 40590 0 40646 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT3
port 178 nsew signal tristate
flabel metal2 s 41326 0 41382 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT4
port 179 nsew signal tristate
flabel metal2 s 42062 0 42118 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT5
port 180 nsew signal tristate
flabel metal2 s 42798 0 42854 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT6
port 181 nsew signal tristate
flabel metal2 s 43534 0 43590 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT7
port 182 nsew signal tristate
flabel metal2 s 44270 0 44326 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT8
port 183 nsew signal tristate
flabel metal2 s 45006 0 45062 160 0 FreeSans 224 90 0 0 UIO_BOT_UOUT9
port 184 nsew signal tristate
flabel metal2 s 846 0 902 160 0 FreeSans 224 90 0 0 UserCLK
port 185 nsew signal input
flabel metal2 s 34426 7840 34482 8000 0 FreeSans 224 90 0 0 UserCLKo
port 186 nsew signal tristate
flabel metal4 s 6417 2128 6737 5488 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 17364 2128 17684 5488 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 28311 2128 28631 5488 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 39258 2128 39578 5488 0 FreeSans 1920 90 0 0 vccd1
port 187 nsew power bidirectional
flabel metal4 s 11890 2128 12210 5488 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
flabel metal4 s 22837 2128 23157 5488 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
flabel metal4 s 33784 2128 34104 5488 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
flabel metal4 s 44731 2128 45051 5488 0 FreeSans 1920 90 0 0 vssd1
port 188 nsew ground bidirectional
rlabel metal1 23000 4896 23000 4896 0 vccd1
rlabel via1 23077 5440 23077 5440 0 vssd1
rlabel metal2 1709 68 1709 68 0 FrameStrobe[0]
rlabel metal2 9023 68 9023 68 0 FrameStrobe[10]
rlabel metal2 9759 68 9759 68 0 FrameStrobe[11]
rlabel metal2 10495 68 10495 68 0 FrameStrobe[12]
rlabel metal2 11369 68 11369 68 0 FrameStrobe[13]
rlabel metal2 11861 68 11861 68 0 FrameStrobe[14]
rlabel metal2 12703 68 12703 68 0 FrameStrobe[15]
rlabel metal2 13439 68 13439 68 0 FrameStrobe[16]
rlabel metal2 14175 68 14175 68 0 FrameStrobe[17]
rlabel metal2 14911 68 14911 68 0 FrameStrobe[18]
rlabel metal2 15594 1248 15594 1248 0 FrameStrobe[19]
rlabel metal2 2445 68 2445 68 0 FrameStrobe[1]
rlabel metal2 3273 68 3273 68 0 FrameStrobe[2]
rlabel metal2 3871 68 3871 68 0 FrameStrobe[3]
rlabel metal2 4501 68 4501 68 0 FrameStrobe[4]
rlabel metal2 5389 68 5389 68 0 FrameStrobe[5]
rlabel metal2 6125 68 6125 68 0 FrameStrobe[6]
rlabel metal2 6815 68 6815 68 0 FrameStrobe[7]
rlabel metal2 7643 68 7643 68 0 FrameStrobe[8]
rlabel metal2 8234 1248 8234 1248 0 FrameStrobe[9]
rlabel metal2 35006 6640 35006 6640 0 FrameStrobe_O[0]
rlabel metal2 37766 6368 37766 6368 0 FrameStrobe_O[10]
rlabel metal2 38141 7956 38141 7956 0 FrameStrobe_O[11]
rlabel metal2 38318 6368 38318 6368 0 FrameStrobe_O[12]
rlabel metal2 38594 6334 38594 6334 0 FrameStrobe_O[13]
rlabel metal2 38969 7956 38969 7956 0 FrameStrobe_O[14]
rlabel metal2 39146 6589 39146 6589 0 FrameStrobe_O[15]
rlabel metal2 39521 7956 39521 7956 0 FrameStrobe_O[16]
rlabel metal2 39797 7956 39797 7956 0 FrameStrobe_O[17]
rlabel metal2 39974 6725 39974 6725 0 FrameStrobe_O[18]
rlabel metal2 40250 6368 40250 6368 0 FrameStrobe_O[19]
rlabel metal2 35381 7956 35381 7956 0 FrameStrobe_O[1]
rlabel metal2 35657 7956 35657 7956 0 FrameStrobe_O[2]
rlabel metal2 35834 6368 35834 6368 0 FrameStrobe_O[3]
rlabel metal2 36110 7065 36110 7065 0 FrameStrobe_O[4]
rlabel metal2 36485 7956 36485 7956 0 FrameStrobe_O[5]
rlabel metal2 36662 6368 36662 6368 0 FrameStrobe_O[6]
rlabel metal2 36938 6470 36938 6470 0 FrameStrobe_O[7]
rlabel metal2 37214 6725 37214 6725 0 FrameStrobe_O[8]
rlabel metal2 37589 7956 37589 7956 0 FrameStrobe_O[9]
rlabel metal2 5750 6334 5750 6334 0 N1BEG[0]
rlabel metal1 5750 5338 5750 5338 0 N1BEG[1]
rlabel metal2 6302 6334 6302 6334 0 N1BEG[2]
rlabel metal1 6210 5134 6210 5134 0 N1BEG[3]
rlabel metal2 6854 6334 6854 6334 0 N2BEG[0]
rlabel metal2 7229 7956 7229 7956 0 N2BEG[1]
rlabel metal1 7084 5338 7084 5338 0 N2BEG[2]
rlabel metal2 7781 7956 7781 7956 0 N2BEG[3]
rlabel metal1 7728 5338 7728 5338 0 N2BEG[4]
rlabel metal2 8234 6368 8234 6368 0 N2BEG[5]
rlabel metal1 8280 5338 8280 5338 0 N2BEG[6]
rlabel metal2 8839 7956 8839 7956 0 N2BEG[7]
rlabel metal1 8832 5338 8832 5338 0 N2BEGb[0]
rlabel metal2 9338 6368 9338 6368 0 N2BEGb[1]
rlabel metal2 9614 6028 9614 6028 0 N2BEGb[2]
rlabel metal2 9890 6368 9890 6368 0 N2BEGb[3]
rlabel metal1 9844 5338 9844 5338 0 N2BEGb[4]
rlabel metal2 10442 6368 10442 6368 0 N2BEGb[5]
rlabel metal1 10212 5134 10212 5134 0 N2BEGb[6]
rlabel metal2 10994 6368 10994 6368 0 N2BEGb[7]
rlabel metal1 10948 5338 10948 5338 0 N4BEG[0]
rlabel metal2 14030 6368 14030 6368 0 N4BEG[10]
rlabel metal1 14030 5338 14030 5338 0 N4BEG[11]
rlabel metal2 14635 7956 14635 7956 0 N4BEG[12]
rlabel metal2 14858 6334 14858 6334 0 N4BEG[13]
rlabel metal1 14904 5338 14904 5338 0 N4BEG[14]
rlabel metal2 15410 6334 15410 6334 0 N4BEG[15]
rlabel metal2 11493 7956 11493 7956 0 N4BEG[1]
rlabel metal1 11316 5134 11316 5134 0 N4BEG[2]
rlabel metal2 12197 7956 12197 7956 0 N4BEG[3]
rlabel metal2 12466 5151 12466 5151 0 N4BEG[4]
rlabel metal2 12597 7956 12597 7956 0 N4BEG[5]
rlabel metal2 12926 6368 12926 6368 0 N4BEG[6]
rlabel metal1 12926 5338 12926 5338 0 N4BEG[7]
rlabel metal2 13531 7956 13531 7956 0 N4BEG[8]
rlabel metal1 13478 4998 13478 4998 0 N4BEG[9]
rlabel metal1 15456 5338 15456 5338 0 NN4BEG[0]
rlabel metal2 18446 6368 18446 6368 0 NN4BEG[10]
rlabel metal1 18538 5338 18538 5338 0 NN4BEG[11]
rlabel metal2 18906 6647 18906 6647 0 NN4BEG[12]
rlabel metal2 19274 6606 19274 6606 0 NN4BEG[13]
rlabel metal2 19550 6640 19550 6640 0 NN4BEG[14]
rlabel metal2 19826 7201 19826 7201 0 NN4BEG[15]
rlabel metal2 15962 6368 15962 6368 0 NN4BEG[1]
rlabel metal1 16008 5338 16008 5338 0 NN4BEG[2]
rlabel metal2 16514 6334 16514 6334 0 NN4BEG[3]
rlabel metal1 16560 5338 16560 5338 0 NN4BEG[4]
rlabel metal2 17066 6334 17066 6334 0 NN4BEG[5]
rlabel metal2 17342 7065 17342 7065 0 NN4BEG[6]
rlabel metal1 17434 5338 17434 5338 0 NN4BEG[7]
rlabel metal2 17894 6368 17894 6368 0 NN4BEG[8]
rlabel metal1 17986 5338 17986 5338 0 NN4BEG[9]
rlabel metal2 20102 6266 20102 6266 0 S1END[0]
rlabel metal2 20378 6266 20378 6266 0 S1END[1]
rlabel metal2 20654 6266 20654 6266 0 S1END[2]
rlabel metal2 20930 6521 20930 6521 0 S1END[3]
rlabel metal2 21206 6572 21206 6572 0 S2END[0]
rlabel metal2 21581 7956 21581 7956 0 S2END[1]
rlabel metal2 21758 6572 21758 6572 0 S2END[2]
rlabel metal2 22034 6572 22034 6572 0 S2END[3]
rlabel metal2 22310 6572 22310 6572 0 S2END[4]
rlabel metal2 22586 7269 22586 7269 0 S2END[5]
rlabel metal2 22862 7269 22862 7269 0 S2END[6]
rlabel metal2 23138 7269 23138 7269 0 S2END[7]
rlabel metal2 23414 6725 23414 6725 0 S2MID[0]
rlabel metal2 23690 6793 23690 6793 0 S2MID[1]
rlabel metal2 23966 6572 23966 6572 0 S2MID[2]
rlabel metal2 24242 7269 24242 7269 0 S2MID[3]
rlabel metal2 24617 7956 24617 7956 0 S2MID[4]
rlabel metal2 24794 6640 24794 6640 0 S2MID[5]
rlabel metal2 25070 6538 25070 6538 0 S2MID[6]
rlabel metal2 25346 6606 25346 6606 0 S2MID[7]
rlabel metal2 25721 7956 25721 7956 0 S4END[0]
rlabel metal2 28382 6606 28382 6606 0 S4END[10]
rlabel metal2 28658 7269 28658 7269 0 S4END[11]
rlabel metal2 25997 7956 25997 7956 0 S4END[1]
rlabel metal2 26174 6572 26174 6572 0 S4END[2]
rlabel metal2 26450 6572 26450 6572 0 S4END[3]
rlabel metal2 26726 6572 26726 6572 0 S4END[4]
rlabel metal2 27002 6606 27002 6606 0 S4END[5]
rlabel metal2 27377 7956 27377 7956 0 S4END[6]
rlabel metal2 27554 6640 27554 6640 0 S4END[7]
rlabel metal2 27830 6538 27830 6538 0 S4END[8]
rlabel metal2 28106 7252 28106 7252 0 S4END[9]
rlabel metal2 30091 7956 30091 7956 0 SS4END[0]
rlabel metal2 32798 6572 32798 6572 0 SS4END[10]
rlabel metal2 33074 6572 33074 6572 0 SS4END[11]
rlabel metal2 33449 7956 33449 7956 0 SS4END[12]
rlabel metal2 33626 6572 33626 6572 0 SS4END[13]
rlabel metal2 34001 7956 34001 7956 0 SS4END[14]
rlabel metal2 34277 7956 34277 7956 0 SS4END[15]
rlabel metal2 30314 6572 30314 6572 0 SS4END[1]
rlabel metal2 30643 7956 30643 7956 0 SS4END[2]
rlabel metal2 30866 6572 30866 6572 0 SS4END[3]
rlabel metal2 31195 7956 31195 7956 0 SS4END[4]
rlabel metal2 31471 7956 31471 7956 0 SS4END[5]
rlabel metal2 31694 6572 31694 6572 0 SS4END[6]
rlabel metal2 32069 7956 32069 7956 0 SS4END[7]
rlabel metal2 32246 6572 32246 6572 0 SS4END[8]
rlabel metal2 32522 6572 32522 6572 0 SS4END[9]
rlabel metal2 16606 1921 16606 1921 0 UIO_BOT_UIN0
rlabel metal2 17066 1248 17066 1248 0 UIO_BOT_UIN1
rlabel metal2 17802 1248 17802 1248 0 UIO_BOT_UIN10
rlabel metal2 18538 1248 18538 1248 0 UIO_BOT_UIN11
rlabel metal2 19274 1248 19274 1248 0 UIO_BOT_UIN12
rlabel metal2 20155 68 20155 68 0 UIO_BOT_UIN13
rlabel metal2 20891 68 20891 68 0 UIO_BOT_UIN14
rlabel metal2 21482 1248 21482 1248 0 UIO_BOT_UIN15
rlabel metal2 22218 1248 22218 1248 0 UIO_BOT_UIN16
rlabel metal2 23099 68 23099 68 0 UIO_BOT_UIN17
rlabel metal2 23690 1248 23690 1248 0 UIO_BOT_UIN18
rlabel metal2 24571 68 24571 68 0 UIO_BOT_UIN19
rlabel metal2 25162 1248 25162 1248 0 UIO_BOT_UIN2
rlabel metal2 26043 68 26043 68 0 UIO_BOT_UIN3
rlabel metal2 26634 1248 26634 1248 0 UIO_BOT_UIN4
rlabel metal2 27469 68 27469 68 0 UIO_BOT_UIN5
rlabel metal2 28106 1248 28106 1248 0 UIO_BOT_UIN6
rlabel metal2 28842 1248 28842 1248 0 UIO_BOT_UIN7
rlabel metal2 29723 68 29723 68 0 UIO_BOT_UIN8
rlabel metal2 30314 1248 30314 1248 0 UIO_BOT_UIN9
rlabel metal2 31103 68 31103 68 0 UIO_BOT_UOUT0
rlabel metal2 31977 68 31977 68 0 UIO_BOT_UOUT1
rlabel metal2 32522 1180 32522 1180 0 UIO_BOT_UOUT10
rlabel metal2 33403 68 33403 68 0 UIO_BOT_UOUT11
rlabel metal2 34139 68 34139 68 0 UIO_BOT_UOUT12
rlabel metal2 34875 68 34875 68 0 UIO_BOT_UOUT13
rlabel metal2 35657 68 35657 68 0 UIO_BOT_UOUT14
rlabel metal2 36347 68 36347 68 0 UIO_BOT_UOUT15
rlabel metal2 37083 68 37083 68 0 UIO_BOT_UOUT16
rlabel metal2 37865 68 37865 68 0 UIO_BOT_UOUT17
rlabel metal2 38410 1180 38410 1180 0 UIO_BOT_UOUT18
rlabel metal2 39291 68 39291 68 0 UIO_BOT_UOUT19
rlabel metal2 39882 1180 39882 1180 0 UIO_BOT_UOUT2
rlabel metal2 40763 68 40763 68 0 UIO_BOT_UOUT3
rlabel metal2 41354 1180 41354 1180 0 UIO_BOT_UOUT4
rlabel metal2 42090 143 42090 143 0 UIO_BOT_UOUT5
rlabel metal2 43017 68 43017 68 0 UIO_BOT_UOUT6
rlabel metal2 43707 68 43707 68 0 UIO_BOT_UOUT7
rlabel metal2 44298 1452 44298 1452 0 UIO_BOT_UOUT8
rlabel metal2 44843 68 44843 68 0 UIO_BOT_UOUT9
rlabel metal2 874 1554 874 1554 0 UserCLK
rlabel metal2 34454 6725 34454 6725 0 UserCLKo
rlabel metal1 1932 2618 1932 2618 0 net1
rlabel metal1 15318 2618 15318 2618 0 net10
rlabel metal1 40710 4590 40710 4590 0 net100
rlabel metal2 35282 4964 35282 4964 0 net101
rlabel metal1 36478 5168 36478 5168 0 net102
rlabel metal1 35558 4488 35558 4488 0 net103
rlabel metal1 36570 4488 36570 4488 0 net104
rlabel metal1 35926 4216 35926 4216 0 net105
rlabel metal1 36662 4250 36662 4250 0 net106
rlabel metal1 36846 3978 36846 3978 0 net107
rlabel metal2 37674 4335 37674 4335 0 net108
rlabel metal1 36662 5168 36662 5168 0 net109
rlabel metal1 16054 2618 16054 2618 0 net11
rlabel metal1 20148 3910 20148 3910 0 net110
rlabel metal1 19688 4454 19688 4454 0 net111
rlabel metal2 19366 5253 19366 5253 0 net112
rlabel metal1 7222 4760 7222 4760 0 net113
rlabel metal1 7544 4590 7544 4590 0 net114
rlabel metal1 7636 4522 7636 4522 0 net115
rlabel via2 7038 5219 7038 5219 0 net116
rlabel metal2 8142 5304 8142 5304 0 net117
rlabel metal1 7682 5270 7682 5270 0 net118
rlabel metal1 9108 4590 9108 4590 0 net119
rlabel metal1 2668 3162 2668 3162 0 net12
rlabel metal1 8786 5270 8786 5270 0 net120
rlabel via2 11270 4165 11270 4165 0 net121
rlabel metal2 12466 4488 12466 4488 0 net122
rlabel metal3 12420 4488 12420 4488 0 net123
rlabel metal1 21574 4454 21574 4454 0 net124
rlabel metal1 21298 4794 21298 4794 0 net125
rlabel metal1 9614 5134 9614 5134 0 net126
rlabel metal1 18814 4488 18814 4488 0 net127
rlabel metal2 20838 4046 20838 4046 0 net128
rlabel metal1 10856 4250 10856 4250 0 net129
rlabel metal2 3634 1802 3634 1802 0 net13
rlabel metal2 11178 4726 11178 4726 0 net130
rlabel metal1 14720 4590 14720 4590 0 net131
rlabel metal2 15226 4199 15226 4199 0 net132
rlabel metal2 15042 4641 15042 4641 0 net133
rlabel metal1 15732 4250 15732 4250 0 net134
rlabel metal1 15456 3706 15456 3706 0 net135
rlabel metal1 15686 3910 15686 3910 0 net136
rlabel metal1 11408 4590 11408 4590 0 net137
rlabel metal1 11776 4250 11776 4250 0 net138
rlabel metal2 12282 4250 12282 4250 0 net139
rlabel metal2 35190 5440 35190 5440 0 net14
rlabel metal2 12742 3842 12742 3842 0 net140
rlabel metal1 13340 4250 13340 4250 0 net141
rlabel via2 13294 4539 13294 4539 0 net142
rlabel metal1 13202 5270 13202 5270 0 net143
rlabel metal1 13846 4624 13846 4624 0 net144
rlabel metal1 13202 2856 13202 2856 0 net145
rlabel metal1 15456 3162 15456 3162 0 net146
rlabel metal2 18630 4386 18630 4386 0 net147
rlabel metal2 18906 4726 18906 4726 0 net148
rlabel metal1 19090 4250 19090 4250 0 net149
rlabel via2 4738 2499 4738 2499 0 net15
rlabel metal1 19642 4250 19642 4250 0 net150
rlabel metal1 25346 4794 25346 4794 0 net151
rlabel metal2 21942 4760 21942 4760 0 net152
rlabel metal1 15778 3162 15778 3162 0 net153
rlabel metal1 17066 3162 17066 3162 0 net154
rlabel metal1 16790 3162 16790 3162 0 net155
rlabel metal2 22034 4947 22034 4947 0 net156
rlabel metal1 21574 4216 21574 4216 0 net157
rlabel via2 27646 4811 27646 4811 0 net158
rlabel metal2 17802 4726 17802 4726 0 net159
rlabel metal1 20700 1190 20700 1190 0 net16
rlabel metal2 18078 4420 18078 4420 0 net160
rlabel metal1 18124 3978 18124 3978 0 net161
rlabel metal2 31510 2890 31510 2890 0 net162
rlabel metal2 32522 2618 32522 2618 0 net163
rlabel metal1 32614 2346 32614 2346 0 net164
rlabel metal1 32706 4454 32706 4454 0 net165
rlabel metal1 33856 2414 33856 2414 0 net166
rlabel metal1 34730 2414 34730 2414 0 net167
rlabel metal1 35006 2346 35006 2346 0 net168
rlabel metal1 35880 3978 35880 3978 0 net169
rlabel via2 5934 2397 5934 2397 0 net17
rlabel metal1 37030 3910 37030 3910 0 net170
rlabel metal1 37950 2448 37950 2448 0 net171
rlabel metal1 38594 2516 38594 2516 0 net172
rlabel metal1 26358 2516 26358 2516 0 net173
rlabel metal1 39514 3910 39514 3910 0 net174
rlabel metal1 40250 3910 40250 3910 0 net175
rlabel metal1 41492 2414 41492 2414 0 net176
rlabel metal1 42136 2414 42136 2414 0 net177
rlabel metal1 42918 2414 42918 2414 0 net178
rlabel metal1 43470 2414 43470 2414 0 net179
rlabel metal2 7130 2057 7130 2057 0 net18
rlabel metal1 35926 3026 35926 3026 0 net180
rlabel metal1 39790 2958 39790 2958 0 net181
rlabel metal1 34224 3706 34224 3706 0 net182
rlabel metal2 34822 6375 34822 6375 0 net183
rlabel metal1 20286 2040 20286 2040 0 net19
rlabel metal2 9246 2057 9246 2057 0 net2
rlabel metal2 8510 2125 8510 2125 0 net20
rlabel metal1 17250 4012 17250 4012 0 net21
rlabel metal1 19550 4624 19550 4624 0 net22
rlabel metal1 19918 4590 19918 4590 0 net23
rlabel metal1 20700 4114 20700 4114 0 net24
rlabel metal2 12650 3774 12650 3774 0 net25
rlabel metal1 21160 4114 21160 4114 0 net26
rlabel metal1 21022 4590 21022 4590 0 net27
rlabel metal1 21574 4658 21574 4658 0 net28
rlabel metal1 22011 4590 22011 4590 0 net29
rlabel metal1 10166 2618 10166 2618 0 net3
rlabel metal1 22218 4624 22218 4624 0 net30
rlabel metal1 22632 4590 22632 4590 0 net31
rlabel metal1 22862 4624 22862 4624 0 net32
rlabel metal1 23230 4590 23230 4590 0 net33
rlabel metal1 23414 4624 23414 4624 0 net34
rlabel metal1 23782 4590 23782 4590 0 net35
rlabel metal1 24242 4590 24242 4590 0 net36
rlabel metal1 24656 4590 24656 4590 0 net37
rlabel metal1 24932 4590 24932 4590 0 net38
rlabel metal1 25208 4590 25208 4590 0 net39
rlabel metal1 10902 2618 10902 2618 0 net4
rlabel metal1 25484 4590 25484 4590 0 net40
rlabel metal1 26174 4624 26174 4624 0 net41
rlabel metal1 28106 4658 28106 4658 0 net42
rlabel metal1 28382 4624 28382 4624 0 net43
rlabel metal1 25990 4556 25990 4556 0 net44
rlabel metal1 19734 4046 19734 4046 0 net45
rlabel metal2 36570 3910 36570 3910 0 net46
rlabel metal1 19458 3604 19458 3604 0 net47
rlabel metal2 18814 3910 18814 3910 0 net48
rlabel metal2 18538 3638 18538 3638 0 net49
rlabel metal1 11776 2618 11776 2618 0 net5
rlabel metal1 18998 4012 18998 4012 0 net50
rlabel metal2 17986 3740 17986 3740 0 net51
rlabel metal1 27830 4692 27830 4692 0 net52
rlabel metal2 30498 4556 30498 4556 0 net53
rlabel metal2 41538 4845 41538 4845 0 net54
rlabel metal1 38226 3638 38226 3638 0 net55
rlabel metal1 39882 4080 39882 4080 0 net56
rlabel metal1 39146 3604 39146 3604 0 net57
rlabel metal1 32706 2924 32706 2924 0 net58
rlabel metal2 32522 4284 32522 4284 0 net59
rlabel metal1 12374 2618 12374 2618 0 net6
rlabel metal1 30728 4590 30728 4590 0 net60
rlabel metal1 31234 4624 31234 4624 0 net61
rlabel metal1 31510 4658 31510 4658 0 net62
rlabel metal1 32246 4624 32246 4624 0 net63
rlabel metal1 31832 4590 31832 4590 0 net64
rlabel metal1 32108 3026 32108 3026 0 net65
rlabel metal1 32798 3060 32798 3060 0 net66
rlabel metal1 33074 3094 33074 3094 0 net67
rlabel metal2 40158 5015 40158 5015 0 net68
rlabel metal1 16652 2618 16652 2618 0 net69
rlabel metal1 13110 2618 13110 2618 0 net7
rlabel metal1 16744 3502 16744 3502 0 net70
rlabel metal1 17434 2278 17434 2278 0 net71
rlabel metal1 18216 2618 18216 2618 0 net72
rlabel metal1 18308 2550 18308 2550 0 net73
rlabel metal2 20102 2176 20102 2176 0 net74
rlabel metal2 20838 2074 20838 2074 0 net75
rlabel metal2 21850 2108 21850 2108 0 net76
rlabel metal1 21022 2550 21022 2550 0 net77
rlabel metal1 21620 2618 21620 2618 0 net78
rlabel metal1 23782 2312 23782 2312 0 net79
rlabel metal1 13846 2618 13846 2618 0 net8
rlabel metal2 24518 2040 24518 2040 0 net80
rlabel metal1 25254 2516 25254 2516 0 net81
rlabel metal1 25760 2618 25760 2618 0 net82
rlabel metal1 26634 2618 26634 2618 0 net83
rlabel metal1 27324 2618 27324 2618 0 net84
rlabel metal1 27968 2618 27968 2618 0 net85
rlabel metal1 28796 4590 28796 4590 0 net86
rlabel metal1 29440 2618 29440 2618 0 net87
rlabel metal1 30176 2618 30176 2618 0 net88
rlabel metal2 1702 2108 1702 2108 0 net89
rlabel metal2 14398 3400 14398 3400 0 net9
rlabel metal1 34776 4726 34776 4726 0 net90
rlabel metal1 37053 4590 37053 4590 0 net91
rlabel metal2 38042 4029 38042 4029 0 net92
rlabel metal2 37766 3791 37766 3791 0 net93
rlabel metal2 39330 4267 39330 4267 0 net94
rlabel metal1 39330 5270 39330 5270 0 net95
rlabel metal2 39974 4063 39974 4063 0 net96
rlabel metal4 37260 4080 37260 4080 0 net97
rlabel metal2 38686 3961 38686 3961 0 net98
rlabel metal1 40848 5202 40848 5202 0 net99
<< properties >>
string FIXED_BBOX 0 0 46000 8000
<< end >>
